��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ٦��i ��R_�>���C1Y��?�"c��m=��h��H�V��v����[�vL#KZ�"��\���#\&W���Ӯ��d����(}H�a9:���a'�C��d�{�f �[Ge)�	r��#���ԝ���==��H�V��{!�oyؕA	��#I�bӍ��p�D�-W��c�ح�*ы������t�y}�9�*rѹ�z ,�%�}uDgt�O�����+"A9e����t>��-q2���.=��rv�Y���zX�x�2�6|����b'ɹ����-��N�~'[���v�s�t��g;��<��/\7�������;�
ڶK~�v�3,9�� F�4*�Wm�.�y(嫈L�V<qg����i����De7�D��<Y��!��X��c)�Ж��shr.��< �3���� c`V���9�`�=��+�t� bu'��]D�(�;|�%�%Dx�%�[K;B�{߈ ~l�d>�Z� $I������;�lǜw���]�ft��%�5 ֣���	�	���5)��V�;m�k��y�p��٤h�Ba�0����u�;a�?�H���Iq1��2-߸T�3*��y_ܺ*�}��/�T�<"J��*qֲnmM.Dqi����W7N-�K���:����X�WLѪ��I�㛵ehx���5��2�F��f��"s�Q��Ӣ��pg=U�6]ǇG�j��h԰��,�^t�,Z��Q�O���T��L�$&�;JK;���
g��n/e�v���zl���/3Mw�p>����v��@-�j��ț�!״K����?�^-�A��e�p,O2�A�h~6=���wVH0�{U�7��ˌ�Ǎ�����ŶQ����)�����M�Թ��+!�È��lBe���Y^<1�jXt������r`�y�b�rOQ��0�+�:@�)�$��u<�GT$3�?ӳ�e"�K����S1k��4�l�Ә=����"����hܣn:lsY��}!���'��+����~��LC���C�Y��d}�(0Ȼ���;j@=����%5r�@1	�67�u�����<t�&�վ��=�������0��8����Fl�G/o��a�q��g���7c�����\��B?�C5d��X<�#�i�����<��fr]��>��8���������$&'<�����K&�e�cё�p�a:�7������N��v�ӽ��q���`� ���O�2�ܤ��X�'�������edx����0<��4<sD��a��jГ���ථ �|����͢�LG���We�y�$�r������n��������K%6�P�N�~��8��ۡ��ҹ�؞�_��U�5�􈙯��\2��p�G���g;]"�#J��1	��5ism�%�3���(��)���T�K���2!�W'�KǬ1'y(Y���_f�VIY�I��M��=�f������V��R��L�7p��Ex�j�ˎЪ�ۄՕM��B[,{n����K���i��Pp03&$�}l E��a���$%�k[ܹ"�B�|ZCu;��VF/���9�*���� z� 7��z	[��T��5ݝ��*�B
�A�~��n|(��M'��E40�������-�qgɮ����H�-�S�ͫΤ\f%�)���Ⱦ��&+��So��e�L�	Y	�X�8_
V)��IM퓎�����-uhi@b���6�ף�c������!iF���%!��ꎣ3^N�3�ƂAR���s�J���P�PD��×��t9y���ϛ�Q���m��M�x9�z�����0�.�3i~�A� ������	��*D��;{����$#�h�oD�U�U�ض'@��
R�>�|���6�
�^<�?��1���C��
؏bt��O]�'Mɉb��$�ʈ��&L���{��<^ҕL���+��bf&6�\�Z��)O�W�u�	�{Q���J8��H<������f7����i����9��ԷP�?��O��}�7�0_�m�O���*�>$i��OZ���n�C�����OD��7�����t�1�#����a`ROX!��u�s�b�q�6��rvN�RΩP�lg)�"^	���xd�����6�_���9�Af�ޜ�	go-Sf"9���CȦ'D-�i�
����~{�kQ>�u��'�?��B�L�J�xG)��L���u)������<"~&�xR��l��jR�沃ν���uNA1�|q��H��G�C�3#B��M�e-5.�^>�� )x'�T��z��J���
I=��ʍHW6hK�ԥ3�)�IP[���8�ԣ��vӳ���R*c<$��W��9�ʹ6��o������.a���6��Y4���b���Ug׹j��&ߘ�Ä�XY�z�������Ӝ���[��xZd�����;���"�����uʲ�E��:秞G��&��~x�Ύbg ���V�c4B��V��2ؾ%��	Yw4^�Mo�s�z�~pˠ�]N:ۡ���{x��GiaS�����|�����8OrC/զ��ո�MK��U��:���De��0�D��	D/}W�,�� %��f@J*����'uю�㞠�(@�v�Y.�@c�6��x�h��>��=��l���6�-?�	�8{;����6
�dT�ܹ���p=T�ɍ��yZW��)#���ʹ8�����4Q�lf����H@�`��T��H�<ӆ�s�iyu�9s�.�v[+�2ԵM�v���E��Ž�&��v�������Av~��r�� �뤫ưø7��r���l�R_~��%;EFl&C��k�l�?����x�ΜA!�5�F�	f��7�K?Ճ��3�~�Gy���`H~� ^��PL���s���l��D_J�-\���DQ �G�pU1��[ �#`���e�"��6�4\�z�*�!���*[�����42a"��}ˌ�qٚU���[R�����Gf���O�e�T���G��W�&rX�,1�A_G��>
�>0Z�"A���+6��C�	�㍺�mnC=�#&����މ��1ꤿ�v�鷾s[��a���1%B������.��(���`@0I����YC��I�z���cBxF����=��!% ���ˀn���RIv�?��8�#����S� M�4��]��)�_�����	�ry"U��Dܖ�-<6��ۅ��S�mRZ��Ч�S���
��u�^}+��J{�g#�u���xc�m*��J_�+�����A���G�e)v�:*���g�K����i:m�Q6�������T���ПV��H�]&n{�~E���T;S�	'{���Aֹ�N(b�O�Z��S*�!�c�Q�bpv
�W>փ�D��vމW�o�K���S��)ܶ�҃� cL�gA=��Z�F�ji֨z��T����/�p��A�[m�ŗ�5[w��+�]f�h�-�X���$)��|�ݙ%�r�PnpHm�9y;�~�f*Ns#{����NƩ+)L�zdc4��'�2�wL�	�t�R���)���p�Ȁ�����met�$m/����e�^�ǀB��N�9@O� kF��:&	�+��j��(Y؇�hG�-[@9;���DlY�Bz:4��R�a �Ζ�(���R��u�K�����_˹�ʩ#A,��$�����@�f	B�KĽ�;�[�0�����H�\�DCd���Ǎ��j�9�K����2Xm����2���k#���Z ����FMH)����j�k�*�s��>;�bВ���^q���������y�땁���,�t��E�sT���VC�w2�G~�J�̽�׈���u�g�>=e
&����)ζ/�[$ʖL����������5c��N5��@O��8]\̻��f%��1�Z���c�~5UG�_�:�=Y�T���(_#��Q^W�u�08�;.�)TCS�uX7���I4���|ʁ� ौZl��ͩ�ѬaC�J�h�:��}�1uc_��G��s���Y2������*a]��"�l��Y��
 �[���.��AE4~ς_�
�^vp�#͟;�mfi��Hb�j9��w�.TvjI�K���ѵc���k"^�F�is���x�u���-=@�����i��9M�5�n�rb��+P}��b!&���F&y���81M�W⎳��Ⱦ��  ����p�`�M%Or.ˉ������蘜i�3C��w���RNcP��=�u��a��;�涷4�A���h.QV�km����ɮ�I\l�Tq	�aj�@��f��P�81��Wb# fܨ�� Ʋ���6>��l9Iy���9ɲD�a'��^~�в��c���Wm����IO��H����k��${W�G�����\��׬?��Z^�kv��:h��{!CGxB�;wZ�HO@�������tف��6�t �Rf��IՁsL3b���N�ڒ#O(����ߍ��(�ŷC�F��}}0g	P�O��7PN��+�;�N���X-�c���	�;�����{�M��B5�i��&��n�o�Rrʮ4�Y�/zc����R���a��U��lY�"[��e0hf����anM$�£�_r���)�i.�L��B���Z:�1��Q���2:�s���]��C��i\��}c����tНVgFN�q��J8�����',�G�UI$�(�3��h���Q�%(z���?��R??æ� ��}+���%R���*7W���1��٦����ѱ�:9E��}�r��b���b�1�^����N��;"U<)��E�=�ڬ�`S� �.��Y;����u�	s7�F��S�������HŤ�+�}�s����	��W��҃������!�2k�J���Dsl�M�I�U� @�a��D10�1{�/I�\"-��oc(��3S[e�z@�995�C�����a�uX��(�ȕx'��g��|�|��/j'��l�//�-~���^\z���a�Up�G[���=,I����U��I��f`�?�ҽ�U���� ��er)���"����Tg�1P�r�ǚ�c{���p��Mw����[7�|i/8�F`�Ͻu:�?GP���z��m�e�=_آH-*�gB�6s��u��$SH7<��c1�%a~Q��w�
�q-�y�*�vI\_t��a�i��.V�#'�[��9�ȸ��qm�cw�˟e�/:���D�S����7'�͚i߀+�Ld�.�F��|���;t�ī���F	!9tx��Z�����H��e�"(���	���Y[��$�`:6< OO灳�\����7p:���٪��!���E��T���}�=�p�M�����J��I8�������z�rz~=kʰ��N\���v��hh�ꚃco������`1����zpU�H?�fp 1^+H�i��h7��m�k�~�XW������g)���vT�n�Sۖ�6H�
|����'���e?uB���ϣ��3�������ci�E^��7�6�'L����OU7w .�OLT&	y��]��=���G��a�qk�cz��9����
��~m\r�8�9�;�}�#; ��m>0��'�:��ڸQ�R���h�e܎ӃLn7-	q�W_�K#$�����W�����u{�
��Q��j�֚��S�هnyK���1��0��x�����`&��k��{����e�� \u�d�rq����ia�����9<9��,��E�Zc#�.�bդsx0�N{k�~c8����j�X|7Ejۼ��sui#Vt��u�ţ�����k$7"�~���Y�I4&v�Mvk�:7�N��F\���|�6$m1��B�6�7��Ԣ��	.�u�g�bs�%�mC��W�ߊ<MX �7�^�/���Q��W��D+XYݖ�:�>\~��*EmUIE�"��鬴�(0	�N��Q�C�`��8�|����+ݔ�?�����NČ�׾�utO�ÒkN%lR}��^�m�cBn5j���z���є�8�h�
iW_OD1��d!�;g��:>�:]�R3P�^���:���{�}��C_˛=��Ē�7}O�����ޱ������D�W���u���uo�'����ͽQ�Of@�gz�e���9��C8d�(��w^���0j����o�z�#1�ԣ��)_�f��p/d��eByhs]�&�/-ޟ���V`]���[��;�Nb��a@~uز��&n����܃��i�_�{�x�!5�4�`��t�m|�������t<*�aNt�2s��}r�W|�9�us�pzU�rV�J?M�΄�Zgj >��|8ۏ���
ѫ[�����|!^�|��cţ���!On3L��CJ�����Q��D���g��p��9���Z{�c���⹆ql�G��Y-�;!I��M��{t1e�~�ODX__Cs���=�0����ptus
~GOdiT�P�L]Qg�H�8xv_�U��<폽S��R�M�A;�}��7�{�k�s�_�W��>�������9x��aQǂ��K�N	������u�t\~����`�~��,Rx2�q�5���E��l����f�RG���z}�:�E�q.�rvavܣ\�����2��]�@�s2P[�`:�
D�O���7�ӂ�Ԋ��Ք���K)�Ա�zk�ک�L�`X��$�����2����+��˲v�m+K�f�A��_7��&�SEES�ʝ�^��Nb��꺢�%��z�����l�$��.�B2��9��cFg9q�K��h�pH�/bP5�>b(�w�P��F��{zn�^ƕ]�E�����"5o6���Uׂ�1���J���NJp3��