��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ��t-�Y�
���?�O>�	�P��qC��_���b?M|/F�!v�n,Q�S,C
^� 0s���A�}����ͨ��o�d�'%9�vL��?܆э�n5�h���6��Ĕ����p�SY� �����Q���'2�rQ��'�l�psJӒ�A�MQfx�¿��ޮ�����z���"=$L���>��ۣ0��Bo{�cJ;oF|L���P�BIf��~��/��'�:�$R�d�<r9ā�Kl�͡�VfO	ǰ?p����)c�0T�h1k)�s�v���A?�e�ni�&d��#t��܈_�q�y�bc�}L\�nhd��6(\�l\T��iڄl�k?���d���A��"��ޑ�F��+��{@�.�U��a�-O�کr��6}�ܒO/�'oӖ;�������ʹ␏sm�N�+R����B� ��/����6	@8f+մ1C�%�H�2�DC0!d�՛r찳<J5*Yk����R�9ˊ����J��y�T���'�ͷG,OkQ�Wf�F��+.�۶��wA%�ʜ��(��ZN����
��4�E/�vo_�R*H�+�e�z���������}�稱�_=2琈 us��.-�;� 2M�z4�fkgH�%�^V�,�$��m�����HQmK���K��`�o�e�q	'���[1d:��ᨓ�Wl`Y� @�ڝ�C�R�<S�78tz�*��)�ˣ�
���ҩ�4����,h<��\d�Ƿ��s
�vi-��Nw��}�jc�t�-�x��xq���c�u��R"_��Y��3<�V�����yeɆ�$�I��+��a��H��@��h��L�<�0�	�/� ���dr1�$��tE@�g0�����5�;?�$+M�=��3?��MH$�nKl���r-��0���'P{��%���S�h�p����^)�F" p�(�I��س�xz��!�Lr@G�onء��h��"ӑ��P������ ��Yb(�] s��c%P:����'N�{nԪ⢍����l����/�!{�  t��Cx�kZK@�QC+<ֺ�|0A^�fr�����3д�s]�`ˡ�?�����f�ˋ���I^����B�Њ�Ē�-����-X�e��@���:Z�LCH��Z@o8(S�Cc0�n��=����t�]���l��ov�s]#ҋ=��=aNm��B����8���q$U_����V׬�5�_y���CIo�?���W�:,Oc��D�J��������
�J�]�7��f3�!�ɣ5�0pUsQOj�e�@��*&! A������9��0���v��Ll��'�0oi�S��`ݐ�y���B�?�nN��4����`a��[������l�s���Ѳ�Ǯik��h�0J�f�Q}_1��_���L|,�������5N�kf2ЛL���cO��\���O�o��u��^Uj�����L�&��H�?�2$�{qz��qډ÷�,��$�v���e+o��1�:G/����z�V훰�F��|�	K�G�:�Z��2�L��u��I�V�c� `�FA����t������{{8���,�d�*�k�8�&����qoN�<�N؀��6Ia�XgK�I`�<�&Mg�Z-O��V^]Mڞ8[�.:�|l�qy��n����w��i}��ϙ�~���5��%Ij��h:ܠ�[ی��nn��vi m��l@P��`����@Ɂ�<6m��)����zSo3�db^������$Z����2?�uoG���l�Q�_P��l2����gx�%`��ıZ�a�+A^4}�����bG����ؚ%��O�4#"�gv���z��S�?�y�w��X�D�ԙ���&��PS&��&�y�^��,�h�x[� ��G��`������BM��ϫ߉���A���MV"=z|0I�{~~�6E<��-�u$��7���s�&D����u����h�����ujͤ��>��je)�00�Z� z9W���~h �_r��fEܪ�E0��0������XHƬ6;,�Y;����s�u�/�M�Ï�I�;]���FX�b�M+\��|v\C�*7��X���4�1ن�,�	5B�I��X��=�)���L�dz|`�S<�\t���{ßG��0}>ޜ�;��3.��z��E�����@#"I���/�l���K���Np�l�U:�h��Zx�*��RE���ϧ�P��cZCl�.�˕Ny�">}���{%3�P^��R[�eg}���<�؈�~K,��Y�SCИ+��\9��Q|�s�Wb�F���Qt��Mu�.�F����ئ�=�uM�42)����O�/<�Y�2=w)�z]c��,e?LD����zy{�2~��rNC��|`I��f1_)L���Q �rsL�(�0�,�D&����A����y�����Z,�&�0G{��i�RF��W�:"�S�.�e�����dJ]�¦(;q�`���<�;�������0�|�DL~�b�s_���K�g�'F�g�%|�{�%�њ,���yG_��!����A��'�� ���j�+����
͢n��k��\�Xf�O#ǔK�@4�O^���)XݕP\�>O|q�Ld�̽_�/��֒����?Ƌ��شp��Ϣ6w��jFI�3�Hf���ұ#P�#�_%\��֢2�Ϛ���g�ŮO�sO#�4`r��<��Gʇ<P�w67���R�tgDB3�^�,��� �:#@��тY!�-@m���Ǻ����"�o���9	�ڧ�<�"�1���C����I�k����n�Zب�O��{$�|�&-܉��` ���"�p���2��k;��~ �O����#��!�p%W��y����D�NQ>�μ�:��w�"!O�N�)�7Z����j"� Q�%��4�F�~�%��JP{2����PAٴ=��g�Tep�L���Wb����[�~��
	�~��1ޕ�z���!0�F�"3��	ӫ-����󸯢$ �U$����+<9�8����IX4_kvg?U�,}�R��jӎPF���9�;��U�^�"}����c��hR>���UW"WuZB�+5����� )�7���oW�`���-�����G{}���2i�Y�Ϻ��O0�{�kÝ����p	`Z&G{��:d����F�}	�Y�A�d��SS�1�juǤ�x@�� �]��MP��/�q�L�)qP8C���1]M�S�����ފڜۧ�Q�љB�GM5�����=��c�����ޏ���d(�A�؛�j�s�i)*߄�T	����Ŀ�j")|GON����D]>9��gf:�����;��Ce�����:zm�ݭ�W����m_��:M�i*͒�D�_O�tc %Z)��e�.Ζ2��kP���@ _&����bA�ӯ����{�<��� x0��Pİ9�
~���}��"�j��g����������m8T��� 3�?��OAs%^��g���h�¯x���=� ��q����̔�V����f�9�����j����h�-i$��7�ף����?�7�Kv�<ɠDh��o��?ൣ�D�07j��̊U�!�k=�Xuq�['�Ө�o6	�F�'~����l8@��h�HuSi�#H��&ʈ�t�6�q:�ڒ��\x,(2 �z�t��j���6�B�.�/9�-�%��m��v�S{��q����{�=xT1��,��_�K�M�p�M5qo�1^MN�lsd�����Q����Ε#/I0䫃���'+]�C�w��?5
�$��C�E�7_�Y��2��e���J��,�;���
ku#���G�/��P���g-`g��C�࠾�>=�zR:�?	�;���T�;>��>�Wq>8�T�ɗ������*ĭ�5]<ھ#Q�>åO�.N�[�v�e
c���a��O �, (Z{`H2�s��(F�h_ɟ�#
l;���i��xME[��^0nۛ�ﴗK��;�{�-��]ɫ�_�F[,��|e˜���9R05g���+=��ˈ�O5��ǈ�%@��W���K$�UMT�?�����,o�1Z���aCn�&'�E�:9�1p��l]F�����+o(�r�?���>s尅R��5����qGv8� tñ����IY���A��92ka�b�Qjb�3ߙti
Օ4�`�z��
;B�H��܊�}���޻�]B��TuN����L���YJY�+���<Q�R��G#��O��4��Im_X�hi��/��"��ON<5kFK����h*!�M7!
F�l��;[����Kz\@�������c����,�=�~Ɔ��?6�y�b/�={�'���E���Ơ�nq�A�����Zu~w�B_�X3��b��Hl�ZD�@k
刿��z�Iw
kE�O�ğ�����I�b�A�F;�`�`��Vn̼]ͧ�GT� b7 �e�\��l�`��x�.3քCc�1�)�/����녪'��$��/qB-�D}��
/�ie�ig��}�!!:0a&-�>���y5S��7u��WO�x�ûB���e����Q��7�H�X�1#p�y�Lr4���Z�I�"n����"�2H�Y}U7��U�tӆ�d��B���&O���%%���*Ԥ4���9L�2HB�ﭚ��l1p3R���z:���1L/�����C2�JK�@H��@O�����n5�]H?�e�.�,R���K׌�BFo��=҃�"y��PĂ{K�YGQ�	��r�	A$�8��⇰�_��_�ej͋��C�D37���1��X�;!�`
�,�坸��K,�,�-}P��'��glz���kc4 ��5*�>������|148\� �9�>|ŉ,�F^x�,q3���IhP
>.Q3}����c/��Y�oR�d�!q6T?D�3����y�/)C����	��L�&Ԙy�7&9�W0Y�vG�ķ"C�[0{���j[>� $ :ܼo�5Uk��&�@�\�U�Վ����OL�8Z�Ͳ%C)�.����O�5�j�,�_fNI:�z�҅� }�A5BA�v}:����%C�~�A`=�-�D]~�9U57�v;L�n��=*d%lpVe������v�:Q�6@�I�|�P���m��p�5޴f�5 :��+��o����;2*џ��?s$����1�M��EC���oS�]��Ε�{��j���2�����4ژr�lS=fU���`���M�8�QgI8�\'���GkD�`�cB�p�"���\�pb+��Uz�i�/D6��X�=�Ey��p �BCl�۴����r6X}�b��!��!w������X}6��kRK)z7���;�f-%�^��
���? ����F�P>ү�Z!6���e��PU��D��eS|:�i���O!�:NɁ���W�Wdr
�r`��(&�Vv/������j����ǿ�T#7�8#,�_�ӥE�_U�ew)�j��Od�:��ńD^M%��Z<�Îo\�eٻ+�6*��;�7�mՁ�H0A"�����4r�T�\���#��</Og^͞2�$g�� lt��I1���1}�פ���d̝W���l3�7(~�\����rSEm]��J����&�����"�ƽ���n�F �9��݊p�66���(��I�y�u���g	ƍ�g�K6�>[<�6�͑c�$�]2�0)z�5k�[F�9���Q��V�=Il.'�h��ϻ�7�K�r��ԁO~e]+h�� ����x[Oדس5@��
ɮ����>C��#�2�����\J@�ȑ�d?	\݇������u�x�b3G��z�e�y�e�As�d��x[��?#����Z��m�]����ƙ��dH]t��.VIE�%N"Ǩ�qe�wi*�s���4��d'O�� ɬ_g�(l�2	�8��k��d��ي��c���!�E�7;���Y�PL���ꣽ�ʨ��2��IJ�jA��`����y��w�Lİ�<�׸ll�!)�O���!X��:���i��m9#����Pg)b��$&�R���Wc �?�l4��<�R.P[�K�v�6+.>@-�76y�v�@��`��z0k�_�T' b �l�F2����]g��q�@�=�����#v�cև�Uf���ݍa����V��V��U�P�݄eV�$���ϓ.��)���0������U[T�6���&�̤�x��xt�d�8�ڮN�?r�:�ʠU<�p,�	_���ʀk�6vrʷ���N��[��sA'@����by�uO�\Y�_�6�
��bM	�J�Q�Y��,�����������.���f$���T�X��G�[�+^�H�!�y>c�4���8ݱ��'�I������
J�[6������9k��7dƸ/�����L����B6.S^�f��cTz]	Ðr�s��GY!�`��=�L���n��C�h�J������qȮ��Y��=�ڲN�@.r��PӯP#������� �\F�f4)n������!|��as�t>�ȩ��S`���?�ϺW )<D~4��Մ���8�����9ܴ�/�<� D�lU�Q���Z�w�_r�ȷ���l��<Q٢��7w���)*G��u:�����j�c0���>��RϚ'�z#[>:�Z�CZ�ү��e��?�A"��>k�ĩ�kWɀx���^9������� *?/�wޖ����V��ѽZ�Oŵ6봡�ݴs^�^�3�cq�:���0kz��#�>�W,�M�-�2H�e�4��+��0�m>9�	�������`��2�ݥ�,,��e��W[�1E�ݣ�=wH4>�D��.�����lRn�\u"�����7K���,!�̖?.H)�U��g�aS�W�L7�G6UPv�4a��k�vӉ��o� ��4�I������HmF�@QF���������6�Z�H�[�)�=��|���&���9��H�?�78;T���(�[B����-�N���� l�ソu��t���a�[�+��,p��H�L��*����,�5��`�=v-�V$�wp�i�1�̇���(��@�d����=�td�T"ex̓1���>b�����?�)�}�F��Gjo�LDF���,��u�X�{��NCl���ŏU;|�M�u�V����߰�g�C��\��T��n��F5�]�z���փ3J`� 6(�x�#n����<�����x`&+�וlp���e�H�H�����oA������S���0�G�֙T騵�Bӎ�h~z0x`F��� ${gz#�M����G��*�ژ����h꺴���a���!�|R�-Ъ��'I(g�.2J��63`뛮��2v�A��&�g�ڻ�Җj�A8�ѳ?N���Lc�U|{�V�x���)5��A\��~
r>+Ό`E��&�QU��7���?4��F����v@��\����ŉ����r�y�����:��d��A�J+�m۟����XX8�Y�@���-�X���×,�؞���)Юc]dk[X���y�6.,dFM�"�=3��3�>3��ᵏߨ4��9"�g'<���`(H���}���6M�m�<�K�Ͱ8���n�R��_Q�F�#�΂\�y�1��q	v�F� �7��8���K��Z6-��T���k��՝�P��q�PX ݖ&� ������H��>�_�����l`����m�H�=���;�{���S�V��.6�ԪcyӉ��x����y5D�j��ʒ���i�TZv'v~PR�k20���Ln�rG�ܨ"xƻ$+Z)5�,�j�$������lP���uNvjӎl\ܓ=f%I�e7��o;  [���wu�L�Ƒ�Qovr�e�M��y��#�I�S2�I��>��y͈t��#Wء��{*2�KK���H�&Z�\A�c��8��5�t#~�vf�`LA��--t-]=�Xj�hIF��ley�I���f/ h��?�,�^RY�D�~j����:�{lPfC3�P��S��`j�#��i��xg/`��� I+C6:���� ;�u�3��͖;���o��3��[Y���zŨ��HԹ������]����b����nLp��eX�;�B:��aTZ��l���w.�k��J:�K�M˽3�C��V͐y�&в�w�=����sP���[��h~<�'�eX�¡�K0�o�)R��e