��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ���6'����*���Bjɾ�?��کm}M"�o��a�y<9M�FpmBǲZ�^0K�x�gŻ�H��+�#1��0�q!�
]v�� �CW(�敪d�σj�?����Չp��J"�k�����3�6֕ռ�}�HJ�\)̆�Q�	���8�Ƨo�
s�W�{�K�
�cK�7���p�fM/Vx�CN�\i,����p�^��%&�T�Ŗ������D�e�r�����B�L!�S����:q��X{@(�H���L�o �l�N��Ȥ��P�9��-�B���Y�rڼ%IW�1�08�"��������(�i"��#��{��YeA�H�����ޝ(���4�<�!-=���9�JD���ķ�}V��. �P�m
�r��U���=DS�����+�	9zR����(��=>�O���P��4���:��|�T�I &}Ϫ�7k�ўG�2����m���d~I.w
�زZr�]�"��/ᄏ'���?6��'y�!vp¿g��EC��x�!�c��5>��bL'ue��Е�cD*Axk�,�D�~�L��\qS,Q�TVcKO���x�9�����7]��N$�Q��0���N�� �TNMVD�pI㎻V�DF��)(�ތ4*c�������`���1�C�P�����q�E��:N��yMg4,��C���AnC������"WIk.餯=^�t�U=���<�oF��<����k�Q5o
5����Ba�
�"l�&��������8��m���h@�03`�6���TdyOCZUDS�-}o�.��D���8�	e0�s�"mq��Ք�m4a� �/�����06ObG��f_��謀����o�����*�`��4��k�8x�,3)�Y\滕i�4�gCt����L�h��_a5�ٔ���9#���~c����".u ��Hp�4�If��]lV��`\��ù��V=Y��o^���H�~ `�#���ϔ�j�p�ى�X@��pf�)�?N��aw��{-*�f����g������٠��ȋ}&�V^_i��(<��d^ÁF��u�$�̎8���,�<���E����;��Շ�;����Y����G�$��O����>��O��i4��!-��$�T���;]1�v�M��$Z	�Z��w�R	������Z/Ȗ�H��P����T���j���w��2_�v�gĨ ���F޶��>%B��3{g��>�s;�y��^�����A �8f����|&�rOW���| ��e"�돋	�C-
)0�9���@G{&V짺@��ϴ^��ZS�����1�Y̃U`��m5�Y��%��tL���%��)�Ivl�(F�M�v����s��3d{�u�|���q��X��/��R��ڌ����]�!'%ɂ��P	���za|��JC�R�k��6�>��2��R�������g�.�a���	E2v�9�NÇ�?їa5�
(�|���aK�L%�v���NK��Mv�$�-���;
��.�{M��$^$�a%Ż�طt:�k�������t�y'M��;Xv�N����/�L�4i��'�:���������g��^�v^�{,3D+��4���ߗ�\�!�G�[���C~��a�"e4�0����� "��K���z�}�s�CvP�P���r�R�L�X��50�)9>��E�LEc�2��b��1�wU՚�ZS��	�ϋa��Gv۱��爘Ca�ZQ�*�3�YC1N�l��7�
 �ԭ�6b��R�+M���# Qk�y휇��4v�4;Z9A�7�;�g�
�ɒ0��l�	���x�aW����Qԇ�dW˨_9�}8�7`:���]���NԔ�hp7��]z�f�����1�KD���lJzv�3��=�=࿭Dg�w�� a���cߚd�M��<W>��7��di�@������d)�@�?p������+�Q_y�˳:*4(8� ��yFNM��;y�� �i�=���X�r���F���gS��5���ܐ�S:��'R1�#���&W��׋����� Sŏ�2p�"&=��i��`������[��Qs�AK�ݦ_��Q�/G�f�@�L��窵5����iy��X��M�^-\�cI�D�2����vI�%�x��P��[䛉�d<W2��!�A��1}�5E1T��V6�̑˟9+��=ĳ���)w���h�n`�3˫ƶۊ6�S+�0����zR6%p�"jJᵌ��q��t	��\������^���?n�Βc�.z�	{ ��7���{�!���|�BPU����"��K�L-��"��O���DX��Ƙz	��D�D���Zk���S�m��7��\:�6:�V;Ot�]��� @W�qv>ϼ���I|�Ik"�l���1J�jY��&+�`��X5����Q��-�����sc�����A�
�����hTTq��m^�]��30%|b�$+��*� c��P7�|a�'�����bf�D�D�����D7-;���(A�I��^E���i�į��'l�~��+&�	;�cZx�Ɓ�k���Ǧ����t ��8' �J]ǵޑ�_R��[���_�$E?M}K���*�~�ճ5���}g�/���.����p�U����"��wj��@T�m�+Ou�O��O�B�vi��?��I�>2i����� !%��y�tP��(I�_��qCa�hi6�r+�w�w�]�b��"{�*?�Ԙ
Z����Z>J9�N����>�N�H��m��s݂��L[8�g��T�%�%�9�QNU�j)	k!h���u�e��-?0TK�<i�1��M�Y���p��9;l#�3� ��-�jv1d�ZT`�\G��ѿ�Lc���h��<ʝ�8�������Y�dm����>�
['���P�.����UVh�V�?�G���q����+ΛߌWa��e9�����:	
�-eznAѠ�������d"�����	~�pH�(�q=����iH���Q|!�hG��M�:��6�T���c:�܈�8֍��ٺN�5p�7��"/U�qbHB���H��{��R+�[J�9_{�����`�D95���+���OWW����_h��0��MY>l������%��3��&��Z��,�ޮa�&�p�l�Í�.2e��)㵁��`Q�G~�!=@A/ �����=��u:����iv_�+���.��js�⎿��Ik`C�~w0l��!3z�+�Ȍ;���!�8�J
���zRl�Lӏ�������4�hw�6[��Z���#�ܫѭ�TR�LY��#�u�H���H0�G���T�)F5�	�}��bt^#1����Vl'��Zs2t�^�x)�FZ��Rh��,�pSu�� �j), �!f����,�5�	ޠ�"�"��o"�^gC��x�T��~�|���B2�����(��:�o7��ڦVt9�F���x�7��ۂ�}�J� ا���	�Z��@![���eT�;)��m��9�T���BC�kSԡ^8]�۾�S�0����rZ���*t�Fna�e��[���&���9�.4�u�9��!T(��B��
:M�*��*��Cͩ�!�L�TѼ�K�j.3��p����2Mχ�y��,?�(�zp�9Wa�{�6��y�5��t6��NJ��t`��$6�_�Α!%{��{bP.Ĥ��f�:{�m������I���Cm� �9���L27��FG�,�Yq��ڋp&a��c�Vr����W�+����^4��&��S)`�'��<�g��_�ƦO�/��-����
�Cx�@3���R���N�����C$��y���Bd��hJ�h�4Z2}����G���P�y��6��wɴF�od��'��	O�=XO���b�!E�%(�����/�wc��!N<z����#ט6c�Nu+�_ �-�� ��=_=]�2��= ^�&���O��0JѪ�;3ݧ�ʷ����e|N M�[|�^�ѹD�Lz�*g��w��`���s!s� �Ǽ�3�wmu��p�P��.2:��Ꙭ�[D�O�&d1�٩O�Ň2/X3ۊ����(��v����֡\�΄�|:����r�������s�{��n����G��J��M�I�zp?V}���x�9�˪Y�#�����}ʁH�����A��,Hv�.�`ԫ�@��d �Gh9^���YC��&e|U���e�m˗��h;QJ�~l_n n�|��U�UM� ���$A�ql��y��O�ӟ��]ƖLfM������T�[Wg��E���`i��6����W�[�LuQ�ͷR�tCg�oYF�4��������dku0�4YM�q.ت��]zR���-k� ��$��V���َU���Hd�.(�f��Z,+ȵ�O5��3��?�%E)�U��x�3�%s;B��}�f��܀��}����|������	��;��u���X<�RV�%��IЭ~Z�Ck4H��D�A�ە"I��5_�+|	U��K^�@IUXl�fr[��r.���DK�O���e�2mb�+�ePZtᦣ4��x0/AY�`v�U�auP�{�l��'���]��n��S�����ُ�WFԻǷ�����:�1�*�8S{�'�i<,���az�9�J�� ��Y�{^_UZ��( �����b�%�5����0����a�31d���F����7Z�@�m�*��G
�M��[J���Ze�J�	����{�3��|�1�7��g��uq���d� F���,)���Bc��z#�[?��aAqM���ː��,Yq���#�
9�t�,m����N�H��Z1�N�0Z��r�!&�,�� é&��b)��&{U��ucN<6
�� ъo�P�0�.<E�%X�~�%�On��+��i�ω�'��L��ڡ�o��N���$:��
܈�߮�@Π0^Kv
����عs�u�j��i�Y��C�t�AN�Qʤ�J�,���SX�ރ��f�e7JY���M���W"P�nVbF&-�YE�B��"JK�6j��X�yX����\ֵ`�`�� ���˥M�����Z'�Zo��GbNHi�K7����H�O:�6z6��0]`9v��9���C�|�Hd��G�&�vC�c�Ji&�@"�">60�yK,ue���Y�w޲S_�Y�_HFl�n��:!�~��LK�I��ԛ/�㑩\A�Fe���;ؘ�=�4c�Yc
9��#Xk^��=��]Z�٪E�dz hP��+��o�/Ȱ����K
��pea������qf�NZ8I�Y�v�E:��g���c�ۋ�gX�o3
����os<�!�$����E�������@ƣVx�6Ǉ�q59敍A����q�g��)�o�?g/"���>���3�w��OTc�^�nū�%W�K	|��B��ͤ�����Q�����vsy��d&�0�ɛ����*�H(2���z]�\�1eD 0賿*�E�2_�	5̊�A�W��(.��r�۩/���C���$�8\R'r��w�����8)B�gA4X9s���&�n�����t���Z�-��5����k���'ċԵ&��m$;�rC"U+v�8���4>RE�/�#�mDLka�!�e�շzR�K�Z��?���O:>��a��橪O����JЩ]ŋ��d��wMt��V<�g��%�%~�4V��2�*>c!�V��7��Ηo���֟�N[8��fS͢
$É�~�L��OV
l��R�T�~���Jw(��^<��&od6&|�7��0���'M� wRY�q>��\�X(�+p�~T��\�Pj��<ǲ��@�&�l-P 4|��/A �%V���Ӳ��ޏl�9#wqJwZ&~O�D�Q>�2�w}ݮS�lon�׀+Z��(�ׄ���"(�?�X�j�6.�l�u�K�0�E:0(��2[���y�Z7�<�������u4�8'C�"��+KiX�]��_fm|��=�UZ_����zR�A1#�*_�'�]�S˺Y%��ٽ��ZW��� ��Lġv�ۦqG��I`�[�� A%x���h%k�>^&��S�͊��V)�brTo'�UR<���i7��!�p�
Z��pEZ�Ɉ�0��}-q�5;����Yb��?&��YuT"��2����3s�==ѱuc�Q>�9C���,Sb���#��^��A��������Ot*�W$:-�P�)�^�����{��rI<��� @pc��!I������f�lՐ��l�*������T��>Me�������ِۇ�.���C̬���V99��TM'��a"K�x9"��TmjMR���)��%���ˋ�C?��4���M-�'����`\��ʔ|� ��fۡ�&9kr�$�����?c��唥uR�Pd�����2��`v�ѥaa-��y�'�A8�����j����'2-���B�ż�[�Z�E��8S߬�΂��S����0ha��9�v���I�ó} �B"t(�`4C���M�Ix�����qI�k#� d-��&Yi�\��"���d���#�N�Oe�G^���<�/�k�P`�;H�Q��h��M�����a�U^�u=�Pc<��R�V	I���!�Mvֲ�m"��3M�|ɮgc��������ci���ßBa���w�6ҵ�7��_0�����ը�J���ۭ��^�	��D��C�rϷ�j�}G��I��ԉk���/'6iwVO5B3@�Bq��B��97���Ow�R�~�[\ mɀwg�)i�_�����Xv��c?5�7���w<h4���
�!��.}�\��^���� 4���G׿x�Kexd���ʼ�=$�3]e�������l����ϕ~��(�vZrO����E\Ý��.�e�,�T�M^��l|h�m�2.�m��5���8#\�׵���g� "��/�-��䨅{`���@g\�M���b<I��C�m���ݥ���y�n|�N��5��u����n�I��x�u8�A<O.��
J�.�0��p^v�!Y���� �P��q�?��RBB��Pj ^��������1��fb��T�����W ;�U�}H�ɏaj�/���	1%v����$v�4F�����E��Z
�j_x}g��t;�;�VԊ�o�Ab�@�c�䢼�i�h���L ��R������5f0Q�hQXw��%ܚ�7D��hNK���u6��<#8B���t����BQZk�#s�I���Y�[�V�l��6��X�^&���� I�28��,�H;ju�S��P��O�*����e��-2zW1�@c��N����/��칈G�(m���Y?�/Aq��^��	�1�����9�lC��lG�:y�у�D���S���Ai&��1��L/�x�]2u�d�|Q,�����J�Q^@���_	�v4���'�I��)beD�)��Q��tC]P�B&0M�}Q��)��كS �T��ap�ݪ�V>#��&�x�_/�b,&o	a�:��<�o��c3��DQ�Q5�w%����� Ǐ�C���H�X��ge�ĭ�\^H侼rw
��ʿ�/�_-c�s���	GE]���P�2���vŊM��wDR�^5��VvD��D���W�"�����"�p�t 9��Z1A��N�>��c0p{�Q?��tm�>�xTW��	[Ԟ�$$�J�lp��h��o@�R�f�L�ngɉE���9�-D0����O�?��ٻ'k�-{�0�����}��E�c�u.a�9��'��'�	j�24��� ~)m=�w?�}�Ft9�TYѬ��Z�I�Ñ��h�� ��Z"LB���c�&u�n������	�h�M׬0 �2�[��Y2Uf9C��_��*j�X3��uo����ԝ;{������vōP�RDێ__�7=�o��#J�IeG�J�����'����X赎\�-]�3 T��~��	!sQ�����%<]���&`�}zT��G�z���{@���&`���&�Y�n��t<�.]�.H��EuO�6�J�maN��7Av�M{\�d�4� ţJ;w�Z�s����B4EP��@ⱉA��RE�ȱ�J-2��ˢ�~�ն4�t:�BT<�������������U�:%F���
�����-�o�!|h;y齂�6Z����a]�eT�;6��|m':6�M<����
�;�`U�H����d\mK��u�o��bM��x���p&tGp�#7!���'ǥ����

�$��g���)���d����� d��?�a��U}�L�a 
Y��f�9k�,���� �Jl�(i�$�9�W��4S�rw�u�*�b[7e����]5��U� k���9)PɌe�"��|A3����_:/�P�@㏕ת�>����I��=݅�y&������EUQ�f�l��	9�f�s�����M����[]����M��X��P�^�����M)��G#�K쓷��9l=み�[4+k/أ9�uBs.ް]^����T��̀�;�?/ `���	��I�[��P�2�o�7F���_�&�+Ƚ}�}����4���@Ì�)y�3S��	����o��Ϛ���m�Br���h?}���'�xp�ź��I��Y��p&\'p�����t����a��׷%�8�M(n�-�.W^t��\�k�/��YF������7�{^x�ٖ>�&K�����E���E�ܶf�d���>j-xl��q��*�Z;��m�,VpL�J��dCN�R�Ec�Xvt� fݾ_����(ޟ)�b})qFzO�S�Qy�Z�(��P���LV=.�c��c�Z���#V 4FW�D(h���Dx�(�� #H�5ϻ�7' ��?�fj�*��5�-��o͵;&���Z�d�G*��4����8V�J��W��V��;v��8��l)Lnh��yù3ԗ���)C���:p���65�yt�q�*#&����"K�?�nB��6;;L:�2����-.�]ɤ�L�o�Y�+Z�YĨ������Mc��O�\t(~'60N6�ɨ�	�̔L=z·���T�Q�#�gs;٤K!MpPY0��Mo�Ǧ֎ٟSsV��H_�����^��ß��<�c�|��ƺ-du|������X�ℴ�#&$�0��Myh�w8�i[�����u�<���jb�9W�
��)�f���9��� ?wV�ٕ��ʒ��s�ǔD�o^ �;:����v9��O��kn�"Q䧴�'2��&(��5#�R<ͷ��UQRYx�gS�1^{���F�m>� "�)��}��~�f:{Y(�R�����s�
a�n�:F�2^wҗ�*�u�CX�&τ:|҆4ysZ� �LJ�/�P�{
r/{(݋a]~��6��D�9\�/E�A��� l2[HrG�����[t�C{������kS�j��Џr�/�Fˊ��V��#�>����W�	��r��O����[}�V�i\�hBS�AR+~2�a�A�!�k#�����N���[�
e���u	MtPPS�Yl)���|���'��/��-�|� a��?�2%цӕ��0��XL��͘:zY��U�L^B�k�m� k���ʤy��,�h�aɫڡGuW�pf�)#̇�F3b�\�Э�jY6����iQ� �T1^+���[��6�*� [�9Sg:*�n�C�I��4��t%)��7ԅ�9༶���G�sj '"&g�8�;���O$�f�Z������;�y~!*W�U�:2�[�Z[٠��~�W�vܯ���te�G_�7�j�>:�d�'�a��-��W��}������
�"ZE�a2X�=M��'�i�H�@�m�t�Z��Q����xbS�'����q	6��ϋ+����	�A���d�$)���-�-�Do��qw�V��G,���liN�� �I�������SfH5�=8UGF`˕�}p�.�9�s4t}�P2�p��O_6�p�6��4�t���^��}O��:�齔ǅÒ��Ξ���(��mC�ӏ��iN��?2 �vі+�l(�8�,��������!,�,V��H��B�q� Y�/����o����Ϧr��_����Qf��L�g���1:x��N<[n�����c�Z%��L|T�kf�o