��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�X,��W�қ�`Q4/�(g+�f��}j��u��2���Q�+Q�e���f���K�J���q�������u�¾��z;������:�ψV�zn@�޹����z�3*{�>g�$����<�e��9$!�qh�l��#��"��z̎?�C�G0�A�#7E�0����j��"�G1�u�	1>5Jm��3�b���W�?K �e�\~b��L�^E�Ābk]��l!���};t%�-%0�қ 8uTӣ���� �/��d����\�=���l)�Nʕ��/�ݴ�����d[֔��3��2b=�y�"��DM�L����;7��1��D���i	=�4�g�ܐY���c�v��8f�8�屚�&;��A�hჵ�Ȧ��daR1"T��T!�͍JB�kD\=+��kx���@-lZ�wؐ;	�x�Rov����AAr$U��ܞ��>`�B��.�{�s�$�u����LC��?������E]ȷe�� L��6�ƞW�~��K���in>z����_���V�?m{�,֚��%<�c_�w4�Z�8L��+Sfi-�,?�VL�nWB�o_>�T�X-�����?��0�<9:KC��oՏ����D�F��}S�O�h9[��ІR\Z%���/�P;ݶ -.C﫳���$��NH�����S�F��Xub/r�������w�G�w3J(��3�ڴn�����[q���o��GT(�E4��3�;$)�H �`~�ò���u����X��Dm��õ1�\3����& ?@n�L������2�{��a��/�.T�[�]'�G�0�LcZ���{�C�����L��ª�i�{Q�5���UtYR��
�`o ����T7�"�c���@��b��wlz�9��}� $���y�A����Dt��TN���@�Ճ79^��r^w�hQC��
���5#Q����3R|���Ȉ����'���\�0.���2%UVsnw4e%�6���(}�d��%�:��V�{�|L�@�x$�$Aq{�\RQ�m�e���՚���	��m��>MI�/ރ��La��!]�!�����$<	�s'�k"f��������gKA�z���K����ƶB�/a����;3���Ơv4�"ژ������L���5s¹z�]��MV��~�o����k��R�h�M�������L! ��%����<�sg���� ]��^��_�wE~4@�,�U�!:p����m֬T\ȉ���͠B��U�I�'mx��U4E�Z��l*�@���^F��j�h��Z�[$��p�5�[B���,�����s$c���[>)F�y�"UԪwI���W�W��C���g2�y!b��GņN����9��A�L�ٻ$���_=Q� w�����a^w�+�z��<��ٶBLz(ˌ 4V��ʻ��`�ekӞY�+�C��O��Y�/)���u��4ŧ-=u��+_P���)�Uha%q���EL�^��l�+h	��b�@��u��8i�3$"j\��cMsMYP�~7U�tsK��C(�����~���p�f�N�f�(�-�I N����D�Q_2���CZi����@��2�HǲM�#C|�Ű�>_�*h��~����K0�=�~��I��B&��L�ȥ�(�J� C��t�EP:L�'�l���rȵ�����9c���]�֓F�$H�9��_DA{�r�e��G�����jrQTWDw`�v!�Qj�_`ߵ�Rz���)�X�*V6c�k~�z[弬�Nֈ�1M�AoR�ܨ1$�����檪��Mnl����XU�oBQh^-���H�J-Z8_u�@<$��7�t����Ad�o��6>��ay���sD*Ie�	��Ǎ7I+v?��po��G��6��`J*�	pTd�a^h�D^����3R�CK���qwK���˻
*��%��ļ+����&�W���P�QxHy`�s s���H�wY���^�Z뺽�8/p��F6y�Î�!�2.:+e�Jŉ���������P*'���ͳ����#hc(�p1T�o��At���a0���{|���d�M��BJyr«s��{��V��)��T��^�c<�p����6�����r�c�����9��fi��\��i�@���:YsT7�Oi�������[aԢa�u��av�'w`����V�/ɬ䎥��H��=gĸ[R��.m�n/O�\>T΍���1���M�Iw�޹�b�x6
�z��lS��B��}-�Mn脜V3���ݝ*��tu"��SY���*��qA�Z�-	�G��M����f �����yaO��Q�ڀ��gv��]����I�|.B�P�5!EHn�U؎n2fB\�ԫ�`	���H����&2�s�%#j���O<�冲�3L��h�A����ګ*Dd�}���!��ʮ���������7���k�9.��(���
���Q/�+�,��%�a���81�|����<��@�.
6�jl)�͚��,�r-!=�׿ݡG��k��b�O{v�֋�|�j���b	���[H	w֞>7#��H[S�Woe����H�V}"�8J]��7\	6@�X��֮�C���v�zh\�D+	���yH�]����^�P��Uun�\>�Px���/�uZ��j4���z���]�>vn]X��C"Nb��`V[���+A"�,@�	!7�2�m/J�lT]����H�G:�dǷ��~�ʗ�� �hR"��JҲ�R��1!��9��7�F�:��^��Ju�+Rg8S���H����N����N�:-n�D.�Z�͂�cCHRklQ�xn����1	�-}��n��w�h�ps�#l���H��Z�����m�uH���I=�`����wzPC�a�`ͽ������]�F{��/�]�h�Y������Bob���\ز���675���F���R�١ۺ<�h�,�k�1�&��nK`�W�
d��*��G�SND�z��G�B�3*��&<��pɜ���1\/)��>ۤ�澺�;�<o*�q�ۛ'{�d� �Q�i��^�� 8a�iu�� o�_#�g��.�G��f���@���(�N�)3�V�����t���Ja�f+�~�ҳf�Z燒�0�����!~��7��?w�c�����e�H1�n�n@�}�.�cڳ�nG�܈�F��$��wU#1�caZ�W2 �"�+y�&��w��|4�rS����R�[*�k)�/�{CA�U���^&��UӁ���$6�,�V��/��&lI�4��c��]���E�<EdR*L9�+)5���,v*�/33���M*���G�ơ�ȻkuiA�0�ծ���-)��	w��x�El2��P�7+�y���q
~ZN����<�b��EG�u"9�J6δ`�g�h���D�t��E΋͖쑯= �`�"u"�,�ӚZ,�ċ~oH#mp��l���2���Z`R� 	�� <ܮ�4M���K���f:�dEE��n���#t��8�.)�)hU ���Yŝ
ʝ�߾��8�w���7bt-�دc5Oe�;�S��:�R[��ʁCus��������s�8�qT��)��=�iD���Uj�fz�1t7ȳ�7�����6��TV���㘝~�ޖ8{������:��.
N��:G���Y��A ��J�a���.t�������ʙ��$�(\�dX$���ηD͙_�B�sتYĜ�q��{�7A����Y�����Y�消�9���靗��S"��7�**�C�gV��W���BP�,ԺX���Iy4?�n��hq�C@���@SK-PYI'����8�f��`B����R���X�����Q� 7��d�������|������'č]	��y$�!��a�`�x��'Ў�w�ߍ�󥍇�(B��j0�p�A�e��/�Z�3�m�8�u����e�Tyˠ�-3���n��M.�h�<>wS�e<��P\i�>T��q����Z]:/}��Ħ������:�����z��(ueh//h�GG�@����I%��怿'8m�I�^�n@���ו�Es[tK��[
��S��x���s1;�#ӏ�?�Îj:��A����5� M� �kVRpͭ�o����ZhԀ�2��@!�&���#�G��2p��l-1AL��Mc"7��e�P���]�Ak��ɞ"A%��L������!���aK��(؂D"bE{�w�&X�˩'�_`���V�;_��vMaJC�	�t����-������t[��Sw�:A�|z��M��#��C�@"�f�A<�XRG�f:�p�H����R���.4x�Pd�����p�A_�HRtӑ��eVB9�$�뇼��*ʘ���H����m����t�CR��UÌE�(i�Nkx�|�N8d�0����iO�4T�6�6��D�C�3Tv��"ycV2��<h�6��]��?�x��P�R�E��Ci���[ͷ�ժ�ҟ��������`o�C���8�����ER���x�e�Ĉ�D����l|���^t�{[����t.��a�Q�Ċ>^n����.��8������r����z�TKi^�"��e"MsL�(�:
{F˦��� U��E&�8%��X�Н��}�1�GV�0����i�6��]�K1��
���X�2��5���-cP����#���b����x�}y�P�K��`�e���6Q�Wɾ>�Y��e����i�e���Os�  V8�C4Z�ns���B�ײ��9<�-S���01�9��B,�kH� �-I�2/=G;�$lQ#cѦ4��$��H�F��?���ɤ4�7��Mi���\�SJ�ã�/�1���HO�"�^����@U���񖉵���̕�%	�w�Ϯi"��)�
�n�ҳKZ����w��..�-�=�B.����V�`	{�=w�0�cwӪ�cWNy�<��������>��S�	
0X�|g��5`�����x>���&i���[�$�g魳��k�	�@�Z5�����V���G���̊�0|��K�3���KH�}�1�G �@XZP
��Y�ې	�̱��Y
���5�Zd�o!A�Cvt�_x3�<	�V�|�?�[H�Ao�����MΠ��ϵso�y�Y�K-[�eS�ֈ����}����|E