��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ02R]n��Jr� �/�+�8�G�;W������7iHq�D��'�K��u>�8$���Y��	�w�#�t!o|V����ev�^'�O��a���8=�B�Y3�<��s��Tr>q	��=��)�s��.�N�]9�4BZ�4Ç��MFk�I�#-��e����/jϪͰ`e�����(��h��0��z�$�w����b��\ٮ�S�^�#�7ӈJ.]���<w� �����p�11)�k�����b56�2S��<��-���.c錀���R�5�la|�.Y��Ts�v��G%F��H�v��W�O����\�8��ٌϛEx�h4u�htLFh�W����N�&f�+ǯJ�����y�M+��B�؅u<�4�-�Ѿ�}��o[e,�s�l�)�������mY���fU���׌�J��S Y+�#f�[U�d�

��٪�A�]�
c���� q-���H������ǡ ��+�9��~�]*���������8�q!|1��Kh���@��T]M�ԖJ�?Z@��<��\�R���
s�x�a�y\�\1��ƾ�?��E"�ж[������t�E�Ɲd)0��|+�.��y���7���I�lEu��#O�_f�F��{�9��ʂ%��EeXB>Dr��OO��&�D}�:^I��;V{���	���S��mo��:*JuU�	@��f����-S�^
���!"���pQ�c��hA���������x=5�o�����?	�Grl8��"/E�4m9��l�������Il8bME(�@fz̠UZou(��	�`��LWn��������~�?R		6Vj��Nx!��I�,@5�3c��� � ��K���=M��� �(�1��������lW���D`y�T������+U~�t'��	m��h��Te.���{��"ԧ�dQ�ﺕJSe�vS���xg��x�9�|lƵ[����uU�\�p�$t�V8_J�C�na��yiD�!�F(��{W������5��b<�,���@M!
t�O�`�u��]�	r[�
t�g��oQ|�d5��P���O���C~���xlX��t�HAg.��J�# �~�zh��:�]��J�?���طUq1��'BX3�y8ڢ��_�!�)�w��=��(O�����6��i��טT��B
`r�����������D�0�.(P!ROCv��#��:��QG�IyDNJ�yS��PV���N`����-2��|ٍ�T�*����h�j~�?~����Z��2*��0>>���<N���"�e��;���[�k��͘)�-l*��o�$���Z��#;�� *1��Im�#����j�(�Pe�5�]=�l��H�
Iy�@n���}���;����J���0��ȱ:�j��Yq	ew�Q�Hj�� 	�
�8kj-�����@��"/��Fp~!�y� "�y�qS4��Dޟ�����q���&{�ܩ{�����!�@4���U�RV �v�S�9)�7��&jA;|�����S!��i4����Kͥ�)!I���B���(� �pם\&�M�����(۲�*���}~L:�����L>�� �݁2߷[+.b)��O�c,�Wd��-�LG���	��B�:�b:��>j|CD~�[e�{6�#//�>����s���C��
*8�,cha�p���H5f��.�����l�P�����G�仾��o��U}Zr�F�N�qVv��:���g_�{�hJl/¤�rL��+��`�Q�ЛYY :��]^�L���ׇ"y5�mM�Q-��PLyN}>E�x�/e�83z:���ڙN;�}�T�����1�bp{�>��r���eٯ���˄�d/^�(�6ِ�]1[�_����m�.�=,�/��)�&�yh��mL%�߅aO�ۥ	Tw/d�\x���J��%A���,��zl���ܤcjM�͙�p�5�K����~���O3�̖���&篈�=�)�����u���2�i�2��뼛q�x�����&淏�;Kum��u��� �Eu���玭�"��#:�x�ȫ�/	�{ʐ��<��eq�Ak��:
B��wr#	��*d����О�(��Cy�̌'|Om�C?ݮ^�������A�6�M�w&��672������Gc!������'�~��C=F3�-������k��w	�!K���3�����q��l\m�|	���8�� mdMRC*�'��E�z�D��~���=;`S�
�����q�b?"ac��a9�F�F��7`l�l�;W�� ��FN���޸\.j,	5B��Y�VG�;���a�굫ƻ��`��˹���8I��ڣ(�
��`)���N����wf*jI�e���6�{
i�0��t�&�H�̐���}|$2��ڷ[?�7D��L�(�Հ�X��zQQT{�/�[F�١lzj�8��ҁ��ϳ�kc���&����2Ž�Yk-2%A:~�9.��t���Zt�[�,��!��5��� ��f˄+��c�b�%$.���JE�t [�q
�,�;��p8�=1�u8E#�A��^Y����@��T�
��X�""I�{�0��8��oE#�4�
��n�8�~�	|��L�Hz��K�RX��@G��7��.V�ls�yd���-.u�T���[I�+Ӏ��-~gA���X�<
���J�(�W$�oZ٤�'t����&��䒇� ��5/[�܂`�V)V;(]�L���F���oF�N}�N��]	�{Ϧ�J:yr�)	T{���0�+ƴk��aG�yvZzX8��,Nڰ+ZC����u,f1������0�a?s�==6}`��հ��u��1'�{��T3�s�ޓ��E��*�����	�-L��~����X�@V�6�lo�#1�!㽁�_Q"�QfI�I�po����a#z��b�^�ye�PI#��D�X�����Lc�}�%������M��:43��+Pʕ*��Pʘ0���<���434��m��O����w���HMn��wZ-@B�Ӎ8�@Vo���hu���ͱ�.u��)��"��c��O��t��I�N"cV�\�u���J�-��u<�}A�s�_Y[�^zZ���;���Nc����>!,b�L��u�	�N