��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ/F��	�zVQ�6���g���3���i6����N���j6һ���j�>.|�|�g�eb�.U3fu�）8���vJ8�����ś�@9V��*nh_P�D�*z]��;�<�k4 1,���ԕ�����+���]3�X�D�O��H��y��?�"f\�jh����E���0�Fc�n9'����-?�]5�AoΛe�rHW��u��l�q�YaZN��)6�߽n�[L��4�cT��%W�dg���X[�ę���i���P5�6�Aݵd��1�?�}b���^du�T���?M�`���ڈ���w�_����l�$ujɦ7���h�@�1e�" ݂�B��~�j�����p$R+#ʀ�3��J�Q�F�Y=�hR��倬I��rb�>%e��AabwRⓌ�v�ie�u���x.C�M���m�f���0(�n{W玲š�"�Qۊ����˗U��!0i+T�`cM�t^�P�2=�љ��'�%X8�w��c��#ڢ!:�@�=�I�Uu�J�IP��I�~?�V�/����SΜ霟��Tv7�b`��	0��ێ܋�FK;`\$��llӽZ1w2![XCǒ{S0b��)�^&�w%rG�K�����s��X�&z:E`6����<�Z�8R?�D�
�;y7˫`����)�4���R��:%;_��^ӠYh����2�
���hC��P�fk���)@�\r�����N�V(��JNxV�eg+��~���z�V�O
����x�����`%�2��*`��tn���`�o"*�uCy�e�vơo��Z'I2˓|�����B��T2�1nA
�.+�qS�"���HYN�NƤ�G��x��!�9�������ffp��1�7� -����M��%Y|z ��
���%L��Gz�f���+�M<���3��Bhb��=s��6�H���</c�W�x:F(���E�%������0}�v3'@nY���Ҽ3�%�F��G.�$׭��i�49��E���J��Q>�d�ō�/y�j���7���l�&��|y;c��i悠@���yDNg��..c�;v�)��r�4xu\W�jF"[���*�=�扊�����<ٰ|F���{=}��O�&���
�����M��J���_�w��E��1�GkZh2��KMص��6��Za
Ҳw%�)Tip��m�a��74�5�R�T,��R�|���
���O�bM��1D���'�Xh��,�w)�3�.����Ϧ WWmc55���������Q��u_[���Ukx<��*
97�X���YӉ/b7<�ɶ+�]u2t���M�e�أ1�� ����[{�� �q�<��O!d�?�Raъh�
�`2�H(�%���vtAY��nU���Đg¿7A}�rĕ�2
E��=0;ze�y�z�>:�ͭ�#c������
�=ln$"DheM{�ɔ�9�B�if�8ܥ���P|����'6�`?M�!{RT3D�I��8 �hnvm����#M]0]eo�/�}J�/e$sگ>���zg�#��xs���\i�A,�W��%��V��������������;�wuV��m<��?��^�C��7��U#i������>������[�i�0����5U�O8���l�H�$���(������^�K��w�]���6P����{���Ʉ4d7�y�:i�5�'�Z4�wqr	��^��7J{��~Z7����1*�)�`���Ƣ��&�V���*;9ܓRo{9�����jY�\��k2gp�cU�	E���TÛ�+�>�l�߼AD�|�:��-��e1�8z�s��z���*��0=(U��s�p�{�Vl��a�W!l��ɏ��I%p]t�m�C����;��TWrt�C�V>:�O��>�9�|�54�5�\��+!�~DJ(ǕJt1*!���GiP��14!j�����Fڽ������TČ�/�K�v�g�pľ����aɝ���{�� �7R=L	gX�(�[7z�3#AT�T���f�;͐�D�%�U�w��w߯i�`y/���ߺ}�q:
�)�l����|�L��Ai<p�{�M	��T����;�U�|+3`Ȧ}�q�eQNn�i�y�Q��0�.e�e�\���$x$+�6��K�;TX��T�b�̐��;D�.>+��#~P7r�d&���=��z�;N3���Ia݃OHuj��ng�qYg�mh�<Wb$tY��ѱ"�۴\:���@vE~]7�b��O���ퟫ�A��Z{������賹��y�ROV�p/�������y$�U�'T�ᓨ�$���ѐ�j��O2�_ۂ�Yܖ�vmR&���6ǉ������Ĺ�Z��.����D}<���ܟ%��y���q�����[���(�B�nlC+!0k	��¯u�}��wN%*5�ȓ�Ϲ�,$�C�K+`�C�xW��/Vw�n��ha*U*}E���P�)�e���R�Xnn%۔��%2'�uv�w�<�i�͑��w�Vt``"����'*6ټ�=���XX�Wq���6�,�TdpP����F��o�ƭ;o.�ٸ1��"� C���G�;$���*g�C�@sie{��xx1�I�m|��1j���\6��R�kL��(w*�q�ny��$�y3hF��ˋ],���/QG}��v��;w� )bR�m�bb��}����R��"��؍0%F��Q���U�(B�7�kRs�<���h�ٛi�3�D*��$쇘��YC[��e�)��+���1�e�Cm�� z����r�=�����
7̵% �;�L��ׇ���FGO�J�{Ag��q2-�`R�� (�o��H�}]G��
��O��I#Ǐ�q��"_��9����I�؋����Q������ɽ���z_��l�*�C �0����Ygx�l��<����_W=����}D�
 &��d��ξ0�;�|�����`�ØOx���y�U(BeM�ZxɅ�\��ꔔh�ȵ8�>���0��gl�1��T�E$��,R&_E*$&��L�-�/�5DK�Q5q"����_�RFu8w��w(�4� |hft�\s����觱�a���W>�ӑ� L����������������W�������[��s,���6K&g]g?')_���D����!�N�ă|TH8c���b�h�j?R�'�e�7.�P�̺a��������.$Ǩ�	�h�:Zs�k�OL
��[L����`���S�S�i�A��4N�N����ҏ�z�HD�FN~�	����L����)��C�xcPGX������2�U��������E>8�p�}�]PV��+�Q`��3�;��m���T���(�������K��X�r�,G��x<���Z�t+|��������F�T�����j��(#Ex���1r62��}&
�2���dH|�>(�Ƨes����~���7\ّo)����{��Τ�;���U䕓c=h���_��E� �~&�!"(a�q_Å�,w޻�[�HP�}G7JM�j2W�2g�j�U:Q3����A}��$�a��Hn�2]�=b�Q���+�g��6����JBf��q�:$U�B���.��ȋ�q"A��Q鐽�G	)���Ʒ�LWשz�>�|�p+��7B��7X�f(q+m9�?t�N�E�5sN�WR����4�b��5[aDG5.�[Kޞ�+f��B�5�dG�~u�~N�7�9��PlO �sYá̧az��E�9Zi�농�s���
k�b�d���ʛ��Rȡ7�E� 0��YDO��cx�V�v��w��������M���¹���Z��:��i���5���K��x�3383g�d�-V �4f'�������N+6��_��vw����C1@�mhh�x�:�jk��h���Ol�<������3���S&�,D��f|U�����b���|�d�5�M�����Ebw��1,�A��_��H�5A�iVYֆi�$p"� �� VIGG�{o1~eBȣ��#�fe�jR줩j|��*-�̵�ȅ,����,QX}s�6V��o��HAMp����'n?���.,�v^��D�FS��1>� 3�!?^v
/�qD��Y�:8q�W�jH?�:�eJ���o
u'�D#�jg��"R>�lT%�Az��)�duD6!��=U���e_)�ղ�+ ���"�oo�����K�u�����1�!v�����IJ�VIs�c�����~#%��U�'&� oI��s�۵���y"���o7��f�@=���ߔ� s\Wl��..,�u�G�ݙ�������c�/�=���wL�E��XT�i���U�����>�Pxi�TϢ����Ė�C�M��FBV]�`B��jv�paCD��sq�*%�ނ��#=��9��k7P֡�n��`��<�j<O��V����uE�ӹ��E��:*�^���N�dJ��?�0��[����8	����S,I���Z	�2w��H��ϛ
�.�zSoh�.�'���E��u�KE1�O�T`H[�p�m����A�!aGXiT�U(������@�ۻi�VY)�%�Z���&�Tt:�cQ=�?�MeHy�x�P^H��_�U@%NH�:�*���Ϟ1��J�-=���i2���)&�}S�?�]ӑ�Jj!T�J�r����z��_2��~���J�8�+��Rq���&�V��@ؓ�俞�B�����(�.������AAgȈbz�&e9i�K�W�wn�>[�:� �!z|��H�h�ۈ~.�w��ч��ŻO���9uȉ� ���QS����nPl�PEI_��s�jc[oU��O,�޸�K��bCR��C�>喸?�][�;1�Cq����_�W.�U7ymA.���s�I�nE1�A�~�f?�S�Xz���F$N|�. �'G��;�!�X����D��"xO͑ .�雬-J8[>}]X�!dY�w��n����8������
XZ�[ᜨK4�#�"��{zA�lW�@��O��D�����U{��O��/��M�Y/���"�`�k���{b�TR��?�Vo}�f�����yV㚨���af��&tԩ�)%��l�2��]�{��hq%c&�ؾ��?`%�.3�J;���u�Q�`�L1w�O�J,�e�|���^?��+�������jǌg1u�jC?Zh����,����%|���ԹY�/� ����Gm�
*ŗ�܃+O=D�K�����)�]����b ���3�8��dޚ��mix�Ou�Ae)=!�Ù������ȱ����`�Dnu�����`���6�\0�����$Ly<W�NE���fC��L�2��]$��\�5\�h*�}�m����J���ݏ�2Ύ/��o���X>�W ���`S�&R�`�"䱱���NC׌�c���<,�?I�L�v&�����E��2_��\��^��%J��`�>?���Y9Z���-�h��td<��1����(���R.B�ʍ��#IZIi,[lm�㺿e�D�1��oAĶ5;�A�@�k?����8^���������o���.eE�^�;b�����7�v��)2~��5��I�V��98���s�u�5i���r�s@}J;���U���,�S�^]�d���W���:`�Bo&��_�h���~?Y�fdયFp�R�1������3e�{>ȑ��k,u��B~S2z#a��	$qU�敷��E��?�m��t��&;�Ӟܕ��_F���|_������96�O�6;.�Kw��4�/���Xņ
���_��Z��6�}��� !��d���]t�]����7l�j��Dͬ5|Y��:����͜�ɰP�(a�R�ee�\ؑ��^&,~��7���_	����16.���~w��w������ /#��w]i��I�����'ء������wϺZwc�HƱ��4D!�,�^ɋ7oȉ)F*L��>C]�X���� Fq�j�r?��_i~q��,�[M$Dr�)�Ĵ�^0���g����݆� ��|áA|Cd@�:�w�|��y
�u�Uo!�����Y���Z�mQ�v� &��f�k��j4�P2K�� a�k��:�,����X�	���
n�x��2�%,��k�#0BN��a�bN�y�gFj?��Zj����p(��ok��!����6ٸ~6oV���>�ء]���q����q��.`j�����YU�^T1��Lh�&���R��8Hww��x��إ3� Q���X��C\�j����W����5��ݧM���k2ӅU�i�e,��B�T88$�ߒn��B�~>c�1:�P��D�DC�YV:N�~&��f�����r�D�M7:�f��->�c*��U ��Tg���ƷfL�B�<l�05ᇬ焉F���r�^�BBu<��[r��^$8d�T����'�	�1'uX�a��?�gq[(Aۑ�\���!I�]KE��H�!�����z�Qy��jQ�����br�`�S�ҿ쳀5!�Jv:��I�[FE�Dp�]�;r���=��F�K2��~h*�,7#��W���y1�c�)�C-Q�üp���*=����ԕ>�Ĩ
��|�7�������j�k8��zW�pK���{K=in��4F	���ó�O�}��od-�N\"M�f-��w ���s؏�+�v�D��ѿT6'D���x�aJ�w`	z������#��ȱ	�����֨h�����F��0�MRu�|�~�j��|2��J�Dp��|�K��-�[Xo*c׊5�i��[��F�-���U:��B׬�����/��T�!\�_��^g�ב a!��{���o8���{θ�,��j�G^ɒ�*���2xf���MϺj�w^�q���C�oMS�S�Ch�v�IG�SX�VBqv��dh���B�~�k�{��܆��b48���w
��O?���t����r!B3�B�1d�?F��ބN�0�c���z�@$p	��^Z�COζv�Z�>g�T�sm��-Dn�#�u#���)8A�lm��ka�N�8���jE\��@q��d<��cĺ�1������E�Mz5V_����Čs^�FN��/#��=��W�z�׳�>���!��ܿ���o\�Y2�#%&y�)���5@V*���d��D�]��f����$T�^��` "�J��į�ag`���3���)h���/ij���O.�� C�)=9�P�O�ig+)`���HE'���׮6�Ke�/���ٽ��8�E)�Q�j�=���*�%h۾kw�m�Քoh�8|�M���!��G���6,+6T��ҏל�U�7��,j1��)=p^V�N�>�~���X/���2!�]�5N��a��yOyC�#TԈ���+O���w�Ke?��g&њ���,����QP�98�� oA����
�Ʉ�����Z�GeIW0U�����"�R��f��=)����8����Zl0��0��3!��,/���٫��LO  �X��[+�l�95}'�B����Z�����r8R����o|;�`�h{�o�!�L��Ӕ~�|Yᦂ�ⲯ���ۤ�7x&CB��#��ʝ��h����$򷢃�	4 �}�2�4F9M.�A�uc��GA%�x�o4�(S�a�� l��=�I'�>�O[W�^~R�ڼW���$fE��S�*��?>�0C��B���L�6	K\H�l%h9���t3�ΦO���'�J	�+���8��������=���b���*�DC@L��L��u	4FA5�Y�P��.b�	����.�`z��wd��qS�RC�L���"�{](��NP;"��X|�:� ܺ�e���V��ø��u��G.�D!~�[��Ȱ���:C�B6�S��q%U�}��emH'@C��>�=A=~�V"/�r�\Jᑭ�
�%��%��3��'�����8Ti�$��0`��h���L���>�h�jf����FA��9����������'~(����3������a�ń�`AP��y��>��c��+կ�)�}�A��,#�b��~
�`Dd�#��n�iېS]�a���aዋ�h4����X���4��~Q����3$Bv�����>#����ERB��E8;�l�#��R���qb�f�-�r�*�c#�|�b�@W·N����c��R���ޚ�@L��o �VK ��>j^i%7�>��;[ld��3Un�<��h��F*�T�4�]��o�m/�4`^z�k<�|��I98�89E����u���,�C_"A���X������}�ˣ�[?�юS�$}�3ms��:|��P��q�,2��@�[>����|ee_�������j¦G2����$i������$6�=��du"Q�%�1NEr�:�D��}������H����p,M�5%L�?�iWў�z3c�ȎT��v &Y3��k�[n	SL;E�u"�oW�a�Nć<@�z骣@�GM3��}���{9�इQ�5˸B���H3m�g�R`B=�ْ�}c�i�AdnT2����`�V�M=�m���	��>�f״���x�JR���� �r��oN�Ui�S7��8�X��;�!��}����k���*8�+�	 �@��ԘH��*Q�D����s0�N������W��G��T(��+��Ke�E�Zs�y�F��qINa]
Y�v��xi��lWu��
�%�1�]ӷU�'��z�i�q��)�u��ve���AD�k���g�� �_'^�u"	��nSh�#\[��q�3��74�8�gQ<Y�Y���Pl牖��~��l�YT�Cb�A�p�gN��z�w*��1���n1P��'_y/�1q�!��Cp��C	�c�Qa��L��`!�Ű�,�%{n�@����% o�w!�,
�X�G"�YƐ%f���趍\�.v��p�>3T��u�Y���ĝ��*E&x(Ge������6^D�f����O���M��
����84k��9$�:ZW���r� �R�&�����axv��{H�з%�ؽ���N�X5� ��?v��-�->�<�&"�q��ͪ8&y��٫��N�H�@B���L<0_#�KGC\L��;��<�	���]�6ᦰT�K&Ҁ����T-���ޡ�{�Bt��|.+�m��n�����IY��;����r�1PR���[�FB������0=�8��		��0���jVh	.�n�	t�t��rKcJJ�f�!)�kH���-}W)T��w�����eT����	�Ǥtw'=�NW|�9������Ȟq&��?�:;�.u��JsM�J���iI��)�Őވ��Q�(j{ue�vw7B��$��ҍ��,s%3�]����{$q�mVeA�w�8���\ఛ�/Ł�K+g,w��W�f���ʾS��D�0�f��ʣ�?�����3h���T�_c�Ќ��KzpZ>fn�2��$��BG麣C
����1G�������<�;UZ��('���"+o��}ga��&�%{���$c�6�L�X�6�����+�_�۟u�%�`F���k0����#U�ֈH-h1��	9�-�2lJ�����'i��/%*�T�D�]<9*�8��i�ʤ�� �`�ĬV*���w:�F�O�����,PR��<T�nDj�R�dcp�C`J�T�-]��R�>��ҕ�DH�T{G�ԟ��+��-,Lx8�p�����6�%FH/���B�`ŏP+=W��Z��6��q;��\c�S�t�u]5���}�B���vMRb �/JV�%��5Ã���Q���\��)e����Sq�_p�S?�~�>�qe<�@``��Vn��H4%mKpǈl�%{�-��N��Y����a�����ӓq�+CA�]5"���r�d�����|�%i���",��]�3�b7�mp E�ΎJ��ޗ�3��?F�s�(�z�DH�&��H��vJFʧ
dk��ޖ�=�~;H�5�!��^��y)��U�G��������h��0�p���j"��o���++� ���_��;� � ��Լc�Lk�#XOt���Q"f�k�i� �Ҵ��ϗ�u��膈�C;�t߱O��Rr���&@�J2L�eɕ^	e^�1l:����`W�J`63Dgp9Ym���GZ3fp��`Y�	��w��i�R��/���p�
륖�x%��A�ɺ�E	7��Tȏ��P�g.v���@ :�����l+�ͅ��<*f�:��v.1Z�leQ�D��ȕyO�Q��"@/k�����.|�$l�2�7A�c1�XTA�'؎�"8�l� �{r7�����<ٽJ��+F��_��Ta'c�+S�J�G�
Û+R�eM���#YW���3��z����nC�l�H�R������|�"�'3��{-/D���C1{t{nNь��K$*eM9�\#W�)Q
U/pw�����3,��_��X��W�틻�/��y�?����R�@�w������N�U.`�9�̰��<qd�����P��(Ӹ�/\J=������������_�0"�82�d ����MD.r^P{c\L��-�j�;?q���'n��7�X3=El���
��W+G�#Ob-��÷�r��fFw69�{��*��6Z�Pe[���͑��Oį�Q��� (� )~:��i��+U����;���9<���*%�3���i_�
`�l�I�-(!���/M���I*�����ao�y��s<�M��4����C�zſ1�S�͢<$���ۿl�0el�H�	A�#ɿ���� {���:u�[S��'Ȟء\�e�
e�� l=eC�6����y���۞�KU�E?""Jrr��OR]\�P���m�\5V ���nI5N!��\Bx�n7� K��W휀��H�P���R�&�P�nk���D�ot�6|jQ�tU�>[x�����[����� �i#mP�H�3)��.Pʓ��L&CY^�o�2�]z-Pϒج�u��N�!!��^b�q�b;��7��aކ8|C�P&�|C�Y!��2�u�}��"�ʿ9A<̱[�y]/N�	�7�b&=4��)h[D�Cf�c�Ѡ����x���L������s&]׺5�	��O3�X��Y��8܇���G96;�����NT�*�]
�e�i�\�_�[�}���e��g\�?z%5�O�4D��"��V�v|9*rk��}Dgp:�?���*V�h^�"����J�������:S$���^��w���C�Z�U�L���_;9���J�Fa[5�{��]���7]�5�����ش��ZMo���VQ)�Za�g�,;�BoWDk��ܯ��U�yXV^�j}4��Z��ں|	�$����۲AyY�X�ީ�Gm\��/��(i�&�����S��x�Vfp�SW���(���� ���Y�d�����~իG_�'�R.�V�J5�i�V	ϔh]-�'2��5�:N|qo�o�4�iA~s��,�l�R(Ψ�b��]KE����y�̂qQ������)�{%{�eNˠ }T�T�
�4k�� wf��l�c�+��#�d7e���M3J:�����!!�(�2ӡL��^9ݶ8��W�ilL�
�`��|�U/{�\5���&uĭ�,6��j�B�Vq0)�{�Փ.����@��3���i�)� 򬣈�[����A��3H�&'ĉD�ϸiR�^��
�^��s=�j;2�(�LP�;��jo�ͼ#�H�j��L����j���	�c�C��Em?�.V+�pO��/�R��ܰ!�߷@��D�r��s58���7��yOk;c.?a�b�e��:�p��&���Ь+ 9����j`���aU[8������2l���Z���+q!\��E�2��w�+2�+�"B�xC�Ș���Xw��W���5�[�":R�R��~2�sx��\���h�!`����1���ϗu����Q�|�"r�w�}�����GӍ38���	�}�M���YG����Ky�>,����������`)����ǎT�q�|s�hg,^��V��6�o'h���m��6&�u�`�iɯ}+q咥�L[aO���,vj�
�Wzœ��Fp�ј+�vEl	�;#�i��$B���]ل7+Ê�Lɺ���l�k�4�2�章�G�Fx��vYy1�uz6�c���ǅM,4�爲�֚�8RW�C;E��}���&���<t-�ê0�8\S�&��Y�Y��R�~��X6@ݴff:�<j�Ǧl�ɍ\`Տtq8�����e��,��C�W������s�[0
�U��6uAċє���8YI�(F�1b���"wE1��κ[�%�cE��\T��
���{"�.���<<�zK���K�ַ�֞�a�N�n-������k�С��H�"�6܈j��]tD6]�`���PcPB��t�?�e�t���4И��L�	�ŲQ2b_}g��h�d�^i7EΙ�N��j�![�}+vz���5��D$kF�H7�}�UoLd����e���O�����rJ��K�|Vwk�LY4��f�p���,̾����+(X��n�uV���{+��57)z�%����K�X�g`7
�Ҭ<Tx;">-���ί/��k� %\�jd����U-y��i�&��dq�/�b��V8 �r5bcwc�1�:�B�����jAp��x8ː0FV������A�Î1o��.��H���$_�WD�_�;�mG�.c,E�Y҆PG�ť���` �1�P/�x��8mm����k��r�t����ٽ���RP.��0�^n�^*by3o��:�XzU˛8|N�G�ۺ��-�N/g�S2����-w< B�>�����ơ�7�j�3�~��Ue{c�5��`��o)0pbgo��<u��z��n�Zٝ֙#*cR`%`�Q5?���,G�_�z�ӿO.SQu��-�8��9u�����|K&Ԙ
EfO�f���U~_��~//;�b��S6��n֖�']�DZp�o���d��$h�ӳ=DZ.wg���ۯ��48����;ѥ2s�Vv�Х�����Oe/H}�h
�Q�{(�DU��]���(�$���F������l����,��y�a��'	Ⱦ�?SnR�ᩚ.Ύލs_�5%f�����x7C�y�x��ж0�vE���v9o�~s��]b-wUs�0WP�NN����	��9��,����8S�B�s:K���ơ��n��=jkD��G,�������h�6#֘�b;-����}�]t7�)��rݺ��9�'�#�'~�1ʮv��?A�ƴ��j�O�p���v68�_����9����rr�
%:{%�v�䢤&�]�z�>���I���:���G����t\���5����k17Y�'$��Y>��}`��qI�\����W�La��3>�)\ؑ������PϤ؍,kg��T�~T������t0�Q����!@L"��N����qq�.�v<���_x��G����V8]��N�×A���ΛoXD�RG���sNi�OG�&T��x$X�`�gHU�_ʷ���z�Z�KJz�`��f���w��+>Yb�Y{�
�-�xZ
���N������^sU{ڤ�j刊���S]R����i! �٤�JD���w���
ޜ-�d&S��p��6�T1���#|9^�X��Y8F?�-�`��j�7f=���:��)�����3dCOG��.̕2��z�a�%�G�,[^Jd����A�0�!v=���/�2ӻ54Lb�W|ss+@�}C�U��4M�.��c�4�@3��F��.�+hb���8�>����'�brc�Q$��
��a&4�Ek�^�M߄Fp)���!�D$�����ɴ=%ږ��*#��z��d�^��:�Y�8v�"���"�F eN	r��5�"%<�_d����u�� DaT����_�$�c�'q}Z��ք*/�dm��ϝ�_���
�ŉͫ9�p7�5�L#�,5(h�n�)��@[�`P�P݊��V3e�l��L�v��'�bA@8a�0f�}�>�5*���V@s�Zį'Z,B�����#�>!��}hZ��l�5���v��@�&r�A�`v�=M2�����d���D�u1��7��a�:�Ҧ����+�_Ճ�~�QI�%�4�"�Pn�pW?"8u�m�W0�jY�.�S��㨖����=�T�%0�yݾ���]6��)=	�Z�,W�>j����.�/"���bO=#�(��5 �{�[Y�����C�����~^�%��F%N@�+��E�6j
�@�@�ֲf�ht,U���z������t@��Wegh���.E��n�����{4/��J��f~G��4��GJ�|6�X�	��I�@��[�������1!��˞$U����֬s(�EJ@��=*�Ҟ>{S����~,5b����	 �ʜ�S~�z7;�������Y�@��$�MG�P<���/rhaS�G��>�W�C78�Zu4�Wڪ1qE��W�P���b��߇��/�Vphܡ೐��'Y5�-����K�x,i6�	Ҩc���/��y���:����X$�D~A�������
�--�r�ҋ�d.���SH�u�����芻En��D�vV4�Gh��3>Z��=�a��\�Ox���y*2��S* � Zo�A�|��9��X���PzH��*��<s��z&��I�����<�ݑ��Dv��g��?s�Pz�9"�"�ʬ���2-�/�<sơD<����R�EU�N�J7׺����nB��������I�ayM��UUx� ����
1m�n���  �	���bv Պ�\�fՁ[�D���r���m=UC�_�J<���XW����Z���|(S�3(�:�mܠ?��m���߆,�l��,ﹾ*q�kF�% i4� g��/ɳ��[/$g؁�}/��l@�w���s�)�o���i��fͼ�'���>�:>�g+9�w�&�8�]1w�1$�bo_�
,������D�J�:_E����u����Q� g�]����ͳs���E�#9w�5%DN��C�]�b�i(��44��x=~�N��u����+M�E��7��T.��]�x�����GQ�m��P�[�OD�p��|����t.z�t�h����n4�ȭ�7���Su}}?�"�`�$�U����3 �u5G��[zh�%C���N.�{�����E@����E�j#�Pa��{�S�1�0{��k�݌�>��<X�^)J���,d2#%�(�TȨ��(r �\��Af�BJ�޽�Z����8���|�:Y�����_,_13Z�O�+=	��HڵÏy%5�Bw�6�H��{FJ�9ZC��?��3?�0ɥs��褿VE;:ĳ�^�^J�̖tNKGc�@���^L��gCYd���(|k��u��l�������ĭ�F�?&��s[P8uxl-TS)4<�� ���� ���0���j|-w@PC�C����~V��΂##�$����Jŕ��]B�G�l��&�r(�L��N`@����v��:��TOt\��&Q��F��n�+d2c��o�G>�e2��ß<�� H�Z�v	�Cͯ���z��:��R������&=��
�>�eK����¬;�~ک�"�����4C̠d�V�z*��Э���{��S��6 ]�
^��p��]Qp�¦���e���Y'g��{�L���"p2���x����g��m��pl$����
� ����l���U�0�A��	W��";t�%G랳\}5��"k�Iu���&.���5xT��&�/��:��U���|@��'�tYj��kE�q�Zu���Mk��`C ���!�5ْe-}��b@�)��F���B�}�һ+��Q�7^�m��VA�(d7�)Kҋ��	�{B��Y���pd	�<��u��xͫץ��#߻f��O������X=��!�	���̫l��f�}��b�"�0.2kl�����Q��)�p{��-�B��ur��[���W%�7d�fl��Y�(a��G��L<�����Di
,M	��%�b����Xzfd������iT �_�>��qQs��&�"ˀ [��8,���2�@x9�?uϽ���1�+��=��}�@`�Ƥ��GfhMD�m�X��"\�r[G�2��^~P��`����������-s�{]B��� "�9���謔F������A�GK�Kq5oA�h*bJk�P#J��]as������,C��,����}��c\��=ߨ�z �'Y�}i*4E��#|`��X�K^�OHN��MFQ�z��RJn�؇)��_��۽�!�Zovn)�F|��X5Z<d����/����s 9Z�,U��jF@ڎ�gO���^A�e̠�t)7iHA	����*�l��u��p�F�QF���w�Xbԡ}���Z�,z,�{��v'�I��f�7���x���#��pZ��N�� q[S{��?���?��~�4Iݨ�X�xTM����`ӋC<�0���w?�ıE�_��ϤJgk]Y�@�\" a�R�̵3J�X��!��(�JW:���F���.�[o�j]�k1�MW���܋)j�+,�%�;�,X�_5ꃽ��p�	|��oĺ>���`�n㰞w��{x���y����Y��o|g�n;����ib`�Q���a?�-�����k�Mq�9`!� ��hr7B�9��t) cM&�S��
��f�9���(�K6�z[����z0V�.D��~��A��8w��t����"�3?y��:�
>l9$qZ4s��vK2�.�I��]I��4�k��몖���ۿ�]�,wB"i�'z��b��?�C���z����q�Պ�V�v�'VW#�T��ӢhEN���jz��_�(.##��z*ݣU��Ռ+����Z�,��#��<��o�����v� '���R�����`�8~�7�)�	���m\�h���E�.O{3} jlj@%��}lƈ�~`�e�O��bV�S�o���ru�
����\xoI�0ä��
��E���*Q>��l�	|��>����8� y1��XP,�����	�I����MƝ����_���_�Sh���1�sY����z#��G�[��6~?lt�g���k�>�g�ձ��kE�D�q�����9^f?�;����L�����lX���ͫ1�ݘ��'���o3���'B�L��#�&���ޢ�կ�Ho��,�?���� `H+��^T��Aa6�p�	w������'�O����; �)���,Wd��)��qh5*33�]!�; ��0,i�ڨ�j�zs�}����l"x\4��3�頝0:�G=��Ju�K�KC�AۿЮ�."�oj���`@��[X��E�o�/�[���^�ߵ�!E�R�:{�������=��ٰY]��M^�8���3 �_J�я.���N�*G����.�ݏ��n�����/��l�iR���{-���u�4����io������Sd�Rt?��;����[pDW�G��^FU<
I�˳�����������G���n$�j�'v��U~ϑ!s��Q���=.�J�V�J��){z�~U�����LT�	O[fs���jz��}#�mp Mo� �������7P��Q�[)��`
����?
�JĤ��>�m�j,ل�6Q�dse㚾����=�]��ZwC�0��r���m%{C�daB��-t�u���/I6�ߺ�f���Ep�W`Y�tMK�F}NC���o�$�Ŧ��ɕ����g|�E��-�,#��bݐ�����G���<?n5T��p�t˼���\E�d�Q�B�{�ф�ęb�e8���b�:]�x��U.�b\m�p����$ �0{�f��6�'�s��Ra�K�ͪ����6�f�_����c��/�Ś����.��}w!�F��j����LϞW�p�!������,(Xy0����+\��̵�-Wá@{a����V|̸�x?t��q�i��d����THB���QL�0k@tgn���'�V+�64Q�ӻ��s�b�P�v�+s��|�-Ɇ5b��Q۽�����+��1� gO<���+k�R����oJ���e�a#�A���*�S��_QG��z��4S�G��Z-���>���e#��hA��E��ޝ��G�,o��k6��<��������]��l��X����T�m�H
I��}B���SA�>�HG�p���ߝ���Q�L���ѕF�ѵA4���1/s�s�T��
�S-ffr�}iY�^�Bӂ�w=��I+D�����32�U
�W�]�������1�(�F� ��X�����^&t(QO�,� �2Q?�C����>e�Xr���x��j�s���6?R/�	}��#�X�W�x�Rif��ǝ>����ѭ'�X�� &z�������׽�"恇S�#�wcZ_������"�gHx��g]�`�}�,�!+&Qm�5:�!�����q7�&[�m�D��O���(��:<F��'Aq
���+f��3Ny�X�3��ҿ���DP�W���x�b�0�c?�U���;:q!D�-�?�ͭ���Q:`�hI)P�䴷��n�dvꆥ�KW�c��7�F�M��q�ގo]��9<��s�/���˥��n��^�=f�E�2��|�Y/8�.�B9�}��.'�03�Vf�w��(Km�	�#fx�������Z�Ë�>�=���iF�[z'��#�%9�"���BA��i��Ӯ+�CP��^����I&%Ʒ�c����s��U�D#{����Ӿ(D�+X�
'\�;�2��DinQO'��'��B���Js%_��of�e�aVT#q�"A�ϯY�8�,�`Xi�� Ʊ8�V>�$�b���>.���ͧ�'!�w�e��s�nw$�8y�f˺����N���e�����0og�c���kт�T�)�,�[��q.P�畜���i��kS��BT;q�_M~�����9�Eͤ7k�zR� �I�E@1��^����|�b���M��"����
|`��!��Y:_��h �T��G�Q�E�ѥl�Ȁ������b߭ꣃhH$I{�ٮɷߞ��h��}�����
͕?��A �&c�s
���k��~d�v����N��ۙe�3z���G+u��!;��r���m|��0c�ݾ�2#;��K��+�V7;~���?�9���9��`p�����t�8�a�xM�BN���6��igj9�
��G���{!5�q|��U���H�\�#�B�eYTz�.4�2��Qo7�V��%��ۭ^LK�t��G���ؼE?�qn�O����C���ŵ�@p�̈���S��#U�I�$�6I:܋A!>�h6�6�A�U��xaH oӦ,{.2eZ˃�Qu~k�uvj�[^K�dzܝCi,����N�%�p(�k2R�y�/��4풒k�|��� ��`��Ԡ�����%֍w�k�h���{��W)���8�hS��B�o.9%�W+�dB�zs��dxW��\��8�H߅#��3�gz���w q|��`�;�"Y�~�<�������&zΝ�����~  BN�U��6�M;a�*�@�E�K�4���fg9�7^�旴1�I�d��E�j[��l%k�$�r�e�!5`�Xo�vI��.�"��}t�э��c:�K��([o,��9U�������p�@���nF�
B��d�$܁�>;�e����j��"2�M�х�j�4-\������ehզ���n�k�[Q�:=�����F/�#��~Px�I�B�b�<����-s�ޥ�uh,qu,��E��fF;�'et|����ߧt��/5����Q� �O��˼�mXU�9/�����ޔHZcڜ�&#��\6(Nd�O�fNMQ��,�˅��1��V/r/��wx�yg�J }~��C�a!(�"Q��9���A�p�����*2��j��B�m�$v�`2�h��q�C<�9?j�k��0� ���_�'3[&�/�%�3kP�m�a�2�9��On��>*���.D��|XI�&B(��Z?�>\5��[� 7g�f�|2Ie2�X���z�K�r�&�a�j��p�T0Z���rG��|��u�5�J���nΧe�������ѝ����Q� V�~ܫ��Ϫ9_�E�0�=e]�5�H��ѷs�b���U��w?n�/��ə��R�������k�\��m	ɸ՚��⥪�E5���y��{�H+ܹw�~(�fl��̈́0�h:��ǡɐ��� *��1�����nc�ުI�0wp (��f'�� �?8���j�bZc�O�R����g� ;ؤ���?'�M������+�}n��.��t��fSJʗ���x��8�TB��Q��\�_VsE����#�ȆO(m���b{"l#o�l���k�sm�]Fd�y�K���hmJ�Z`�b�D�5v|P�l^\@�WTx��"<���(<�ׄH�`b��2�&�����8-�z-A$d/�&Պhչ#��#�y��k]FC��S~�K��k@� n�Q�7"s�yK��%P��J���V?��O�^@�Ƶ��Y��#��7�$3GKL��Jڊ���ồ�h�e�$����yǢpDxVmi�y�}���Y�0#W�@4<h_�ƹ����U�wm��F�]�P��\�h:��n��O(����v�5g@pEi�a���ѭ&hp��Y]�,�SLHXt�k+��8����I7���X�9���j��`G����+���*A��#X�Ϲ#^.Lom��f���U�hD�`��t]yw�Rb��Gʙ�,�
�\h��u��i��!~��D�G�0��q���w�܉�(��NaJ�Rnת��P ��Y_�%�/e���8u�H$�A�{ߘ`C(��`
\����5o�����̾��olx�_qDf�¿:x�.)G�AL�6�Z� ��)�����������̟8I��H� =9Z6"��_T��N����An@�.���506��j��I�����5���K��'p7������2��+z��n/.g�� .���oЫ[�I�nKI�Fp~����F��*y���e,:�����F�WkqhyS���ϖ��l6T��n������/Q���gZS�U�'��4$cb? �(Mﴐ����Yى��'����b�zB�y�װ���X�6sC[�+;��2��7�;�1W�W�Eu5���[i6�ǆ�Ip��џ@q20�xE���,��j�����gZ¤xe�2�'[@y�� �vݰͭ��E��ۤ��.d�^�\3ksUO$J� � JtL��`���;�7�Ц��)�� ��V�-|������/O��`�B�|B�.ҙAb�ۀtc��{]�UG�� �EK���o/��R[�1������d2څ_s̠k���������O���=����}�>m�	�z�e�#L���n_0t��U�hV�,�?��;o;�IK�MH(aKs�N*��<�/r��ɫwu�7@Xʙ�=�T�wظ�9��2�$��L ����nTYW�+	���A��t�:Z+��	|��w�|�\ms(X�lî_��C:�F:��������������\�ͦa�=#�lb�]��C�~�@_�
����W�H���
��CX�j�ש\���Y�����`D�{�b]i�ϖ���yp�����~�^٧f�/�=��������N����l�v��ӰL�����R�s	z��Ȓ�_�l�߬!n��Q� ��ϥs,���/��?�\�����/#�W 1�g[t%S&K0&Il�!�-�K���D�$���3���$1Ή7�O�*\-֨8d�@��v׎������i�2̜�tc�?
4��}��g�ud��ZtU1ɯ����y�q��_�%y�.9IG�2��4@��+�zm\̋�s\˖�M,��mXp��u�Ή�"�L@AԄ�����ƃ����7�*VZ�9�]��U�7%B�S��Ί�W<u�x@3�0���ռ�=P���0ci7a�L����g�c��4$��ώј����h���t�RQ�I�@߀}y�:�CT�^(S�x��^�щ#����DY��Ȭjőþ�=A3{��j�J'_̵U���%�R��i��zn"r7j��?���; s���,V��iܖ�0x�,]��-㹠�0�3�K���*_�7�G�}�8���̩��	� ��N��À^t�Q�0�#s�Ib7�G\o^㦆�k-�0}L�Vs��Z�eg�Q\A��Қ�I��^�$~�jp�T�.5�-�@��2�~�^}$�(�.�Çs}�=n(�ƽj�0�!�(r�:�E�Զ���t��As�T�ۖ�@a�K���Yb�Ma��+.�e��v�C��ѣ��S���	�%OC�]�!���]!��qQ����������5��6�����ɋ�����P���tc2|~3
�����} ڔ:"D��oJui���U�e.��M����[��V̽�)I7�<���Ϲ�̱����ك؁��HN�T� �d��穫�9��}�B:K�:����ε�ʹ��.�Z�+���x��7�פ��������Z��֣�pB:�X���d���A �_8�s� �b�2��M����v"SX<��|��sg��`�+�jC��`$x��6�s��j�~uX�_g�At1@�q��oάG4ʧ(��p�$ɪ�g4��k���J�]Ų�}���r�a�К�h5�.��	r}
m��C�������Y��s`i�ds������ۼw��ތͣ�8��zה�^2�ӣ���'U$�q��J���E��@��§!��G7���.I�2f	�z���#��g�����\�tl�θ>�$�@�OS�#�O����:n]��gԳ���2Bf,�V@vᑭTm�������-����>�q�F*�R�Z��|0g����Vl*
��U@��Yf(�N�k��J�鵧+ی|��������[�*;�~�t%�%~*HM6l)/��7ܰ$��b�������f:2)����W]�fN��W�cʤt�ůyݮ��}G���|��*��Dp�k��;Q��|��Zr�!��Ժ��kGJ�A"#M���y�����\����+�}���5( ,���2���r��c�j%�%�D�%/�ߙ���,�D�*:�� �_&���B~�$�%��xV) X&+�f$��?rk.W\�t
>�@Fn@�J�V��=�NB��w�t�5 m=�\�)��Q� u~���o��b���v�r<]K䲙o�o�x���Mb��}ԇ��*x	y��:	,�9we�Kc�J-t>�u��lՉYx*U��5��v�,�����0⑈X�m�b�M��U�׊�N3a7���9K� t�a���5�R��{N���ݚ���JC��3�.=-����j�{�����Fwzg�O͢�8���UB�q�J��t:5���*L�U�ne���X�k0�q�z�㼡&i�T^��n&�SDZ!̜�p=2_΢��U;�����b(��/�M���!ʊ��J��rZ�����p6Ҝ5�ӷ3S������5���H¨sNA���?���ìO����%(-Àڑ�O���@W�]FPKϨ�90�O�j�yv�7@aR����
��Cl�@��g�~���;:<m���5X�D���Pυ�n���vg����b����^��Gq\���H��Ƿ ]�@��0���b.N=μp�c���*���"��$Z� ��Y��8Vg��R�'R��EY0+U�o���In\�O~�) ʫ���~0��)������3��.lw��V]Z������6�#-�~̮`����u���{���,G��W��$<Q0#�{�&I�@��J�ȟ6ų�g�Aؿ�x���`Δ�|/��C���m_�->mos�����z{f�@J�S�����+���]�קqzS�aE��k��}/���?\B�_�X��Xq+Q/7��%N��{^'��ez�k��)��;%	�F�� !{KB��ҹ������f���s�[��[��Eu��m�]���'���(��]�#a��MB���O~��*z���9�U��&,��'��m�4��PH��"#�K�T	�7�v6��5JޗϏM# u-�Ā�Ee�x��7��*�38yE�2�K\?�u�z[�?)w����-.;���5�n�3Ⱦ�4����TN��|b(�g�f>�΢.�O,X��q�o)G��qE[��s+�e�`�K#���ꗚ�|8�[(�l�����^��/T(��v��H)�'�
-���f�o5�Q[i���SPp�V�c��C)]�e�)�1��� ��-�!P��g2V2ʰ��Z#U��Ё�Di�I��4|�/����`O7��а�G�ґ[qj-}ԧG���:���@��F�^w��p.`�$ 0#{�D�e���wx'������MP Ò����e_���I�bQK��C��Q�0�G�fg���=t���
�\��ަQ>��@U0��P�m�d�"�6FWlS����_��hE�6fm#�����C 3-<��8��3��N��5�igZ'4/��g[q���j���P:��݋mA�ע�_ǫ��kշkNRETv�~نJX�{1m���ܳ/����I�5�X/�	4�D?K~��g�����:����Y��ŵ�cH�")�̖3�UTy��Zx��_�Y�z���D�z���]sd�f(u��i�\M�1����!5vN��[�BBU5i�a�K�{ѐ9j��4v�3^9%�)�s�0�6��������� |#XP 7�g?4��9b����Pd��A ��W���ߧQd����M/�"gT���L[o@[����`�?p�r��bP�OZ�����)���G��Ő���3��@	�&�qFzѦ2����4����+�`���v�L��/��/C�i���{R�� _���7R�7��I^]�����;�0`���[M(9�l��^@GfA�0�WC�fhE�K; �,*��v���jV'(�CĢI?8�Z^�ڴO**��NuHܞC��o/��i����־y�UD��Ԛ�(���^C��%��0�XʰK�=<L�df1��y��9��j����=-�8uߞz��GA���^�4�%�7�_?T�^eiX0�0�Q����B����!Q�����	9s}8�� h �Ӗȵ�ph0e��AV��v��!�mWJ/,�4�][Q�n.�@&~m~���Q?����=��8@�0rw��{��K��`hubG(>�����&�@���B��)�'�u~���F�H�b؍�pl�0��[��8ބ~���{�˞���jB]��L����]kK@D�1�V�@C��̌l-����B5 ݸd�z�	:��*���_ո��C������{�o��5���5��75Yܓ�A�&'8 ܖ�VX}��&����i�@�wK�� �_�j�s�x0�K�/��m�����8ْ�l4��OM"/�ev�׌;c���<3<�0[x�ɦ����[�3j���4B���Y��/�&�l��P5y0�b��5@�>�]�=�
s۱�B���3-�|B�P��[z$2iphW�i�a���W�����4�V�p������;�b�0�]��d7�qf��Q`��c���-�D��)���t�����8�62�nD�b�3��^m�0��:8��P74&�F�$JK��g��dx`�?��c��z�'I���K�#t���6�XS���_;E!m}���M�N�>1w�lq�ɞ�|D���a�:u$A�����11"���Zx��'X'�N���ww.v�h�m�?A;�G�gq6���hD�������>Fta|�W�M�*�ɠ*�L3�-���q�[�g'��^�.���>�;��{yo-&�<
�������l��ts����1u�Q�׽5uw�3����A���Nv��f�G��(篣��::���~}!^ꇡgL�8b��;�|��񢳋�p��� ����/��Ɉ~9!g���t$��&?/�A	yR\�^,q!}\j�� �y+�d%�;,5Lf"	��6^닩�:ډ�[��nU�C|{��zuH�}�#�@?�LiE��y�L�^�O�q�s̈�ޫ(����X|%}���%񤟷��[Q�A�=�x�*yE]3�W[����pV�B�B�!�h9�T&�r�Rw[�m��r�ˊ}�̛��� ;�_�$jn���J��n�xl�6����������ϼ�$e��Fm�A�\SXݰ���*5��7(�(�q��lCy�A6��0�Uz#�!|��| `)�gD�� ��gNg�l�<`;y��խV���1�5₫!�{��D/��Cf��.�
)�]����g��}�cmkEw��� �oW��Q�|�F~�\�,�R�d�E�R^���`z���O��JpbIY�
7�d���P�#8�ܒ�T���{��c���	A�C��ڊ>y�0 Z���qr�}]�M7t����C��H��u��t{`R�F���˭uFD�^�vb,�[ ��M�l3["�e�ZֹLhkM��'��Mz��; ����dJX�|衑A{y�S,6ŵko�ż_[� ��`ү��.�(L91��)<:�If�9�V���%a+<�٦�8�amה�X�Sw����w�D7�G�6&��˰�p��[Zl� ���A�Gc)�@o�0�⪼xt%����0��F���ȯ
p�V���u�ܨ��{v	-6����xj6����a��٭�o�d����Ґ��r�!��(P;F i~%ֱ��k�w��$x%�}y��~�h�&��R˸.?�=Δ9��Z���X�Ĺa(%.G�0Ɇ���.`dSR`�r�QfX��6mMW�qVeJ!�w��x�)�yBgػ�M��E���kD�;$6��XS���mC��U����-�0�%�6֝G�j�����O�\Y���^F�y⤤&�0K��T׫_�[yJ�*Ǿ@�5[T�B���$�$4�k�@έ�����WuC1Δp�@��lE@>i���>&�=Z_�.-�&�P���q?�;��pM���3V/���ktq��Vצ8�"C���8��n���D���:�l�nL��e�j(����v��t��2�F��i:8��[:3< ���m6��:�~6Ve�ƿ�r�����xf��h�˗]~�m�<3:w܅�d��gr���p\pM��
mG�-3|��P�ē=_�AK@S�n��.X:\��\q�#���mo��w`]@�M#V�v`@�&_O�H$܂�T"�����S-�{_���H˒�CT�ch��Ľ�?�3�4A���K�cE�*N���%B�f�I���<EۣJ2	)�U��Y�.A5O{\B-ml��P|Q�v�B9���Jln&��&ܵ��&�2�
,��pi<QH6��4�H�N�<��A�"彁���3�$� ��X\�
� �҄Rh��;b�.\�k<uM��x���,w�D�\��N�MD�r�������q,�Z�*����2������������n��.�Z��Maչ�]q��}xMZ�-��2	'��+3���ʎ:ܜ	��[Rux����k�Lk�`��&���h��̆s��H�DN�Nb�Z�ʘ��iʧ'�+��̸�j[���S`R����Ff�f�	bxb'Ot'�P;�;�z �J�m����!!��66�����U`��dL�d���=Y�ӅW3Y��q�ӟ�\�3�Lv�}�$�
���}˽��!q��wIΕ�N�}�|%�鮒��u��꣣�oA�q��$e�y�7�!-p�VeUK��;c�ei4�E�9c[����R�s��]�����`�����A�0�#V�`� 󑕗�z�6@�J�����N�ЭV6*�d�|3�_��Ǩi]�C�o���֟�rҎM������\��B���h'U���Ysm���)=���r;���:�Y?�̊�S�ͤOs���m��v/<�)0�w�J�T�Ӳ��_����q��y�tq�J��d%�~/{��<8���fD�^�=!�I߸����%�M��,qtW�V=��W�%�7��_(�z��s@�33CnQZ�n��l�m/�������̼��t1�I`9�-����fK�٠C�N/_'�@� ��g�@�=���v�a��2�D�@)�w��I��%�mEȩ}�t�H�M?�	������9�� q�g�6%���1%��X�3�s�YD���Ѣ{�ʾ���}�&��?3�jh6��F�Bm�<�r��I]�Y�>���^����pNZ	Tj�DƷe��}�o9 �s���dWc3�rrp[��Z*��]��>;�,E	���\<9 ���6] Z]�A1n�#d�jN{[3#�V�!U�$2q5�G{��?G���k�v��Y�ݬHd����洢��롊9x��_���t�+g~�6p�		%��济K��%kP0b��"��c�����Q��e�L��5�hp���,� �gX�+�npP4 Qp�>N5��Kf>JX/�(18��TB�fi#n3T����![�'�T��J�s��p��Ì����tf�D�V�R��9����p:&�Q�7�MS�B�c���\�^�F$���~i�i�ϵF�?b7.a���	�Õ���)���/��:x�OzE��b��Ga"ip��\֕�\pӦK��Xo+��]���o��s�r�X��0���ǲ��;*��P~�\
4Rw�Hj�K3��m�A�kl%v�c�� O[Қ
�� ��>�Yd��Е$1G
A�q7Kn�G���a� ������h����;�ͨ	f)J/�I��Y�Pw��尙 �6�AE�;�T�-4j����Bu���F?�[� Ga�*̹Ĺl�Wizۑ��XS�l]��G����-�u6�9O7'O���[ױ��3j0����)f�j��(�!�٭���4�[����>}f�$
�)%K2m:����[3��ʈ�@�~$HV|�E��� �#�^X7
��]- �ĚI91�Ϳ\Sq�mi�NP��1�7:)S׵��j/��K���f EF5.�d�RL��].�DI8q�>�hB�0�KK���}� �a�o܀$�o�|3�cˤJ���'V=[��Hv����Γ�"�j)I�H�sE���,�z_=y2�0"2���%�aC��C���hu��ȕ�A��'8�ܴ6l�k���g�I��� �)�%�]��T ���oѭ%K�����\��H!�/o�1��W�h���.��l�1U<
��[��������.nXx)s�k���׬�iW���P^Yљ/+�OC�<UC{aGb5�H�(��aE-c*�gaf(��vK�G�T�Ք�v����M-�#�U���$��-�E,�Fwl��"����t����S���I��¬��c��k��ɲ�� ��N}�sp޻�2<����=T�$�w��>k$c�ꌈ.�,ڟ��<t~�X�s:�B�:�kp�?m�����n���阆e� N
(�#o"�T�x���1���|���І*O���Y.��>���}e�x���3�!t-��+�_��6{Z9� ~Qبײ�6�!������%�}=}+�e��4W�H5V��Pb�H��a����GX�}�m���֢�j{&C���zW�"�j�R�ޖ�P :-���o�M�gf�w�*IC����^�UN[7�����7]�V��gD�a���;�	jF�b�q�i-���)!�S�a��j�}�v
**]�<�րk�=��#�8Fm���kX@�����ꘛme�?_��h�1�O�X�a-��'*;KI'*D��Za��}�u�.��p�3�Z�<_=DVg�;�_����Z]����x����)Mӆ��]�C�^�N����Wl�#[���v�U082 ɳ�q��DǙD>�}���[&�|�{랚�0��R �����۩2���s�ɍ��4�נW�آ,Y����p������2�R�Q&��_5?��W�j�,�p�����빿De�W��R��ihG��A�ނ�p��KX���gn���C���l�!^�����ZjL]ؙ������Q/릹���V��^B=�&��3��F��(�+�����	哵���2�{��҂j'LAGa�w!����v|�=�|'�� ���:7��+_��ճB޻�E0�x�0i<���;���d���8X'TÓ�\�G��L
�|ݽK7��(�S�Mx;�e�ˎ2A�rQ�� �ՇTOM��E�hk΄��)|�#`az��s^$�^���m�R�	�+����NlOk���ճ����ڒu$���̰�#,U�Z�N迧'�{iY�E<I�lP��=糍��[Ts��=�ނP_S�k�Ɲ���eh�p��6ᙎKUG��>�,�����n�A�C�������EmR�hC�%�U�d��n��*m��4������K�x�O�%��:����c[�"Y���m���N쥭��n��y�}QO�o�m��K_�j��|�M#<�A�k(�*Ǆ��b��_��J��ř<�'V4$l�ݣ�4M���Wq'q�C�-��k�@����c��2xo�\-=�����`%��]��yG2�5Ե 5�����ǻ(� ��ȱ�+B��qO ͬ
�'Y�-"x�W4�Y�����CR��'�C�̅�d�K�a�8����ha�<�n3bd ��S�:���O2��ٞ��U؜�����n}�1��[�Rc:	�4�)uvɔ�1 �_��I)B���B��&u�S�b6�f����(y�����vl|��1õ圩Z��K�+�1ͭ%3' �~���=����f��MM�f���(�$�YI��&�-�8L�Z� ë� �x�<������h<V���i���&��4�F��ɪ�@a(���f�ښl�b�d8�!r���]:�Hp�q6C	������Z���P�XݑdJ�C�ȥo�2~�9��%:~�[�Ej�cX���̳F;�|��k.���+��/,�z��-�{>����M�CW��K�|�5���2km�ߕ`9@� ����g͋W�v�\~r���f�m����H�!�z	xp�TC���Ԅ�弇cH{l��G��_'�n�2�+<��P%rpSU�MA\�/*����2���}���Y�r��ِ�Ⱥh�k���~� h/�?o@MU�d��'������锘_ޮ턧���dyNW���g}�F����Q"��;�01՗\I��@	�ӵ�z
;h1��6u�m����L�Z}g!V�OF������º9��z�6Y;�dԒ�k]��ف�i�^���W�����f��<�����Q[�#��7�r��|���1���*�tm_v�f�e��ʵ`|����*���:r�!\ހV�t�q�m�e͠�m��8��<"L���8��u�qnF��_��X<�J�	%��Yv�'m�# I}���tz�=�V"�����I�a�뉾��V�x`�V�`���O�x�驄��$1�]}X1e�VD^+)�rr!��y�mݾܞ]��5������$@�E�j�ͷ�@:15ڏB�L��R�y�O�����<O���ǟQ`�Vi�Ec�ԫ�ܧGD�ۚ�*�d����U
Q����B)^�7�H���==�����RM|�C�
]%,l��i�<P��g8E�Һ�mLc��N]L,��cd�5�>P"�ܩ �!L ���.�@ ���-ї�k�M�/h8��}4�οj`�&��J˗0�I�V�I�l�k���MV�4�v��ǳ��V�R�&�T=r) e.0ȅժ�R��X��Z$TRQv��`�}AXa[�SQ6�C}y.���t����͵��=�8�I����}[�.9�3 R+?�Xu�|&���Rø�J8B��lB=�1��I��cIH?�5۽��f��'��,[f#��?F盩>)rM�5�qي�U hbs7%Ѷ���E��N���m�ŕ
�u�q~8$�=�Uj�fF��t&�ޜ�*���l�_~+p��3#���FѺ�ܻ;�?�4��P�;
�ס�(��1 >��qQ��\{�GX���+}}�S�:I�/Op�BLJ:��V��j�U6uf
-)�I5�6ӟ\;��=��b��L��j ������w�hN�o��C"Wq|��B���!���AC�Y�y�{��	˗V=�K_������K-K�����qS��ԅ�����[g�hV�@%�"�q@b��$­3Bd�{�� Pl͐w�/;�:26�t�x����/.�uC���Lw�R�D��	e�L��F��PVd_5 cd�a�L�;b	'����7;Y�!u)_m����	ԵO��P���|�N:S@��G���4�P����("������a��5&��_Y
4"�ڽĻ�]�W]�;�$�2����F�Q��23＾�5����&M�^Y�<�(��u�N9˼���_O-FGO=�r�W�)R� ��}� B�?�V.t���4<'Iw~��J�
�Ǜ��8�52���f�~���
0�N������2k�-�`��./r �w���0Ș�m+����Q���g�j����˳�:�:rʴ�d������Q�=bii�$���LN�CzW�r8G5�ِp�̃=��C��0��u2�LJ��/܌����{%��U���=�
����*,Y��[o��v�T�Qo ������,@j�:���#�:<��T�6�x��	�ߊm��V#�l!�5�J�̿5���F���'���@T��U�	V�0	��N���u yW@]�X�ܔ���C�z.�ɯ�gJ��w/�>�Y�w�ª���C�҉�գt�H��eޚ�ݍ�ҁ�Iˁ�B�Ž�Ԣ��*tՇ�����/�aj&�W�\�r�A��+�Ӥ�$#�KQ�E�����7Y70Ŧ��Z�j��z:���T�F�� �l{�����m�>5��,[�;�e|�A�	�M
��]�"���1�H�2+cKRm�T2����J�ț(�$(����!������!�Z^ �:I�|�9�(A[.J�
�jqdc��򡟉DΞ�>,�mL�[O�ɂ��@�j*-Y�&$�Fǫ����N�s�2��C���h(��3�64Mf��-��s�Qj��o��է��ժS�Q�N;��Û����<���6�h�ᡦ���9۴_�'
'�^�g�;�x�,��������+h�fJ��H�W H�_D�a�l��@��X�V��E�V�.~�����q�?�c�K��)R"�Ǆ����1&��L(��w��T��{�H���]�2]��V6��ڼ�^D���+w!/͞8�����0��f��h8O(�^;����Ì�����Q�m���K�H�Ά���X�4|��S����Tv&YU�'T!*�@o�B�ȹ���=������p�RQ#�=��W����w��>-��ϖ�W<�fV����H�e��`�+���#`� 'q���_�\�W���c$�Fe�h�*�(i����M��t#���iO�j�b�\��i�%��+x�J��P��I�����ך ���0�!�s�H:b�$s��c����;����z�.;����!}�\t�_f�<=�4힤�d�<�� �]�1�z� �٨e:�hL�fV�I�	kQD�Kp���6���:�:�InM24ަ�&%X����,�$Nt�B��׬��Ԡ����h���L�W�>����'lz�u�1,O�;]���_R,i:&��Ͳv$;���*D���i��H�S�Q)���P�w�*7��t3�����$�V.p��Ƴz�G�శ�����w��yB��(a;q�G����<[�����}��⸒>�_�_tZ�� yD�5���-����T��a�m��shF��מ��?�A�4X�'zx�t���¯/��y	8A�S�Y��%����U4��z�R����i^�,R���� ���w�#ϵ�3=j�7�T �{����-t(��p����~􅃏��'k��!m��4�P��1�g���N\a'�e5�u�t��x��%)�Mx�ִcE���T�ku�����NdHz�۰*|s�3��<?�i'��4{4�.�a��SZ�1qax�,\Oa!	(����O�F��n(0�x|'�[$q8��i�XChp؂�3ѠUpB4��V.�C�h��F�0��E�;+C���&�Q7�'�W�U���e�]U	�!�0�/��#��l�b�� �{�1��w%	����̗Տ�fڽ��(n��,�Xq��t��8jS�\�xЁN��?�HM�Q��Dd�����٥�u.��ɠRr�_qFѷ��D m��x��	�:�ׄ��&�g�!57_��.O�e���M)K�@J�Y1��9X5u�O�3u�9ي�q��[�RR+N�t�H{�8b��I�k���:BE?g�F"��$o�
�y����!�H��cR�Mu�2'��#�ɣ8�s=}����2�@Д
:2 �W�r�;_qa���R����/�s�2IE'��Tb#��K���Y���o��JAXͨAp�`̭UM�T�#K�"3v5\Z1Z��ɑ��@Һ"���t_��1���}�3E:���V��A��Y������y�T��:P�P�ޣ�捉��m�|fd��)Ť���J��5�Z�<s���tb>�9z�$l��ɄX,���	/�(�:m������ii���x������6�@M���mm�]kw�^���F��bҕ��ҟ��� _����9����
�9�y�H|9F���#�"ٽY0;�v�)5N�����&S7=R�z�YҜ*������w����W���t�i�4��^�AG*a�6@!a�`4��F�+�0��r�/S%y�������U=�D�A;zr,
����fŎ���s�����Y�y&��X�+\9���c��6q�p�8P��?�]a�<o�*vU!��W$}�ls�����{nW/ڒ�~A'/VZG�רB���Esy.�Zv)��dw��TB;�v|��]E�5���jCծ�����ПV�o��qcE��.�X(�,�1������|gH���ʾ�S�[X��V){�ˉr�E��F��s����y��?��X�牍��AX��h�
�y>R�d"sݪ]���W�]ś����{�b}��
��資Sb��Z|�k�Z
���X\�����_qj^Rf��8ٰ���#��rf���x��G������:c�EBG�P�����VDW��������w�9��{0ײ+������&$G
�kZtS]� .:���dh��Pk��P����x�k��U���E���b4�9�jO� M��+O��R>�{h��WOm7��U�`蒭� �o����Rob�(���Q�`�������qc�/H�md*�w<#Q�Ϫ��W�V�Ђ�a7:���5��!��T�L�ԭw���|f��3�����O�¾r�@ظ
��u�T�k��"l�`JL|0@�Y1*F.0>S���
�Y��Ӈd��0�QG�H\���H�΂evh.�+3��J8r낃Ta�K�6~�������s�5+]����A^�?!~���x�Ix��qe+c�h�� �!&t��*!w��WК�Vn��ڃ�s5��­��ַ��uXr�	�x`&�k0ʏ���[(&�F�O�>*!$�w����|��c���PV����:xW�ϲj�^C�ǦFFx$"����r0B6�q�{���*�F�r{@�&I �|+�`� ���y�7��S9�KK�8����[/� ��U�c��QA�˷���e2�O�ԙF��Y;j+������# �-��&��G���ͰA;!C"$9'��0�sC�����,+���$1�����dm��;<['EE��]e��W=t*�9d��f�
��ic��JS=h�Sw�|iR!���찭
-_������U�9:��]ۋ]ڒA�Mw��B�~q�$�#6 ݻ8���h���v�:��V��;/�S�����=�ѱ���EV�溵k-J ��t��x��M��%J*��*����:������ΟгQ�?�}�~�^A�N!�/OI��8q���\�V���Ȕ5�mY�'��7iﵱq�>od�,����n�8ˊ������ր��Vt ,�2�<���״�V��׵~z�69:H���Hn����?�Cq^�g�� �_@�҃�6�m~X��.*"W��3ΐ����k�,�k��l�T�8t�K ����!�����(���\��Xá�=Y��"��F��J=�2UiL�]�jP{�Xr߻��,j-)�b�Q�$�S�b �'�\�+�ԡ�*�[k�vE��
 ��DE�}�����,˼�+?~��*�	U-S��jl�%�pa;3;W�	x��d��`dz��D,�
����D�����f��ŘS��V�u�;�����������4Q8����[�8��M}���U���з��R�[�޷��W*%>��,�)��kt�H�<օT�d��uť�����K*R�?��?|�2nh̿�z)w�gi�,��2\�,t�Uo/Tѿgvde(H�	���B��åV���#kͥ�LJ.^�}��ksˈ�R�*�i���}� ]���ӹz����맘< �H�����;�A��i�gC�wݢF�M����ي�a�4c�KNߩ�ǆ�8!Q�(�L�{�`���U_�"�$A�b��D\N� ��^��̌*/����s���R<Jחp��B��2�����f )�|��9�H��U��e���[�TA���Q_�s�����[�2N{j�����{�HdtC�9L�u�H�������g��z��I�n�oH	���������C����"�R*�h���غ1>NQ�%7\�(�J������(8d2�7���G7([������>j_�~�A��%k���p�LN���n��;}^�`��O�I��WyH���g��&}[��"���U9A�`sCg�n�1br���>i(��f�R���W�H��l�Z'䈃�������c���D��H.U���/�1�ލҕcg� ٲ𕌿�2.8ъDp��#������N�D�|�_i�dܦ2� =#LE��AԖ�!���Iթ�?'X ��oDT6�����XRI�_�o������h;��o�:�ƿs��c�,�r��}	�q����1������;������[� i}�P{�X�=�=��^WXωl�n�6�{&�l��M2���%W`ߩǱT�����;���%�Ǵ��bp���� ������s�Q�t�v��5QZ�Uv]i�M	g�ILK����y#�)���t��ft�3]tj�ez)�T��!�M`c�K��/C?tW����$�}�~Z:c�!"�r�M�j��wP��?�Bp��:h�Hm�</��1�;��k�'7ܑX�f��ȡ��<�S����\7m#���Qܫ���/�����`x�;6b�ç�u$u���o ��g�Iw�L^�F>�yܢ7BS�Y�&;�ރ��I(�����h�x�i�)��ѭ�YCR�Pzw�c���x�d��?��e��q�+9��3\��`Ұ�yz��&a�M�5�&yQ�Ն��Z�6���36���0��_��oh5	pƸ�I��m�[�E3tp�M{N��b,������_Um�B�$-��iD/P|���%�;�!p,_%�!:	�g}���u�q�T�|��،�]lf# �4#�ȕ��Tl�Ϋ��~��!2�y���qb�6؊��c?�3W-I�C3�"��h��={4T�˧	gHur����0��9~����6@K:�հ�孒R��G�H[���)�"K��T����H�Vo.�X�\+@'Q���,m���K�QN��] /0zw�Wb&n�=/J@�O��K�����Φ5��JS��l�m$۝$��$	��d���-�Z�΍�B�_,WݣÎ��V����C��]��N}%��R�u�b��!cT�;b"��^�"+]��*[(��-8T*�]
<;��kX'r9���L��^�M�?�+$ �\�Vl	?t/%������e�+z�?��zmd%j�n��̰�� ��N`�Q\j�V��""��K^��{�ם�S�;{.�ǭ�u)b��K��Ujw鹎]�ӷ
Lva�R��B�Roo%W?i�pա]�#X������Y�uq�5v�%���9~�V�K�K#.{�rjK�]G0�s��R�:�I�؆�=7�g�2�7³2,��6�r��H�xVbڍ}�;Yu�>d^J�!4�k)��!�b���DM�={I�� �P�qR=�7���XC�܄���_���.���
�/)YI��� 
�)��������K������v�ش�^%����+�&���f���mrg�WA*����ϠOA/��噣}�qC(�� �8n�������vm�0?Vԫ��=�ut���*X]2�8jѶ^8A��8`�E�D�b�/F��tO���;/z�#��Di�YJ�a�<֠���Q�M��FQK�>�fԐL��`�� S��`�� },�o?[-�F��XM��*Gʇ��w�N��S�	�ZY��'���Ks���^c�O�Hܰ�c�ޒȮ����G����q�T�W� �_c���z�2�ƹHNx��dW)Sr�LO��jL�9wg��1�{GQYUy�P�)W�[�����gŋ�Tz�*�Q�_�z�϶�9zhNN�o���ʷ��\�m#g�) t/�Ì�Û6�O����J͉$�B�V�"aД�� �G�=��dI*c+�Kg�������~��Gn��G�<�2�l�$[uܼ���W> P�YWL�ߦ����I�[�M���.q���$-ng�N�ά�1�@�P:U�~l�(��4��t3۲&ȏ��QI5���	����.mz�Y���7F{R�,��a��|�Ek9�`J�Wb���f�#�ieE�����E�-<E�l�G�@c��P��ͨ3��<�B��s��p��Wu��͐N��v@1��H�sj����q"�󠂏��BO}Q������1Gă��nk����\g�a�[\��kB$�ܦV���K��@Av��\�mη�+v+�-*��4��@�4$�3q`DJ�S�PN�5�m! �r��?��k�LB��9@�sTӈI/�Z�n�_�O�	�]5@�Y�.xle��|��P�:KF�{�S��ѷ��q�*���,���Tk�:��X�
�X��������k�3"<���/��{cYBO�6��~L���)����{v�n���SCU\u7���Vb@c��lVQ��agb��m�J��NĤ���V_�m�"��ȯ砉b�a�&��Al� ����L �+ze/�n��YS���h9fE�Ùhv���e�Dm?��]^���!m�'��X�U�/�ytt�>�=�����.1�=Ԍ����#�D�fd�� /�~ ��}����m�x$�o�/��\+$b��	=cb"�����BL�=���q8S�1��'��V��F�{
��6�핷X%Y��cWQ>_�A����b���m��&bZ�T���v�Bt�ւ��TDfD��N���v��^��`VOH�x�������ӢQ�輯˶�8k�f�Rǚ��]9�>�|�P�פ��ٯ��7���sG;Y�,* �]�\���F�)��݃T-��~����"�]��b���څoХ��(P��D=�*�&�y�ိ�T�	m��%�!,\�����F��<��K�(�}��}�[L�]F� C��s�q����l:��E�5�έ�P�Z!��^9tXU2��.��kx��p�3�hv�J��K�Q�����7O�\0�4fmC>k�G�N8�Ly2�	�wA��L9��8�#'њ?l�I���Y�l�������h���TW���������Δ?��b(�ޛM�Ǥ���u��hG�������o/e)��Uc�>L5Bs��Ps��BcG�v3��?d�%n�"�fn=�~�k�:M��}u6Տu�̈�X�w�	hH嬧�Q��:�0���*�����6���D۱H-�hOF��t2-�P0�Kӏ�`?U��`�v��2h�6�d��J�>f2�4D��`,��q��r!'�A�#Ms޹]�:���)�Էg����4}p�J�m+��8������r�纟�.Vu��������<9gO̎�o���P($�߲@0�����}�:��J��U
�A�A�$��>�i�F�<|F�u[�#�I���1�W��'��tLLDt`u�̱�[����x�|T��ϼb���V�hr`q,R�:�����ͻ��w����w[�8��Ys3�E��/k0 ���H��`Kbv>x�*:�ԷL�ـm���ڈ _������Lq��(��9��������%�Rק>����g��$a�m��p���r3wD�M����؊���aRy� �F���v�Ȑ�8;B����9�4.]+�e̹R1lV��լl0���Ч�����d��Zp����f��� ��s�i�/�6@)!���խ��5�5b��ٶ?E��M�ǌ��±��;��:����s(�N�p�n��C`Q4N�>߯{V�g�B���`P4]��"(
څѓY �nEq��(�.�R�=�m���9����\�ɫH�jH=�ˎ�!kW˄��%:��ȭA�\�5L���z',�j�.%�Q ����`9VV�/)�������h�&D-G� *w*��be1IL�����*�����]�C��Nk"�y�PF[�d�Ii�Ys�6�l�C�, �s7�j���o���m��;���dJn������0������4r���⸋1�s&u��C��_֕���6�΅�F�#������E�R�A��2�~N��wN��T�;���f�L��B�t�'��&G#�è!�,&FҦ�8�#����3�.:�D�h��sV��xA�TI�d@���%	��uۢ㉓��(��ԑA���%[�e�n���:�crTA�0�hr0$�ә�'��_�!��w��j��\1ڑ-,�|~�&�EK��b
s"��%x)aR7݁Z���/&{+Q� �	�u�P��9�i/`%��V����?+Y�[����]��` �3�5����+{�m�I~��%s�Z�`�e��܁��˱�Z��)NCy�Ⲡp{�J���q���Იq�l�(��Έ/�7t� >���#��x�_�lXSH�f���Nm�ȺVj��P^P$�q�U���w� onǐ��N�f�lݧ��Ͳe%��7��V"�J|�~%�a��{�?aL`Hj-e�>�L���������v���c�NE�=���<E�f�Kvn5 +�ò�5�.�y��{S���릒:X��.F߯oB�I{O�>�ԡ�^i��� ��dX���t�N����*�5 �h��mL�����Q�LL�講�a(�Ȕ�#s׮�(����@�ʻ1��`�ݦ��B��L�n���'�D�JK���.;
?��9�F��[E����vNfR�5��`�Ah.�M��9��$�#��L|�M-McLq������V�m�;4�)<J��g�et��$��|�"�	�:�&_��;�%�(���M�kN�m�+[���G��9�	xD'BV� �۱�XJA�L�Ӻ�x����6���E����=��z�ֹ)���{QU�a},bnӉ�J_�*���< z�X�_P�>���s}[1�K�r�黨Q��8�5��JCx}K3}�ɕ�jAC���{��]����c�&��n��]��Q$��]�Ѡ"9����D�/�� RIpn|��)P��y�o�d(���߈�m�@�̑L�w� o�s,=[o����YjT�ME�:LѮ������t��!dZ����B =�e���1��H.Ґ���I��n��]v�.���Qw��(���ȦRL���]pۤX�k�E�A�9f�D�[m!�' x�Afg
q�;�� �W�mظRa���	����yU,tgb
P����fϲ�������ɸ���F��zl��}�풔�Z�?�	���B|׀�@������_q�]ki��&�:�4�-�rD���L�})'�U
贸aV7x�mCF���L��d�9�B�FH�8�]�K�^@�N�1G�7	 ���Q��Ter�H�mSk>�eM�7 r�P�O�� 8�+m����U�Y��B��1�j��:��?�Z�YZ�,X�6_�ԍ)=����j�ٍL�8�j�2X�EV�p�=�L4\�;�J��pFϿ��\��n��i8�6Äx��>�x2��T]"Ҍ������:�x'vV����n�x$�և�:��WQ#���ʌӄ#�<�"�&>�G�G�^E=m�i��㵴�>C ]Ĥ5=?#z�]c~z��ĩ4�����]/�ڟJ�Y�,	u�/�b���^���p=&ܶP��ύ���:�5���8&\*�@�mz�Z���D��Ye�:�?1�&X��⩚W\���ɒP��6��63����`�]�3}��g�N"���(4)� ��r+�9֛��2܃蕝Y§epd�2�hN��T�r���fx���"x�Ju�[;O�[;H;�d��3�H����)Y5���E�����o)�����n��6�~_��j�	x���-���D�b��[��Cl�����H��g�a�qM�Ry�z0�ǵFm4��/�cDa�g>���M���u� ���f|�WS�i�~6 ?+�]��Og�K���z�Htk^�^�PjPxc���/Sdz�P�N���B�9L���Y�04�yJ�μeC"���q����py�Vz8v���CD��>?���W���t9��L�����_{/���ġu�F� J��ɇ��t�}���E�۞�*W�dhQ$}�k�bu�׶k�UT�ʞ�$3<4�F���AX����J����r&���҉���gx��ro&R�&��>���g�V�*���Md�{�7;�Чu&1�6*��O�
�cm`�v5�6Mu��c�B�aA���j�.�%����� ���x|�hՈK! y�3a�2F��ȌS��r��6����}+a�e�A�pڑ#��n�"��9P��Sv��.T<<s��l��r�1��5��ƨ�Sܘ$�ķ���(2������7	XK�*�t� �j�O8�i�+�7�YYP���IC>[Q�dq��.zK��jHJԭ�O�#r��4P�K������-�p�+_F�6g��o�'u����$N�~�Vab�Tvn͖�11��4O"�7׎�I�6��BS��y�(<�%פӼyCd(,�m���Y���"���T]�fM&�x
�q��i*�.��c��;N:�;z�sV'�ȭP4F�S��f<\��}-�0I�{��EI���F�<0�E_�s�:lW׺8fH����h>��hO���8Lɰ�F��˅^��snx!6��� DB�9�<�8�k�EQQ-b�?8��T��w|_ת؍$n�=ŀ��03W=ʺO���y�հ���ʭ�<��t
dl�J����E�7��pz�L�"{��#~�ӌp������f��?���x���{���߫��˸`"�F��;b��0	s����Y�^2��(�u������"$��YmV��E��hO?�L[g�Q�F���O|
�!��j����^�>�'�n-��Ŗ�غ�ǜu�m[K%�g@�$bT��O�nV0vT=�R�腋��.V�e�&��Z �G���"�6�3��چ�P~��,�I��,U����S� wq蓵֡tu��V��ײ
��< 0j�*a����e��d��b�Q	�L;"��0��C��j?`���3�G�#��+7�`A���˔���,k��PC6�����0�>��b��RY?��W�ܲ�Y�x�*�(����MvL�">��sOf���`{q�n�B(!�Jj�wH���g%I,y�v�~��j���d·����?F)���uA�;[̜|���A��֐�%�t�h�*�dV��Z����U�vbO��E��ʏ��7�\�ueQL2�Q���h�5h����&�@ ���8^���p�qT�ݫ�V9� ���D�V�@F�%T35��k\_��Z�s�s��dц�l�S�|�8��ި��1�c 6�"T��Tg��7��� ��3 	�^Z��Po셚)Vʩ��5���j9�e��`A���o:�u:��lX+<�&��e��'� o�"�|��,/�ށѾ �J{~�r�E�9A䀕���\��Iݰ�*w䁬ʫ[�ǿֆ �)��"�6���hۓd��:z�C}�
H���0�������uo��� ���4��!%_޵^����my�N�
Gy��e�0
��u^��r�"��䠂�=�uI����<!
���Hn4�����q�ƊM<Q��[>~2iK�RF�+�"�M�Yp�`ϒ����BF�]1(@)�X��
���{�߳��&A�����(M{cybS���������>ڠz;�(���p��Gq}~/�M��=�0۶�g*�m｣�_/����.�r��pF�+F�fS\�3A�~�h��}��a��y����ß��귊���_" �vhb��W�iױ	 �o踉�a��W�!�Q8�m�d�c�BP~�n�ޙ��ʭp�+��W�y��mj�<5:�k���x���u��0�X�.�ǝ8��bVas��q<iD�,p����pgJ~�la1h��(���w�-�<f#E�������HЀ{4,��J7mOd�_-���	o�����M��V�	��+�-½�Y�{��|;�v�O�$���e�p�r-DAr�" �\�<W�Ǔhn>��h���,��?����`C~2����b� Q�$t6r �4�ٮ�D;�AU��r���5/�њ�]�b\��&�l��Ɖ���nߍ�k��3W��/L�H:^�?���{�$�>���-åd �"�Џ�����K�l�u[���p��_@��t�fJG�ͼ�1����F|���'	���ؿ��A7F_�D�Ġ���E~ �^ 4��oE��[�� �p
�IOT�,[�-(F����C�w����}��`4-0�@�Y]j�U�Vi�t⥶���g\�[J(gI�ĽЃE_Sqo4I�qf�2��{n�(���/ܬÈ�ӏ[���ē���jK�CVfF��[#A��p���E�+�F�J�^���C�j�p�o�����4� �|t��N9`��֍�\��u��9�j�m���lp�[|e���p��`4���_����IwLi6�O삣���mFUQ^>�������5л��MKH���9��m�F��瑗����Og��ɲ�}��h�5c�*Ț+�}{]�>��챮���\Fb�d�,MV���Q5�D=�"�R�f�V��ȗ�i��%�oථ���0l�W@-�+'v��n.FLb�kL��	�c	�%#�p��62NU�c�]7���\˕9�]@���o��C�d�]��e�����zJO6[��TOh�9��,"���3��N�+ᤅ���`�yߌ���S���K&FŖ+P�V��?+�U�~���I���$���q��ewD\�ޮ������'������\���W��ͧA�S�3Y����FhZg��t6Jw��z��D�;)*�|�~Z$o���˪D �=�S�3t��Q��Q���fp���p�mG�w���#�Үh~]j�������G�� ���Z5�7֜e�]^lh֕"O�g�&˿D|*��7��ղ�鹌�0t�0l:ʎ3�h��6JQxl�T rdō�L*]K\����S��)���@�z���k1J�w��1�p�ɠ%�����A|���m��2D�����y����}�������R,�����<�1~��{���G14��x��V�:04g�b�gQ�&��)�.�2{E�|)g�G�(�R]�MO��������[�E;|�l����lK>��w0\l�P����l�4���92�c~��S�� ��ig�~ա�Aqiu�IF$����!�QW�N�閐K#5MڪC
AT~�O�ȩ���̓P��miN<���p�����f�|�ڑ�1��.>@tz�� sj8G�p~�;��;j���F�tT�>�-�EQ-���ڠ����"PBD�r�4�6y��ZE�cN*���uj�,���釽<b?:tļ_�A����Hp[�aP�-;Z�����a
�yH�2�t�&������W������w�.֣���ܨ���v[����Iy���`�̐X��������g5�*�t�kI%��A��cH�����߬�(fM���`[}/�Ml�����2J{MK�L=	%��r�0��ݐG0��覩�!EH�s�ٓ��UZ\	E�V��|ayU��k>bPs\	9�
3J��ELM�2G���}Ou��fCEr�4]���ʨ�<�x�"���=��� �d
8������v��\�c�Kӽ�v�dN�Ex'��wZ�u]�LA�������}�g�.w*�2����� ���c��|��eKUЗ@��y�f�LV\'��>�����hK�>��p\Y���c	�2����۞�ւ~2]˻����Ҍ���f�f^�Ѹs�	�
.*%�+�~pSF�B�L}eKN�{��;�<��%��y1tW����d�#�u=��	E$_G��3�,r$�x�r�Y	��z1lR��sìsM(g8�2~�GP!	�;f[��gA$�����4P9���ċ�U���mZ(�0�O�=
Z"�����9ݵf�Y��W@�yf|y�pN�1��>Ϡ#!O���k��ݽ��O\�1L#�,�K������zx�����#�6v�6�>cF���������
���9��`�ܸ{���W�g�]I�A*
��V����?���Ԉ�%ݶ_�x��o:Y��oV9�$Őu����,��ƿ�F-�o�ڰ��>sV�y�C�Z|����/[�mV���e�GN
��"�pPlVc$C�����-#�0���s`@���A��o�ظH�@1Z2"�ve���tp�a+/z��n���Kv~b*�$|#�]n���y;4�s��v�}D`������RD�\>,���"���������>�b�⇟N�%� ����{��qw����<��;��)���+�,D�EG���(�oɨ�T��{䷁�� �s��$�&H%�q��Jf���v5�_�˭q^� Y�ӆ��#<Y\9���Tǰs�݉��1��~��у��s�	Z��L.�@f��̳���*a�f�˾�z���@��~y�����7�s��� �+�mt�sk�$�CD�?�y�=qr�\�F8��1�:oĂ�%�&��{S[ٜw|��7Af��|d�2��j9�+��5�լ������<K�ܶV�9>c�=��|P�)BK;S��^��}dB�(]������T헅��@�Є�@����OfN�S(��Ṁ��p-U�֏�H��R'Ѹ�K�0IG!�q�A�J�ky=0(),*@fy2Txʹ�[S@�Z���B�N�Plʨ}5����6�����O�6�&�`L'�9����M�[j��9�9��}��G�k|zFյ~�P�g�9�ul�(�KtmW@�6�����;���Hj�ãbP'5xɘ��iCYr�eu��M�����1S㒎�6Q����ؾ��=3h����+/D��R*e�~��K�]���"�@g��Ⓗ6{%i�s��.�6�e�%@�X��% �u>�d�\�����딉�ω��'p�P�[�G��*ݑ��<�@��al��в%�<�U�wfy�����:e,��:����)���3@�[U3��F<Z�9E]�B���)��i�Mn��򎖪�fƢ�����4/���-�5<ʗ�a��עZ��h�=����ϰ�����d-�Z5`����,�H�e��/���?8��xf�n"�R ��k��C.7<ñ��)���zb��G�\-b�c�3�9I��@���9�U؟< "��v��/fѸ�v9�q�?�0��vO�P�eh� >Eg��(,������$k�d������K�L!X"8O��n�Kn������Jdz��|L`�N6r�[]�m�mEm@-���KA��mp� �a�拎y�Ao�j5D}*�Zy�m jC��CeaM�J�B�ʠ�B�L+}ŬwE�;����rz������;
����a��R�|u;���I[Y��g��`=�vf�7���joӁ�f,G�x���*��f��9Cr�:�����mz�GL��A}M5��jSӔ������!���;S����Ԑ"���%E�� G��a�R�1��-��~�q�C؅fwFSZ=V0�k V��=��(7_�.K�����>a
�HL����jՂ��k}[ ��Fldsǁ��񳌶��L���֑;��� 'V	.�m�^���&���d6m�T>_Հ�����l�*�4x����7���2)�)c�r���:˅y<`~��u���\(U��2�*�^�-�l�$D6����/{���HQ3�}�YQ���h6���3���7�/6d�]��Mn��(�5��K��01�?f?��3T����N�b�at���>�7��VуnՏ�E�a��T�J2MR=��5j"���G�(E/��\9��]���4���I��(=@�!�ڑ/��C�T����	�1`�A�DY�+)�[/��fw8z�(I�q�a_1���2y����c���5Q&i�pnn�Hv�������=����"yy�M��Z�=@��L��6�Q�z�L�)�Z�O6��]�����l��r��YmCa�*�j�{�ӭ_�t��i�býf�ʥ-�(e��MrC��<��{�"D����UO���}ug�����Z 
E��]�I�H,c{��@ 9��Z�cX����՝pߛ���&�c,��&az�M4,Dl���q1{T�8�8�1�j�"����1��	H�
��-%�XD���XE�ˮڤ���|��.d����F��)����>��}����eM��&o��dfȾ�`<�V��K�ݹE�7`��#��B5<�A	~�Ǵ)�B"�~���*�^cg�,e�'>����w��$,�z�[�JIs	��}/��a q>+)W8����E�0J쟽쿯�]8>�y|�}�y�<����l�B�S=�./�<��?���b�a���1�#�F��V\-p>:��/�HTW��E�h�� K�7Z�S�:�����J����s�k@<�V����@�~��� A3������������ �^��I��ʨ�J�Pn�S�&�ک�/A4Q���uŇ��i�J�wH��)@h.bOt��t�&����Xy��[l!���R�+�$�ipvp��	:*�pE>�ހ�p��#���S�-ۭ��܌<�])�/���y���K#Ȏf�}��R�����Wt���l��~т�?���4�Gr��|�0���_�����~:���t���i7����a���8c�D����O��%j��_�d�E��iJpUG�u�K� c(�OHy��j��>1"�eӔ�wn��m}x|����,�V!��1B�G=�����h�dTs��JX���Ub��� р���H/���p ����O���R)���0����U�2�$bE��WK���^��4^�-�ת��U$CS?���Z��t�td�>�ʡ�o40��I�x�`CN�̜��������0�1i�
�i�q�g��&~ũ�q��,iG3��  ���A�r���ᚅ�i]�B��b�����Y&�K�����t��~K�"�2�x�(UY`�׈���T�1�}nB�e�Y%��󹩅ܶ�xq�[���K ��H�Ic�@��7���1D�׷N�e�8��9g�Iv,t���2��ێ������a�F�J"N# ��)�֫��[q^�q�j �G�% ��F88Y�(����1�%���3��.̢H�a�m�mz�dE�^ f<�c�����?�i&Er2P���99��(⸴�0i-����4i2hHu��L/�B���y6��_Yk�g���@�}2�$�����T�����h ��A�]|��,.��� ��5��T�/|u�O6ZV6f�ز̕��xM�%�.ޗ��ݖT񳾉�PN��>�Q�B��L�:��6������\�/��(���;t�Wъ����ꕗ��[�rh�b�9�̟U]�o�ԇS���!��HG���[ �<��$$��DV�����Ye 8q���t`pV�m-z5-� �a�|�T�֙4f�����O3.��#�&��=G��cMZy�x���	�G�����:n
��%oPi	;ߘb� ��O㚼��L��sH��(�btVk��I���o�t�*s�0p��'�z҃'���P�o�m����4�nʭ�U�e�툨�����s��}�|�qce�9DT%��̘ȯ�͚�q�����A]��%�M�M^���Z����3�� ���G��bM΄r�Av@*����14��Z��⁠i0-��k� lA����p��5(�����6�N��!�J>�e�Db[�43Z9&�sD� �/E ru�n�Ȉ՚����P�vt��$KST�00���y���ڙ���iw4�i��>D��nI����7	��3]}M���)
�'���w�v����&������0���OB�C�w��sn�Ph��3�N�թ'��SW��+h�vEl}�ED���J��I��p� L�[1�j���g�c*�����2k^��23��zi¹K�A�U�A
4�� ��E���B�$�^r��M�ehA��?���نT�
�S�}�I�bw�w��=��eX"�uU��@�~�y���_2ح�v�d��f�ﲩ�s9�a�7��Jk=��� rت��c݂3��=.Oz��A�3��f�~O�uB`F���ѦY;�^H�W�k�zD�h�3둍
qט:rN��N�ڸ�X(�?d�&�b� ��/ԮK�ϭ}T���C�e�JgV���tbä�Xi��_;�j1�^͜���2���Ê�
*d��O�-�6�xpq9�{�5��7{`֬DHg��ath��a�z��'��E2����mX��1�r� X�P	���vd=��2�x|��$�#��Ӕ���T��w�qɼ&�16��HKʂ2�64�Ě�A*L%=�@]^lޗ��,�u��A��Ǖ�k��$������d<Բ��ѣ��g9WH�����Ay�5N��V/*P����:c�!�S���	��t��]!` �~��ǝ����&hs��
����<��]Dwc�~k'�W����4r.|�� w�z��}@�Q��[ɞZx��Y��k����ޠ���]����½�Q���!.E#�!,�y�빗&���8��;d�4�b�&����g���z@�Tϛ��u��)��I��w�ऋvK"�u��V��\R@r�CE�åMU'v�zt)���-T��~&=PY�^#�Ǚ�Qm&n���芠��@�@��iL��37�Ы��_��5���������3ݕ������6j�?TNU�r�CK�x;H��	�5��#�O�	㱡ѭ��o�{��LxNl�$t�M���� DC���P:�qH〆�;ΉC�Tp���zH��O�S��Bz��ks�{t��nh�`F�������Ϙ��6�Puf'���a=�t��ُ�C�����A�9Y���J8�9�����Qm�{O��R���{LV���ǻ�x�?ۧ��=����	k/	���z��g5�4�e�h���~�^����E��Q�m
��H9qf�L&��9��\`+l���sj��)68�߼胮��qf!E����@��D�ǹ��Y��2��	Ŷ��
tt
�ڂ�u<�x�����}9��M�����Ļ�����<�u
YR�$��R�3f(>�|�y-��y�5��(�%C�������ÐHZx<��p���� ٺ���䶻�ڲꊮ����u��lCU��ʸ���! U�1zU��|��H�@���.��hG*�5�q��N�/�ҽ�9�x�����}g[����,�	L������I�˗r��a��tsU��2r�p���eHI�*a.�X����%����E��P�(��9rx.�� #�}��(:�b8R�%j���4>���NoT�� �Uh��ܹ�@��/\��}�E�?�Q9��=M���A@Ju��%0�I�o�%���+󹉰�.��p*K.�ͽ��%ժG
���}|��z��5L�/��~�3�04��-�K#S�d=F��L<����v���,��]�vo�	��C�`!����P΍����?e�ʾ��s��s>���8W,��	�.mp9�`D�����Řm`Ahe�7�ս�m݊leN;��I�?E��P�ܛN������.�\]��q����7�9ԒG��WH���j[Ȧ"٫@����[o=�O�ke��5y��Xr'�ٹ��S�����asL��YTvNx��N���6��.��.�|�֊�%j�I�K���.B��`��6J̅�_�����Nն*��;�V�p=��d�n�*$��Cx���⊎ޗ�E_E<v��W�Z�L%{vi	5�P|CW���LK�*I�$����뿶�N4��IJMi@�Y�SgH�݉��X �"�V���Cs`|�����QD3�La�j��v������ ��T-�	�$�/���$�<S�����Gy]%�+��,̂��?�2�$�dԖ�<��,��h8�;�?�Ӹ�+W�s{��&��~��u��cX����O0\��<䢔�d۩�p����F�Q�ڵG�0}%{�s�����_���FA��>$Eh�}�l*�/�O��lNmZ���)0G̋⹌��=�}�K�˫[��Eғ\�������|��-(�����3J����^Y���-�Gz�y�w�+V�w�)p�4v��Q1�!���(�ч�~{������(_���`�R�s�/bs�]���"<��*�L�W[�c)ۧ�w�'��*��p�9z���f���2*�^�vf�K�a9�b��~ޘ�X�,��k-m�ޟ�4wK(0�S��d8z�t�<���&"���s��W)/W��!6�G��ԓ�u��Ͻ�D��y.�z
5����P��ʧ�^�h_�o&c$��)�!����U�ߪ��>������ ��p���r�`݉�C�S������XͿ2�ZW`C�2D�)k�;��;Ͷ����mIF`8��3��E$� є�. �Nl�Ү�U�fB�ђ����xQ:e��uwA��tp�y93ǽq�|*���P�d��$=�
���R&_/�Է��-�]�K�Q�#���{柩���*7�}�$��r���"��̯�t��P�v/g�6z�K������/W�5i"�t&�vh�ِ��$�= M.e.���t<CS�*{j�9�𺧺�C��ӿQ2�����b��E�5C8Z�X���,���G����5>o逦_~�@��7�N�t���!yoڦB�r6O�5�,�	Y�YdPh�d-q�T,��Rh=��c��J���u�ͣ=<m'���N�z����)]I�>t������a��$5���L݌!Sl	�JkH�f�؁�z;�@5.ڇ6o�l{� QW;��~囘)B�*]����C/D����ɟ�'�%v�R��;�`���z+	�9�6�r��^<�p��7������IP��Ǌ�J*�B�C���52�+�W�U�V�~R/}wF�P�s�>�K�c�J-���۟Cw�	�E_w{�	����_�7����R����O$��~���
���`�����A��r."�zS�د:۠�����8�(!������נ+͖a���B�T�5³�2$������0a5[m��i��U12���<ߗ��7%Zo�L6Q�Z-v���������T4%Ճ�b$B�'3B)�QՓL��=:��g>x�^(,3e��
s�����Q1��X�"��nC��������X��C,�V!j[�s�I�����ud]/�����L��E������
�mNu!ҦgX�̦O���ހ;R��(�>YH����h��LY��²y\�
�^��ڟ�����6�W**0��w�"�X6\�v�</�},N����**]k⭐�u� nǬ��[�<MVؐt�?�I�׶c�5M�?��Y(Z��H�����O�D��t���.x�wm��¢r8� �;�P��*�<q[<�u�T�6b|n�F� ��e4[M(a[���_2 �ɴ��������2$��Q��cr�|.�8��3�&���ql��z��-?iª�0��֚�	u�<\(DZU�n�~o+ؐ�e�=Fpu������ט,g��U��`�g#Jh�q���R<>g��J-��6�`��L�Ǹ�*�C@7y]��f�W	ɏ6[���Cw��Ѿ�(K ��X������R5Ou��I�~�0;6ӫL{X�>Y#�FYg���h���(�l��X%-�������w`�i�.������K����[�p�(��+���V�=��݂t�
�����_�-E�~���x]���y��K�dkd�I�ֻ�_-th1�9���Ue4�4O�g��?jˀ#�����)U#o�jaŷYlb6������P�������`47�[�e��$X�����m�z?FB�3���y�JP�\/Z��l_������/򖣶�4�xv�O6�^dB<&�1�o�6�	���Q�0]I0u 9˜��]�]��Y@���H�yZ[��{z�W���Rs ^�,�Y�2N�{T�z�G����4�|�����[�++�KY�t����T�T;��A**ө}�F�b�<]2;�q7p%��j~�ڟ�)�!�4��@�S,^�h��ӧr&0 ����&T~���O7��I�������:��J���!>����8b�NK7'ID��<o�,��8?�h퇁�׌9{L����k���s1�O�燮K��n%��'i��R3��"w"`�x��f6b����̴.h@�dN*��2�����O�� ��Zl^`���)���B����f�FS�mu�-Ӣ�-o$H
Y�^w�G�(����<5B��^��,6� S1�s���(Ȥ�`���ʮ��5|��Ҡ�^{�����n�2��r2��^�w��;<��$���ٓg�?�X&�[j�1V]w �4�9^��0�K�-�%qM`�Cs2�s�<���U�?9:2��G���R*���C�����bM����J�wU����q��^}*��qJ�k:�jH��Cd�� T�����ꪃB���z���ia�֟��)�(ݭ�br�-t��T��D�e�и����^6
�G��.��č�*���Z��<{�~C'���G=����;�
���o��D@�ڽ^���U�i���g�b̶��a͎RTT��ZPm�}�4�6�@��60���qV4�����Ɏשpq��������K��k2�E���M���i<X�#i6�_�ş96's6���_Chdo�
[�ʦ���xj�N�N�,Ԏ���R�pk2�-�p��b�����)�9޳����D�1����e|��|7Y�= K����'cd�0^���(�M��y��V	2���Ӊ��ܓt�H�忄�}��D��w��n\�}M�2:*�
����#�������u�4|�`��c9v[����q[ZQ�5a��T�R���e�b�-y�\�ҝ��$�P��. ���Q)0C�?V��)΍*ϯ����Z��ɞ`X�z�,z��4`Q;5�����W��-�dz�zE��
w��.kK��t�"��䦭XN�>���u�(
���`��w�)�/凕�����)����V$Mທ������-��Z�M�M��3JѤ_��.���x�ó9:
na��Q��U΀�Q�F���v���*��ͷ%jC�NV<2��`�t�����Zkhg�B��.mb�����,`B�g�*�ԓ*���:���AN��fw��s�R��$��b8���$���!�`��J\��{X_���''@}Y�^wSX7���{=y�Y��\_͌]����h��n�]>#%W���%Q��M�ߴ5�� -6��e"3$�sB�h߳G#�>$)Aat�� �foBy ��jy���HL��%^Ot�����U*���P��2KS� �9*��[Q�[��W	l���c�i~�{�����h�Dٟk�!R���L��_�����&����>Y�QK?��b�ld!)2�B��0Um�1L�8�l�pFj���n��%����/T�����V����e�o��3|�[P�� ҁ�5U/+�ml��}ݶ�����^�%������DU�z�d@;0�����^
�m�'��C;���O�i�Kn�ӱy]�ޤ5]�$GɠZ����k�E~�<1��,>��浱)x�c����~�*տ��R��D)���m.�wX�=-��7���0����ϗ�`=������n$���	�7��Y1�]�e.t>guq�������?|خW�vNI0�&�@������򿦛�Y�JȾb[������XS�������Ͻ�B�1������m�F��T�E�8��m�9��J�eL��s��HDҬe���ܰ�{c76\~�®H6����X;%g(U�T�P�F����ĿkM�~�uÊ�OOD�]�g?`W�*0c
5��."�
Y�CH��ul�s�Q�i��>��K�#��{�e���:�ZNu�0-�ߣ]��Ht-�K�F01�Z�tF�1�"����6��17� a�s�L�IP�H�cxu ��PӲiX#�p��`@�T�� k�0T��	���U�W)�*D��	�bU���-��Ǐ+ɺ�;�C�&��h���^	��t��|�D���������鬭$�ed�������B�2��S�e	���8���8�~CZ�d�Y!BwR�z��d��\�7���Ax�Q�v1F�n��w��R����zNK	}��1Ʋ�VJ���"��������s0Q��lh���g�	ހ9��*��N�ʱs^�S��R+�'SƝGջ��>�)���hl���V���q�A��r���MjCA�ѽ�
:��C[�D�L��15�H�̽�)� 0�IW�vߊ˥�F��]���rua���P�ʐdv��%��j���g8pd�W!�mTU/U� )��k�2��TL����1n�@S�i�a��B�tTg���k`�=��Pgf�&�2" J��R�P'Gi��"��{���X>��s�J�0�K�L<(γ0��-���(��M�d˵êVHd�*K	�"μO���.����/���ύ���ň���Q���/�r$�� �I�-����ss�2� 	�gsN�t�F�����$ꮔ�~Ww��hF�s*t�~2�4���S6�`o��mC綻Y��v;�J5tVC���:~Jf�k.�#��.~d�\ �Z,/��|b�Z��'�?0�d�g+���D��R���ƭ�:D��I��W���n��(�9�6��>�����&�y�VO�!��\�md=Ѽ�o�hM\�ZJ��F���ԡ♌U�A�Q@��_�?�W[���L����%c��ϕKZH�E>���`�eU�Ǚ|�+�,O~����Ly��ŕ��Kh�:[�� �bb5&��b�+�MF'M]������Ec���c�!1�����G�I�1G�h���&&����7�qB��e���A���^�#��>a�u��0AVyG��'^�x����˼Ǭ�qg~���b���S�**��>����oi��g�����n�y�x}�,n��TRlF�]Ȓ�Һ���zہ����uқ�`s�o��f������0����oˡfg)WQ
�jǿRW������r��s���+#Z��ؼ*�3��1i��q�b��"��(�9yfi�����I[�"H$��>�PX�y�ԛM���er_�d�J9S�jL��¼^���~3t��p�tΙ ���}O*� =��덝z�M�����wX��0���0${��>��OΛ�8
g�+��W�%[���������o�{=/�{7U�|�pUִ?�cqR%n�0���d|�	����K�m-�F9%�5q!�YPכz�1_tQ�
#S�ɔ�S~ɻ/Ǯ�"���WT�$�D��N�H)0���|�4DͨR�Yg:jFn�
���hݍ,�&�T0K�rdG�קx��w��Y����0�����"�r��=�|���R��[:���da�X-e�ې��h?�ۆ��J��.e<���d��kC��o�0�n�cBU,�j�^{���ֽ��{r��x�6 ����	J^
�rZ&L�};���w>W�ٰ�H����M�	ED/r-:2��XrVσ�ET���%X�Q �v�&`4t� >2yf�i_���"<G!��mU{�*w�Pm���G�O�U�u{�U��%��Pdnd=�m�����/x��S�@��D �-V���<B�Ȃr���1���	A�+�{?��'s�f��_�=t��Ӷ�"�.�U1�s�a�O_g�d f5�CmL�Ҥ�`l��Z'���u�&0C��x�Z=s�Λ�b�Ct��r�K�)ޅL�1�J%v���O�#�b����1�f�ښo�Eg�Iya�_�YK����&�P���Kk��bi����n�K9e��K�Ӈ�0>��L[�<�?p�x�Q(�"����YA�{����g��}^MkT-�ֿ2��p0�sX)Sk?��s.�0��^�Ÿ==�%�z )��,`��N�C1�>?��0�y<�%�$T�t��>����Z0�VWpJ^g(�J�0�������D1��"^�nʜ5?6�)��T��e�����T���D�� 1�������O�Be��\�|m�3f�mY�9"�*�2��(���[#�c����5e���-�"��W�P^�� �`k�nP}������b�;�Z���B�]ET��������4?�"����ù��ȡO.p������/�#Dl;�]�3�O&��r�Ă�E�/��Oz�/���E��Vm�Ҳ��������_�fS!�`�[;�8��__���HT®�/6�t�$F�/;ww&`�r�m��Y�>��<��j���ܳ�%�z��˺Fn3�O-��\W����i�����P} �{e��w"T^� }P��P��ȸ�.�1�3��Z#e9��
��Ɉ��y<��tօոVl��O�m�'��|t�Nqh��[h�i�Q�`:E/!�����L�r�I5��>��L���(x����:���hx����!�x$5Rp��Ш������0�Ɵ�u�dI���g�q�!ct�z!XI�U�����Շ�#�@��ӛ<4M"�+����@u?�ۿ�Z�9/�7�
l(��Z���S�c�m�J��ߟ�7�o�U��m2�9��t��g|:ƽ�<�� j��"�f��Kr����� ���CG�Ǧ������9�7�S-f�g6 IG��<��N,������&||��k���"����Ǭ(@��yBFr�MM�����M�1�)a��X��L*��#����.��k�~�k6%z*�
���}ԅ)Xd�\�H?��Iu��Us��CuW��G�Bm��j`r�F���M���!�bD,��P7@x��P�����5Ȫ����0=/Tv}�-8����b�(,�����f1�Q oVj��6X�����0�
�+Z���Ȋ���ﾖr=�Sy����1n�$驘�+��¬}�FNʸ�2�I{oyaQw�qbc�h���{��@��**�܈8t��*us!uu�!�W��}��~��W�.�`�*v�[�fy�N�6�������[��9?h��tHv��Bb&��>�:|����	�3) �Xv�k��0�/ݬ<|c���4�&�X9�,.ΧM����0��'ڃ��[�{Z��ÍD�Z�a�+�����rwlR���]7����xr�ܾ����?^��메�5��#�������]Q��{<m��kǔR=)���Y;59�r_�UUM�J��ſ��:�f�����G�J$�u�P��B��xq��]���\�u��^�������s����u�����X�����S��� d�^��4�,��m������'
���i�D�T�����n��g��j`�ɼ�,D�x�� ���ݧCD�;��@T+��Ѥl� �]/ta7X� �0,�D�D�
$Z|n�KBL7ƊB,���yò�t[����{�[����l��W�]"�����&���'��]����	�}��*$^�tU��;B������`�p/A�>%����r꓉�!TMr,�VeD�ɠb��B�=����:'0�B���E�$C5V���]�u���{5/D��'�
�x4���\e����p�k��
����vx"��O��Rbg�bZ�v���W�c[G'�-jTHp�P%�]�p��7�����y��̪N���=m�a����B����'� �2d�7��8%�a�.��XQ��%�c�a/ġ��(���bz/��i	��ͨ��WZǕR7�z����g(���g5���*9Sܼy��U����}]��b��2㽩���!C��G�ir	�<)X��w�g>��3���egq��f�t�՛�eڄ�Jk��a�LO�q �8�=�D��s��$� ��y�Cվ��Y��!M�d���M�y�C;<
���S�9y�?o��Go�� �W��:N6���ѢR�[�Kŧ���8g��N�
a�B��K<^���eu���5���5b<��}E`ʈ�T��1k�M$^|�*�6�t#"H��t��ߙ�f�vn�J��zE⇲�s�NR�>|�h7�X�å<r �A8��~^�ƣ�~�{� �V!J��{_�׬TG�9f{qh����Q�[{Od�x=��ě������F����e�f���OK��@?:��LQ��xN��z40�~�:�B�2�� ���O�:�z����T�l�Y3z��=шxN�"�[.��5����5m��V���JccS��i]J鍌�)��֟T�i&X�!� �D<���W�pJ�|��"v����:��Ds�?Yѥ��>X��U��3�u�S:�z*@]㴅���o�g�����毀�"�!M��^L���a�?PX�mf+LBfb�u:?�M`��+p��� ��W��	�W��b���� �M���Mz�$1�v��H�}�y���I��է�4՞'�<�[7w��*�����i�^�%c�3��w|y$�7�@�?��(�z���� 
B�5%�ka�*%����빵�e(��J���3.���~v}�ÊƯw�O�)x/����C�Mԓ��-�O�ӽH��s��,)�m{on�S��g��zG����
���s9i�M�G8���y-2 �PN���P�(��0j�(3�����C�K�j7VJ�Y���+S���G�`�{h
�w�r_����)�&���پh�D+�>;�힛;��V��aTƳ!	H����Вk]�S���oX�U�ϵ>�y,��.�8 `�o��?v
> ��{R����op�� '�a%�7�_�{s���EZ���UMA��� E�N[��<�:o��p�v�:������7 y�")�m�I��4Z�v�*N���,����~W�ȹ[@�Ol4����8�35�J�3�߸M�c�UFj���sR��qV�����~*���E�;aU�z,L��_xm��U^bǿzh��0��\���Ŋ�~Dj�K�Q!�e�t��Y �?���)�u������|�iZ����u��/x�3	%6̶��5Z;5�҈zS22޾�rh��~�!RM߫*;�n�`H`��n�siP�%�-ɬ91|u����`- �g#o��5������,u�#'�5���fס�77>��攃����eA3;��(�sޒ��)`}N��5��'�����^f����:zM�����B�;%=��6P��3�x)a���|�]���_����rti�~��CJ�IQ�u����b>�Z <��GIpd"J���=�U�Z���Պ3Ͼ8�A��(��^g"��W�����wA �V�p �dyP�l�p�߻�S:1.؞�]�M� �$k��{x��M6i*��S�F������p�Ay��ܮ%�6�GBu�N2r���������t|�r�~[P8hL��<&�*Z6M� ��rm$�Z���9a� J4QB���?<2�>��}:�p���.�7||��m�ҤR�D��L��q�D%Zڏtވ�ԕ�Ue�f?�H�YyvW,W�"�'Ϫ�	�`.��&*v�v�4)�]�H�Uqd{s+��pi#�(��� �>	W�=�ev9t�-\������m4]�X��^#�i�'E�^���T$����Ƹ��rnNߟ+�[������2�z���^!e���I������{2��Ns�zZ=���l�^�MU��(��'��h������s��#U�A}��,�U�_0~� �R�!�J�ǖnn�7��{����H�o�/J���̚Fq?���ϼ����/+�N �x�P:ȳ���,��2�^��D�*��d�����4�2.�+��b����GeWTD���Oc��^����VgW�8���gP�����I��d��� �O�8�)��?�pm�7�D ~=�� dA�ԏfwD]�Ae�
���;c3�7;C��G�7_�O�	�Fi�`��^��r6���u�
���֔�X��x�F\���L����E��hӽ�)�����$��I���4)+6�Rn']Y�W�1䢢��F
T*������u��({	֕u�>���@Ń��j{�8� �K��W`YA�<u_�ט>���[t^��,:R8d��+����'���#�C��Ԃ$\j&W-�o�
:=�� .��
�i�YC�S{�1ɪ�!Ӿ�����o9<ѵL��o�k]y��� D�-P�=R��<}e.	����Y�dH����d:)zly�	84҈��9D�9�M��L���|��;����~2 ��LK������OoKe۟���ai�DFiW�Ӓ��z�ܒ�b�� �Œ�/�&���Z��	ɞHS{���['�.�W\*B'���JDs��&�s�87(��Z?����Ԑ��D��i>��[][�`�!�j�M�l.�2U���_Y0D�6��K��B,FUˍ% i\��c��;���+�����A�K��N_���1$�?�0���h�A�I��䷻��x�e��@[T��Ex7��ɬ\��-	"Bv\_���[��2VS�� T���TZt�!�!�~�J�K8ۙ��W���vV:^|��,�z$��W�wՉ�IfK���U�����v�(�G�Dz~�����=Z�������Ғ��qKO=K|:4�A���Q��D�tlS䀿��H ��d�R=fQ�c��,�x�[�����t���/V�3+=b][U�������m3����S�,)�J��+c@�b{�iQqf��¤Vd�yfJ�Bn��B���ִ�6"'�ӈ�`\3�]N�âz�a,��~��� .:q0>���k2�l"3�*~�S��iD� oy+�'��T3ڶ`��q�D��f�	�LZT�)>����q�M�w�"ǉߔޙ.F����1�A�Z��ضoƁ�������c|�����`e����)p	��� ���v�-H����c�\"��wdB�c#v�d�6S��HJ�?��F�3M rL�@��z9kg��k7�����/�����_&5I��V��nb�mwy
����-�kRM~
���⨝)�\����(���׼3�r@[�΁����8��?�@bL<�AR7���NO`m�h{�A2͆�­�M�bP��~�#q���KR3ۄ6��@�7����gV�E�x�L���8I��L�i��|������C�@⤀*�8xN(Ii�œ�!������3s�U�R�ؘ�ݠ�O���DS90���ȘV�uJn���Iu��T�x�2"�L�S^�ы6թ���u�J��-:�L���D��Ļ����F�LE4�P�?�n>�G����,�K�~�2�t����V4�&3���02���1�33���~9ؾ�/����@m���`
;S�V4�K�T�"}� �\I�Xx�
m�t8���uJ"d��0�]k���Cy&<�O ̴�4�ض)�Ѝ�~���BZ�y���q�,X��߫����OV�QR�_���b�(iݗe'x�z�����W�B��'V�&̧2�o6���Wg����#�3���O��p�t��&$���q��mS��c1�ح�+���pY�P�%��
�X�P���6�q!��5���dB�ф8_���8��"d��n�,dcl��8^�kN#xp�[K쀹��s%U�/6�:��^A���>R�]�_[�79�����Ք���r\eʜ	@5��i�Wc��	�n�Yw��rĻ�������J���`�ʖ[���w����P<f�n��a�G�oS�:0��n�˛Y�fX�=��:ԑ+'n},���;��9a�"I������D�v�����:��JA˹\f��VDȏ�٫�O0.g��W4�S�I+�Γ�u�\_�s7[r��k�{�?	����ow�*:Q��3��~�N3Y�lKGq�
���1-�H�}5q�ۓ)ht�u`��]���'j�;*Ծ��n���4�ݤps��H���^�dF�I��[��/��A`�!�W����J�ʺ���&x�7vK�����!��^�?�.��{G�V�R�Li޹ĳ?vrL�5]�ܑ״y׃ls�d��Z9ǯ�V�0]G/����4��au��*��7=v���D�Z���>�/���719h��S~*�9y�S��L��M��B�wz=�N�T��\|���W�z&y�	��7nT��R-����>��u{����)�&���?&M��3��:���OO�>�2���B=�UA6���^o������EN�.���5@�L��+%9e�.�F�(�����^f�c���z,��l4��("�~R�W��g�p�Ά���T'\���B6��z������Ÿ�ؐ����]�z��mh�UWT���AR�M�"�5�}�5��T8o.�D�Xߘ���Yx���Ng�%��2 �2��N Ϡ����wk+��-��Onf�&��Gm{a�JB�JJ�'���Α�?���N�ł�+1��XG����v U;W.|͑�� ��֩-� ���ԃ��F�����ֲ~���vL�rM�h�n�=�^\���RT������$ι�e�g�A��۠A~���T�9�b�\�[?
�y2q��m3�+?^s��T�`Bx6�l�{�F��$� ��R���p�o��	�!�L�(\'E�탣%�V�����0p�r��YY�*��!
��4[��}���z���j��!���ײM$��7�Kj�� fF/�@��k��@|�ڭ��	Ү,�p߄?$�>-�WEq�0���"�w�"$���,7�����_��\�?IEe�����O �79�D��wp�Vy�H�U��?�Mg'�x�T3{�{:�D��s�%Y�~�sBj�ہ¥~̲ˠ��=�,3$a��x����{�҈�*w�C�����FT��Q}�o�Q����h��Yʴ�gW���
:ydj��F��}�� O�0�;��Rg�Է����b������7Ё  �d�!A�=�Tɳ��e�U��� �>%c�(x�-��8���v���0h��<����Ⱥ��k\�����"G��H�oU;���W��(͙�G4ȷ�����
�q5*��
\o�J^y[L���c�(���m>� �>��0�����ԛ3#��,6��Ǟ��g�_���=p��s�c0]�{���
zV9M'p�QH��w��)�ƃ�|���D��f�`,b�F����W��p]`����N���҆�8U�"�'����_QI�X/�ͣA���m�)o��LH#�Mt�Tl��D#�t�1�!���:>mD��q��77V�
��;�������4s*keV������o�v�/�fNN:r�(k���~@x/6����`�1$�>��_��t~�u��ry,��~v�q�8�4�f��'{jN������p���q8O�܏&b�p^c��/)h�h��2���&��G��.e4\�6�`ꈝH�Zx�e�M��<A�T�7�&�%̯�3�u�ZΨ.��%Dc��$|)ؐ��,�U�� '��M�ק��/. 󶛌/B)�:���X��������92/�:+G�Ƶ�ߜ'S��}�;b�A��B���������.��L˵(%ﳕ*�}1�y�>���M�k��!k/>�����A�r�T]]vA"*�%�K��4�sc�ݣĜ��Yۭ��Q��x�n��|�����Sk�a�]e"�'������ξ}�(�/���tﭬ���d�8Zҫ���a�J&�XQ.	�܂������V��(���e�����+����$I.r0�R	l��A3*|�� Lx�?�����i���0�Z+��/�)��]#F�i7�͒��s�X�u'zG'�Y�N�)�H#�T?K��1���V�������I3�h�ȏ���):�F�l�ί��J�d���/#�6m�/	r�uo��m�H����i#W�mi�$�mT�����o��ame�o-e�ݤ��?i/��@����> ��rݕ�$�A���|ab��=�- �@����W�zQ(���1�,�����/����@�}zP�I/��^��c6Ʈ�����ȿ���J�v?@Ő��N��H���M d��ƨ���`/���Oa���;{8"3k����V��
Y���PZ&tCT�n��i�B)D�������V� �OB����i`��e-��^ry��|`MY���T�)�e�����xqY&��
��Ή��
�j�I[��(*��3ʾ��5�vx�zC���k�3��=�fV6�<hۡq.w���qm�!?�`�6�j��quoZ6�^
v��!n�Դz�6��b首G�Ɓ�?]����U�-
�Ht䙙��!��`�[�a����2]Z�ɁbW)���ph�m|g,���;p\^���8���y��#n�u�vv�Lzv��\5�|;�O|2�����`�f	&���.k�B~�s2U�c�;��� �z���� zZ��M�H����3��8hz:�e<#D��m���Y,gõs��[/f7	�>���˫R�؛��PN�˵�����t�c�]Т��ĖL����h��E�0=��r��2R}f!�H@E"5�K` �ࡑ�{Z�Q��WB=d.��Y�o�K���1M�� @�\ ?6��R׮a���⋦>�{��D3%��v��������F{��7��2<q� �z�1/7:\�sr�4�n� 18:����.#��BE_^���쵩!Jۗ�.9�Em�+��9ۆUj���w�ݑ ����x�>�G���>�
Ӱ��wD�	G�D �ڎx�Z��RS��~���-����Q �*8�Zd����fWS,Sl��N&�z�*t��5��%��k�O��}�4�hpe��Đ�CHO�	���V�@�Sj?�6�.�|�)��#$�Yڗ5�I�0����o�*#O^��0��X�� +�����&qM(l����R����,��S�K�}�{�|O[]j+�����\=P�H�x�-�'Bx�v�>v�z,��z�f���iN�(=���Yy�u�l�r"zji<��)Oֵ˺����S�v$���w�J@�����,�DEn ���88fDԐ����m _��g=�|D�K��N�Ba�U�F��!��i��7H�u1_ѯ�<4B>�~V�85�����p���&,��B�B�;O�Lm��},:j��-sP�3v��e��%�DL]Z���q���k��6>ʅu51W�-�l`�:}ǯ�*=�k��^��;�+V�F����`�_���`P�����T^P�l�m=hMFⶵ-�EM��]���zf��L�+%>KY��(�5�(8�F��d�O��[�J��t������'hѾ`��>���Wi�S���x1���ōRn�M�JaK]W���>�7�#�s(�>ņ��f	����2�����)딬��_�%�ZѰ=�%NJ'��/gCǾ�?�S`��j#b�hw�-T��zm-��y��,�#d�X뜯�&����@ۼrlE	�G��<LmO�()L�v��ǀ��Y���pŷ'��(�w���$�[�`���E���3�=��튒o��}8���Ԋ�T:@)?�٨����'�RX���qR*�?m'� ��1��	.?��>�Hag��Ո&�
`�{�>o�f|*�0l"����q��ڰ��4����F�`�_�Q]�~F���I���xEÞ��2�Nf�u��@$�Pg�7��Hpa�ԮTE�������)b�'F�j��_�`,�Z���:���◅DC{,��;I���K�HV�t��E�$)RD��(c`�|�X\�h^Ū�G��d���Xe�����Ey�a�&�I�=b��&� �����Me��RS����0ڰ��1� ,��SpZ3\3<��
�P�-�<XHx���m� �7N1߉�Yg����V퇛D��1ѡ�h�\	�]���+n�+vhx(�#�������!�&I��~cj8�;/�̆�@C�G^O?�_D�	���C5���Zڢ�l%V�|�yN�����.��wq�4�PK">����p��/�0��X�}�|n��A�0�=����|�`��>�)�"��>�_>t
�i>p��y�����H��d�d�E)�|9w:(]n�ނj����΁3Xvg4�e����� �-�U������Y7=P_@]IB��E)���F�����P�*����H�.���c6G���fI��4���ap�>}^]�n.
Y���c��C�~��!�8�Gr\}8p�5-v[^�ߵ�+���}��ojH͔Y�+�����{����ŭ@1����D{zJ��>�,i*�@	r_嚔<p��l������hq��%��Z$����$�[���gu>ĸP"q�a$�Wem�u�u��m��>��U ��:��AX5�4W��$�]L����3��ȇ'���h���L� �A�-�رWX����dk��&N�ZT��A�\6��x��	a��#0���G�me��*5xJP�`�D��34'5`��e�)����!o[��5�]�?e�q1-@{'��`:0�[�G)��t�<c|%,�4=���N�	o`
Z)M��VY2�$c�1U��TZZ���$|��a��V��.'Q�Pa#�:e�JW�LWM[�]u�$�B�v�3?�%K*�O������ż3Ix�.@�Pb�%���u�qBuҲRxK��ŷ����p�nAHr��"�o�0��	�[~����#u�ڼ�����N|j��R��m�(�v�k�����!��5�7��X�E�ߕzC�|�؇�i*O{r˵YՕϋ욖�?y��ޓ_B�ڌ}
"��ۅ:�!���>뎏Ms�@2b���K�rK��d|6v|	Ɋ�Vx�v��@�V�ʃ��lSz��+M�3-���#�-E;.N�hJ��&ߑ�ڲr�5.I<�����zh� %���/��,�
�:��[h�o�i"Yl
�/c������Ӷ�nS�G���n�
LP���~;I�@Z�y.m	���{a�\�g��uY;�NY�B�qh�6i������^��B���H}����U"�@4+�ގ���+�� U^
�n4��;�[��Ax�O+�"2e?����E�]��U�f)wh�ꎳ��jV�<.E+�ٿ!$2�P"{x8����?��zn�z�8t�������Kh�[ ��Q�e���������.��
m  0��(a��0+��5=C��Z=�9+?�B�OK��p��`]�sUE�\30�D�K���X��a�nR������3Z��X<
�3MR����S�����
^*5k9�=��kg�ʓn:��4|�M��/���#)��pd�H�ik�X�h ̈զ�b-T����*����ż����'v��M�mfډ��<X��φ�k�ێf	��N9a��s���{����1�;@׋5��aD�F��G�ԒH:D�-�{u}�G��>I���L;��2�Y�p�$���Պd?��b�d��9M)!��u����WV#�v	�4�����1A�4 ���x�[�R�M����t��9�}k��:������@�Ӈp9J�?Q��w)����N�#X����&��%���~EԖ������|���Hc ?[$��s*8��,/;Q�-6�ސ�)ѷTam��bJ���w�"L� �Y4�.G��W��oY�s��[��-�B2>��/}�xh*+(�!� 7s�Vs,���jͶ"��R���lw�3�2$R�C�/-�:��G[�]cM�ޕō9�4�`[��i�~|Y�����p�vs����|W�V�~�fB���w�%F2�C�>�N�+�;��;+�SxT���R[��$�̙O���6��OB3{�{���ļJ�^�cк�ژ��@��R
���nI�[g�Gs�B(��#����l�.��%R;Aen��$��j�Ii�V3��
R��h�\%���^����<�ͥ�g��Q��D�0¤>��j���?��S�ذ���n��ø�D�2Ӌ(�i{����#߃��Q�O������Z���
����nz%���Ӽ��_��v�.�R�j(����`6�V[WE�M��|_t��9o#�:x�)[�x|�`w�1���`�?h�b�il����e�f���ʊ�c���IYM���Q��f��x'1��fk(.&��Up���<�R�r	�鉎F��η��Msˢ5r�y�Z�v���������W�����T�8���������W\�4(�}��`�+,bi�>� ��;}A�QE���IG��A�S/��7�/�d|&���<I',�d�1?�e�
0q
^]�
�	���{�o�B!�J�\�t��h�@���<\����g��~��^q�H(�-�(�b�pJ��[$�g(�Z���g��Ib���)a�5<m�UM:�>���yL/p��ڥx�+��hd��1�R�LeZ �w�C >���/I%�22E�>ݽv��֐ݛ4/�A��s��B��,���&�=�51Lac'e	��$�v�c��˚Ԕ�k?�}0��2.�����:�D	�B�=��s`9��QT��?x���6ҙ�;�o�p���C��3�[�x��Z�����k�Å9En�C<���jc��Jû�`�c��a�\�R-�JH�� v�Q�j��2^
(�+'-��n�>��0tHh�E��ǎ:�m�ۖs�����"�8@��	�I�i�fv[�3�?�z�Wů9'�D9Ē����n������X�~4�	�c�Ei��yq����ie�7�ue�-8na�Oǹ��ev{L�t̨D|R������<��,�d�QM�DĎ��ʝ�;�MRU#���a����R�q�h%�J�/�0�l$^$�p\�(�W,?�_��i��r��p������2_|�s��u�����%Ϣʎ?��aH������K^�7�=��y��3�+Q<�F�Ty��)[I����t�a�<�K^����&�?��*�|I��_��RB�bַ+:tI�kn@$Y���	�%��/����Nȴ�M�ҫg�N�s������!�T���X&]�zlJ%b��	�G��=yM�2c�u����iÉ��"���M��0k����z���pD���y<�e�e�э���}wq�Ҩ�)�?h,�U;���׍̙���T+nUs)�4k?}���+�d��$�����F��.�#��^��G��)�P��t�~���4)<zN`�J���۔�^ID�	�==�Ҙ"���P@�n,��D+�6h 	����u*o@����D�SAj��Z��ϊ]�tCS�v&I3R�B����y��7��Gt�Fkڈg��cT��Ն�o^�b�_yNQ��/f�͎�CN�JEe槉9!�H.%����ǭ
�ZXL��-?�}�����d},/\gq����89R��rs�IdWA�<�f����;��w���Mډ���Elȭ#W^t0��y��II�#l!3q�2��;�b�ٽ���]�*��L�!�6�"�B�-0C*h+Г�ha�*�N�8v#N
�����0��lgK"\Կ�hoҴ:���r�)ɗ�of	ۺ�_\)��.ڃ�0�6k�����|6$�{��}�S��/U�8�[ƁL��ʋ�w���!���|�y�N�T����b�6Q$k�\w�_��w�KbƬ�9�9Iof�^�.�Ȳ?fЮ���q�	��I�m�y� ��<W��U�*�z��~%�0��ܐ�Qy!��ިQ[���z-��-� ����,�"�D��8�x5����ڲ�{�P�����
錐����2#��~��Br�g�1���׮W�q�բ�*����F$�=?/��a @
�?��������wD�5��L��V
��\�z���Y���Q�soN����A��>@�6�3���f)�x@ta����d�a(ғ9�Ox���`���$�}ߋ���0w����+ˮ��לLsd
7;lm�NU2}>�G�
���?����V�׎�{\�Y8��d�ЋE*�OM�ʃ슓�FW'���9-S�?�XN(���*�,�
D��
�=�s�f5��xvg�FAg��S9�p���j�#�C�5�U��~����>�o��;��N�s4�p��~>Y��N-p
���"/N����NKуj� 3m;����q6���G�2Lsi?�Y�Ab�D�� �W��qХK�)��a$�N�L�&����h����2 ��l�	%R&=��Cm�A��+�#�AR��r��k4JgYm`��o.UN����*�t~u�,A��D�O�b.~��߳�78��zM�������p�bA�{3X;x>��`���υ��O�V��*_�dV�PH�4&U^���N򬓿z����6�<b����f^�Y|7�5
;Y���W�=������d�r0�EW�}�S�Ɔ����e �$]��~o���!l�8Ξ���c�xg���b��jn.�Y��aW��F��Jz��S�q�,�Bo~���5�#k�%������h<k��=���֑��m=��9��ȱ>h�^*���n��]D���v�� ����}2�����f�#@]�*�C/`C�.���?]��0p��rRwo���f#)�,
�Z�	h��/o�C�� ����������^^��g��fv�P��0���dz׆���E��O�Զt(�yE�X�c�Bˬ�V:�%�
N��t�������t�y�bk������
��ـB����^�h9dz	��܃q�H��`�\\i�/��Jj0k�>�� ..�J:-��t��T��É�:�uܩ���Pf`~��~}�ƭ|ad�Id�T|̽^nێ�o�R���z���O7!��5� ��	�?ƽV2��25�l{پ7�mśB"Kk��N!z	��(�-l@��Q}\Wv������aY)������\,��1�1=�U~۪�w����tv[%@B�I%T"X�U)����.�q�����Q(m�#C?��r�`���>;�=��M����-�o��B�"����*蟝c��˅9Y��2�����Y����w6���I��`=Ǘp��^��F�BR5f�V�8����Nߏ�0�p�+Q�"%��{�,�F(�gu�T)򰽳L�Z,߶O���H�G�A ݡ��u$߉\aW�`���G�g3�2�R��ުTtGݫ�,����koC+2�Ř�����8�*t��x�匷�h��ܚl����Ɖ�潜c�Z��c�i= �Xe�]����#1����:�M�� f(R��WBL"�
����A�O�u��$5a�Y��R=������#l�!�p s�Zp�IS�ui�̈́�T�4Rǟ�����rN�B��fn�:Nq�qA]r5��N�����f�"�V���Z)�w摂�[_��B��uC�9K�ϫ���۸Aͥpl3E�D�$�T��I���K`	�1�Ύ����tY՘'>�u[��s"*�j	[��g���	z�Q�Pg0?��߿�ğ$"���m�y7N�cj��BB�?mL�L�A�E��#�3J�_�=a��zR:f��k��8�g��t�9C�7��-�N"/�u6{��O���؄?c��#IP��͟	��T]di��L� �x�̈́co�� �I�4��,K��U\'4���$woz����_���b�����)!F����>Ѩ�Mn �<�ӖyΥ&1c��U��������Z� n����ZY<0.�j���4l�yD��2�O#�L_��B��j&�']i��,�h�u�:PW��]f�_��=���z�ٱ��϶RS��~�Vq�Lq�1�@�ͻ2��j��l$�iN��&��:��! l`MZ�lR�y��S���ʢq�h��2'�y�U?J3�05 �ɼ��up�~���K.1�;�:�������u:���=���f�vNYd��=����|[���w�x�OS�i� /��+�=g-E �ue/hS�hɸKȬ�ݢ�$��O��XUXWv�Ե�h��"��c��{N^�Z;�&�{����d-z �FW�~]ڹ�"�s|�X����x?��f��� 託yw��ra5�^��\��G�e����t���@�P�iH�_��I�M;�X᪳&'�ɦ (��h"��9K� �~��O����~�� �W��kÄYMN��}k깅�K��aWxB��]���!�0��ɗ�J�o0<N�R0�
R�=�:2&���;��O��ESJ:���<$�(���mi0�C{T�:�޻ǉ��K�f�cU�,��.�)�t�K�K%�u$�����[�� �V�$%���2?]"?o#{z��)==%иe��Yb<���C-�I$���㫘���v�;�X�)z�%���rS=������Q��+m{Ӄ&n+�y�-�(q���,6���o~V���r �c�ڸ��]�� 0u����dFs��D�Pz��rJ+z�M�ȗ+����,Ϟ��m.ɕ�y��W�3�B�GM��l)�����'<#u���X�g�)��.Ċ�
@c���ch���j��PH��(@I��"�]E��O���#CKZF��$�T��\E������}ۂ�w�����k�C���qD� �c�����1��-�͓#'�)C�>�+[��R֚�2N�_A�ZtY�C�y3�qC��i�͏)n�}O��?��T�Aŭsn�ʬp�v����!Jox��Ie��j�f}���|��T-���!s�0�H�E�(��'XwY���}�@���pl�*w~xglqCLL�3���ĸ�G��1��h�ic��$%ud�~�,4���KV��|>
n}$<��0E��J����gx�z���prQ�Î�(�9�]��#��4��L��!9����� b+��2�38'�d�x���(�Ǌ��i��~�82 އO:�9Ԅ!�ݍ��0Lq?�� 9�}��&��դI�V��"2�}�c�t��#�B�eJ5�x\2{$��e�*�W�CNb8@6U��y!��L7���YX�H�QXV7�V.#  ]��b�N��%�?�%I���b Ph��e�\�@�m�V4o��v��#L/�FO
N��k�� �؇��4Y�҉�(�Uq/�	�"��$�
��Xv��R�����k$v�luɯ�h�p�/��D�&��%5(�-.�ě>��@ĘZ����/���;��Ҽ�!d�w�I*y!A��P�+��#���߳W(Y[�qt�O7^c���=�N�J�tC��[���"��Ig����&='q��v�j-�R�
�ao{�X��R&�Fy`)�pF����܊\G�B��W@��P���J���J�!��z�
D�m<��ĥ]k�D�_����r��$������z����#W)����>/�ԓB����?_���^wƵ��h�X�9�EU�sµ��"$��_��������R��OL��Nsr܇�*z������_ۗ[�l nԞ�� ����i��/s�n�f5��Ar+�R�`�dڡ����Ά�폡��Ӑ�P�;`��W-�OmU>���K�������_�����x5�F<��SPUljgm�G8�b&�a��	��,���ha�¦�=WD�I�ܢ���c�SЍU��u�_�9�9���b�@�@0,��;�AP���~9�5j��N��������N$�M��.{`�yi��\�;/�� &-��@�UqYn��/l�O��`����F����T�,���*?�B�N�p#Ym��� m��aP����q���n `�,1�F"v�!�؈
{�X1�٬����r�
��>�q'E�Zo�?��Q�����v�YZf�&!$}
�Hc6)Ԙ��Z�WQ`
L}�-_i����"���
׵CՇ���ѧ�Nm�����u<��4/4W=�{�*�b0�s�(�j�v��!ݰ>x53���W=�Z���VZ1\lJ���<��z���12��yq�p+xvܲ)��P#2��-m���^�����l@CǼ��>�d�`t!L�i�Ss+���[ͯ�D��$�TƇ�v�v8w-�6vG#���^��Xt٪���r���tR��n�U$�U�P�nJ}��e\���2 󔵖P�88t���[T�1�a�c��,�
Oa�
?:(��j��Z�H^4�6�>�ű�ϝ��_e��fU�6t�/�R���� ���}��)u���G@iw?T��'�[c/���Ô����?:��Q���e�8O��B�<�y��1�$�5�aJ�:�[Ɗ 8L5D��T�n3ER1��BB����:��	b��k�ϔ5}�'�Q)�t&�r����N>iyb��O�>�c"uq�XMdƵS���P��I�<2�t�l�k/O��X:DX���S~[���5%�+����4;Z< Xs�E�/��]�^�z�������S7ML��O��#��#JS�Di�~#\��ឤ�yn�j��p�.�>�y�呼)��2�I_+�+Ƞ�f�[� ����8�D}.�{����9W6�*)��,*��Dڐ��t����D'���`�Łu�-o�1T6�ث�]�&����F���a���a�����pG���"��o��
u�U8Ԯ�g�:v�pc�A�!f q�+����tx�E�۞q�;�Zn�D����7G��K�f��cߘ@�i2A��f���谆�5���k��z�N5.�T�����U�����q�X�C�F熽�]���9[��+}��I��f%L�� Eh�˵^����.F�c-���A��6�$��R�g	����2�:��T���h@�=>h$nj�~!O��c�%�QXP�XM��c
���_2_�N+.��#@Ҩ,x����Ǉ�14�/�%.:[�����"ۜ#��Σ��*BZ䓔��)���HI7*�Q��f�e��W=C��u���x�1����`�"�s<�i���2(Q���bm�es,�gBe��\䇡��}3�]j��k+0f2
���}�ي��=���+}Tm�e��O�s���G��8UA �+�o���xU�῕TL2���j�6��r*�Y�
{3�|��ݯ��専;n�a��%B6�M����F����I�<��3�3�$�,m����_�4_������R'��O�9��r��3�N%Ūb����vKW�ďh��z��?��A�l���n"�bg&ja����r���m;$���:���OC�q��e<UY��N��ã);А�#���{�R"?U�ihMË\y�}���oȖ��+k�\;��� m��HG"��&0�x	�J�Vh��G&���rr�Xj�vq�01J�f#���I������Y�La�6g�s7:�?uإ�8vE��Wi�ٳL�$p�s���}/v�+��*{��9$s)<���ߛ�#�/�,2g�o�Tz��	ܾ�����ϝX4���y���sS��qz��,wU�^5|eˮ���: a}-I
V�V��� ��\�Z�z�(o#0�Z�{Qb��	��"�IYBԢq˓�5[��)v��5쑘���&�s��n9�%-*��N�����ϻy}��5�dwE�@����h��x��ky�H6Zu@bB2�C�(4,�6R䉃e��"Wp_R��/�[=P �f����I��@�3/I?z	Od�Җ�'_�χ���a՟�)�=��ʟ��f����7� p�P�=/�*��&݋�c�����Bd������8}�8e@/���<�3σ��y1`�^E��m:;�y�"���\�:�s�u`�����F�EBX�8�f@�{.Ry\��D#��s�M�Ɲ(��s�du�Ь�=��x�(��'�z��wxcI�z�*m s��/|ϵ�H/�7yBp_�.�qE��ȼ��d@ˉ�*!"�tn�#\�ۤ,^�yYDTx�?l������C�?�!Y�����; �@b��o�f�C�Z~�E�1O���M�ɥ���#U��x���:�Be��� ~KX~<]O;���_qm�mNZ�+Byԡ~+`��O��p�]-E��{�pڢH~Ga���}۽�[e�8]w� �h�@x�n�*<!�ǖ����lx�qaz��c��� c�&e��YCj��e<���y$��-���/�K~��Y��t�-cS���ƪ0�{M�,�b�7�4Y�}L��$�ePs����K����L�t�gNv���HD����h�@#�G¬j3~q�}�,�֯��O@�k�����������'F(��S�[�� �V�̕����7�`�f3jt�mDk��p��X·��+���yk�����3�9ؗ�:��jL'��0�������h�������������MA�?�n��n��9	A֜����3#��?Y�,����È��'��h���
��"�^��KJ��l�GL�`�)��q� ���	�@az��'�/�����^ʐ�J�ܯ�M�]���ؚ�o�2�֥w�gU�Bm�
��o�y4NJ��-PhpJU��x���J�4vW��aN?�!83�%���!���Rҷ���	A���
b�d٬��~g��$�-
E4uO땭�$�[5�3dBKv����G�l�'���P��@5%�z[}D#U����-��/��uy�YX�S�Qt�>*����<+:���+��b��m��$����P��P�U�� �.)���r4�T�����	���O;������G�~_ {B�1:_?�����t��;�6���e�=�|��;g�&O���2f>>�k��"?�6�ʺ��'�P4��	���g��0r�a��ѱ>�_�l,]���-�(`�cz�K�b;QҔ��m���2}�OV3��i��t�D�d���p���IL���L�H/��x�����<w��ڄ��i���ĝ���aJ�K�OAE[�(K�bS����Xp=�=���J�ہPZ���
) ����`�mSKC�Ax��BE�zY9����`���5��ڼ����X�B0)�צ_�Xn��=�p'7B,('�)n�0�ښTa���u�C�,�ʅ^����|@���Y;��D�җm=]��-q�3� v2Z�h�u'h_�B�
��Y�6�Y�@u������\;�g����(f�D�YCŧk��~����w
�ī�����yD��v[�V�ʅ��܆;$c&_���K��K|���P���t���!w`��K�H7�H��|j�n
�:_�T?X�3��bP��ʷ���/ҹR�
��f�*{T�}~����rû�� �w�\��r��Ք�s,о� �_��̓�')��������,ㄽI��,n�'5�77
��S#�|[�+�|0a['�&Uل�˹k�vL�� �%�(���	�h��g�OU{_  �}b�!�mjI�r�� ��L=�+@�ix�D�щ�v�h$ěy1��S�(��8��H��>YF����b&����������̩��s�D�\V�<�ʏvԵz��8\�#K�w׶�ىL-�p�J�Z�٣_������g�v�����0]�N�cFX�Qv����PN�J�
fٷ� sZ�#LT���}�(_ܲ5K�=�;�պ�ĘB��J��>�3�����K'ٚ����6�q��������T��g��f����M�.�u7���.`#���98�a=G�o�?�� ��7��_�[U����B.V���A� K����d)�Cq[3#h!	���eV��
$'j��:Wk�ͭ�Z��*0}����6DE�.n�gs�x�Q��ϋcI��#��S)Qbx�ji�780T��0SL�~�vn���O�r�p��z`X�y,�nl�¦9����â`�r���>��=�x�����(�� ��Y���W����Z�]���v̠9��fO���\&�,�թ�\�?����ۯys���M��Zk��[��޴���{�a�
»Ś�T�M���"%�(�^�d��fO^�uV��AS��i��,Z��������s�~ �c�w���f��	H��'���qhL��ꑮi���2�(�^�Ѝ�`ݖ�([�ّ�T���I*k�0��/}�m�D�tP��);�J:*8�J�"@N���� �<շɐ��Z��hk��b=���0���_B��I�8��F+-�;��O�ר<��ܓ*�91�����	�iw���{�*����)b�[�����Q)��K�(�wi���V{�W6�	�|z_�}���|V;1����1�3Ҍ&�9nT^���O��^�q�_��'-��a��f}�}Jg?��|��u�HHs�KѾ�l���鮂�ɽ�`Q�p�WU�*;�ѥd�{���2�TZ��ݺDP�/=�e�U|�虁�S��H�P|:�E��Ϻ!�`l_��񏤖�L5�� 1�9n3B8���5^3��̌r�?}�(�~vY1_|�hR���U��cɪ�Y�2<�xU��#���w.(�1�Ӱ��'�O����*m��������![���`5i�b�,ΣE%���Q�?�^���#���^�"�]7C'w?i�v���97�QbI��D2���k&�?�txNx��ɅPL� cx7�9$9���4B��jb��r㒦��"jT��=�y�����<���F������_rfu�=��o�w�s�w�r{1F��O/ԯ^U�5_P2wk�q(ځ�v:��vT��l�^yD;N��M#r{" �X�	����r<��-�j��<�bŉ<�I���l8�d�N��]��񉡺�Ț�8��Ԇy�~��/�A�V+�����J������l�P�yӌV��#���"9im9���]�z�=�?>��d㽓GA����3�_bA�	��p�3o̋p�2���Ux�*g2�z&��U�x�~��>��m#�LP�NgxN�@���_1�v���B6�/n��	�c��K$7���k�Nf�T'�]u;�n����Ab����ԇ����\��Srƛ�����[�}��2Ц���QA�e��\��R�r�,��za�cpH��JUY���T����m}Q&�/���'�l�U����Cl{��K�b2�9\ w�}�V�43cd∊���]y�g��e��v����A��e����s��g���tv���_��J��
����EJu�\%�� �G z��Y�T�xQ��������5�+g;��
r�>����9~�}Hxg��@h��'	���bSn	`�y.���=�Iׇ����GQЧ�⋑+���v��������p,��j�����Ozԁ������-�+��o�wh/t�az�qd2cu�[���b�%[��
����X��G�� �E!2 Q+��n�0�êV')�ɞQ�`�㭈�x�n��4�C�Y����,Tc��i#:ݑ�`���`R�#4�U�s�x�?eH|�o�1��R&�y�1Ţs3�7�[G!q��#���w�#�<���5�����Q���y�J�Jd���{��{�D(��4@0�S���
;��7B����w��㎙��� wG���2$M0~މ���߼H�r��O�&g��(0��c}Da���8	n��4l���_�E�٘�����ǯ4~���O�V�f#KŹ����&J7�]f;���y��ܸq��jI��{*��4�#��� ����2�{Uk�U\��Yϴ�.�!@8��Y�`|F���خ�a�ʶ�
dSPaQt��Nz��mxn-��:�,0E��PG�����la@���F/����w��n������'�|�h}���V-��SV�|��S�ɚ+,�V�Q�X"��G#�F�j�F<�m��ߞ��*	I��ۯ�oĹ孖�=/{2�"�\4��@^�*��)Z	(��Y�Єi��j`�X�"�4�S8���䑍���uܲ��sv�-붅���,2�2�p�.�/�)�	1c��ZO$�|���R���'{�-�UmiP�e����^��4k��H�A4�QQ.�XM��8x�����X�f[M@�k��=/�R�����l!c*:�"wѬ,�v�I�jӲk�R�h_%AQSNlG��g���N�s��] ߙ���H4 Ҵ��\���q���'��}��y����:���8�LdÙ�c���^u2���t�ɧ����(%���d\5j��5
Zz9��6h��|�j�������_�^���̠5�WwE�����+��R(�B����9���ݩL$��⠊�^�[z]�'�$��jZ�N�6���'�K>a`Y��KN��KT��@��Ҕ��F����w��.}�j'��W��VԱd���З�ݱ�Ji��dF	�px��M"z`�r�>��)|���K�ܗ'��hb`+�g�r��I�J�T#�������6�Q�a��@o*���J�A�l�[��o��el�%� ���L��a{�����C��4�L��-~ui9Y�<������T�'�����3H�p�
����c�"�+wL!Q\��E��6ԜQ'�����e��W�P�ǔhC��gK�O_<\-�A����⺿�j�&_�;��PHz,�X/��WO��P�[�7ㆾ�@�*6Q[9G0�h-/�O�s(L��h�< ���!Z�¡XQs�ᒩ!o��2M����[U��{�����h��co�x�5�fpm<L&G`��2w���i���%�,	�,��I~F>_��*@V���D�Z"��������L|[�ve���	,�&RU��<ҙ'�Eo^��,FZc�VI���G[��Z�F�T����"�@�M�����i�%U���tO&`�R��9`M�2� �i���<�G�e	�Gx*IR�� �,���qg���~�^��"�ٲ�FS轵��9��@'��Ǫj�@5~�/�i��i��ʦ6`j��j������'&�^a��m����yE�Ǣ�G��7W�Oq�W2%^���\���v�T�X����D�0��N�Q�KB��'9j�F$@f淽$&%�2I�R ����Ӯ�+
�#d5=����X��I�,o��!�EԹ���Pǚ3�a� �g���"��x�I���T�n��:���C��ǰ	FZK$��R2�>ޮ\6�jq���HO�ɾQtd�$��F����y~uC�nL���<S�}������ґV�=4��eQ@���G0���q�i ��EN0��I7��{QZ����r%�܃���W
=�+�M���H��'�5�7G�l���) �B��y������+��N��ْ��1���/ޒ���I����xS
Hz9@��"R%=�-���`?�|p��Y�l���Q����+�<���[w����c_�\N;[Z�1���悅i��RY$����J&E�	.��"
4�4�8���c�������N�Ik�O���B�?�����2�ݜ
�f�ه+6J)�JH���\.= ���{��f@����@��O�$�xs'�&�ȥ��w�+��S2�����玲l?h��.U��y5'H����>9Uz�`;�/�)���,twS|ֻj�w��S�����[�:��Xd�HN��PJC�2䐯�����
����I"�/�Z��h��F�����s,0}�b���O�ykF�A?�Q/=eY���͍��~��|����A���X�(�FW���>'���!�n�S��������	A�j`4�q @ܿf�t�o�z�Mm�x�˶��Vp
�M����B�G%Y�*���!���5��|ŷ�]����X]�w��L�ڦ��M����J�m_ލὸe�F��b�Q�ڸ�ߵ�;S�,�0���:�zPv��D���:�dNSMӶ���Ba3��e#��^�n����]6�uq�8�ӝEϭ�6y˜Fx��P� �C����lJ7{�ɫ����0a}�s�g�Gij�tt�n��d.f�fn�� ��ȕq7e30���86��d�,��� ]������Z�o�zB� G��C]MxI��I�\��XӬvL�h���$�N�h�A��xSu��v�h�#),]I<FF��L'��)�t@�k�n.9R%7ٓ��ғU�i콲�8<��v��\.%��X�T���"�
ӣ�;=��rQFK��X�a�-{���'�8:=�S���/�4��s{�@��4^
ȯ������1R5��(e�;��X�|p���_.��+��yw?�;�T}�̒C��i q�{�o���6�>\J��V0ʋ�1Z]�H��V}��R���&�[���3��H�9a�9������	l�Q?n�Ǒ�B��a�N)cW��ڋsU��!��J��!���"��a�/�M}/���*/�¦��!>�б����k3S1���-R�Yȩi>�-�K3������C|��x��?.O�2xn�_�"D��P���x'nn��C�@$|w!q�����TvT#���*)�	�{�_;��aB)U�̺7�]/|� �
�_f�z�?#�O{�vS��rp���5���v]�B��_��h�J�3E� h�6�OI���f�i��\ה�3�CdP=T�x5�/�Yw�՗ig�"-g��<���oV��*|18Ie�Z���'�ź/A�)��\��)�$���@W���=�SQ�.��
����غ@�Q���{"�D�������mBC�������<((Z����!�/��"�Y�D��^�=�wN/T��^�z�"�Q��2�S�ޭWt��e2#C��Z�=3��!��$���b@@���C��;��D<�E��?�A8B]$�:�yZ�N賍[���`~;-(�/�,�#2�㘼�3�׋V�4%��4R��en��=�S�i�5���a�Y�88>˨����j���C�-��iOZ;�Kⴜ�Τa�	B�~ ��ς�{�� �+�e,�Qg1&R���?lz�c�K�賆!��� 8;�g�=�:i�m�����>��p�]0R�Z	�����.\�=e����(\�Do��1?t���AY�R��*#$��~�M+��N7?������Frs�wU��63�=��X��$꼙l�gN.���6��[�t'�Õ�o]G�N{� ,�s��aa*h�m��DWP�]�P��k�ظE`�+Y-\�}oo�[X�b䢳��m���/�O�ڦR=q��cГ��[^]��O���rL�j�h�:\U�/�f&���Z��`�-�3n�����nN��c.)�p����*.�o��[�?�]3���A�����h��O��&�IZE��gH�-�/��~<�ZX�|]]������Ow�j�oE��H��<#��n(�ӖӇ;�r�'C#w�&=��d�V��R@9{[5Ē'|~D,��@�f��e�!���wc��n�I��῔�T��Ǣ�,g�-������)_��-��R\�K���R;���?z�*Q���&���#F���'���M5Қ36����s\�h,��Շ�����'4�nV]1�;��/�C�%b�"n�l�������We`c��s2#��3e�kD�Mz]�,����e~ި����m���R*�ߓD��l(�R����84�$��M�Vh����zi�kI�Mn�7�����1ӤnUs�̎�n�#	�}�/c[�������WQ��.�d)$��4DC��KZ�~&s�z:.�\�X�kŶ?>�^����Q
��_a���!���m:�$�V��r�D��{	�>9���s�vl��o��oS��R��w�8B�f���.%����+��R�;�n�j2�}?���M�7��#�j;Ў�U�纓u-j{�5UEt�T�>�U�M"���N�0Z��ȷ�a:8�r�魛��!��W3r���|w��VQSdH�D�ܣ����y'}��.AG�w��<�R&�}��'~��X��=�R��� %�U���S�=4���}���`�3ٌ�kA���n��$gD7=C�p�K�O��4��a#~W�(�����M)�E�q��(�
��ށ�Ewt\����=�I�O��۟��/ϭM֡�Ĭ�-�d������U��/�o��W���*I��� ������[�G���n1$E��������O����Q/;S�
�D�傸!#���>o�㩡�D<y��sz�\� Z���&�o�ؽ?k=�x��g��]��=;�6��Գέ��5��wa�[a[��G Ī��"�CO�k��:�N�C����q/y>G�?����s=�����Z�z��gكyO�O,�����N$.{߇��|�Ԕ�D׌���9��O���B8����SU�<L���Iw���	{��4h�r^#��%�wE_Z��8��FW�Ś�����U�%7� ��2���Q����@N�Y�ߚ�Z�����@�����؇Og �A��W	���G�!Z��u�NPdBQ_!Иq��͏��I	�8B��aO�Ҍ\.Qڴ2B4���X�,�xF%1k�� >��F�㎼Wp� �{p_���m�bP�?��>m
��{\�"`�w)��z�!���Dt����^<eK	}f�vr�%���fa*�<x����.Q*�Xz���5�.�[N��R~�b�Ϗ	]2����������+��֛ɰ�u�|i��G9A*$Y�oT-3 ઎��y#��M���<��^�z�,t���O6�^W�ęG�����ϔ�cM�Ĭ!�b/�O��a(�	�+�j�����Ϳ�uo�U��h��FA'�aK�I�:?������1<�$Ӡ��shc���_���ڡ+ae{���|��`Q$�x�Ih��k�_0In�����w�Էb���"�?[�TQkY�΂�z��b�� m}��<at��/<��<oh��\�$�I�IS�:���p��jX!����-�]�,ѥ�W��sc��%mRC�i*�P�o��x	㽀���L��7�	���s�?�?)KjN�J��5���19����K.}J�|�S����UkUO� �LM�Z�����'F��W�zq{E)~u��"������0���tn�.ȏ2�+��]-"��ӴnV�	��&z�w�$�e�PضikA����6�'x �nD�sj�$�S�Z}�£�P���\۠ijv������Hm��{r�UJ=����.f;�����7@�߀�~�_�;.`%�S�r�]��>��J�lO6r/��4�,����.~8
 _����ܓ��ؤ'^�y���Cý�#��/��e�M��p۲9턜��K@�Gh#Y���I��ɂ�[�U,��8�4PZ��ބ�)�n�����%���!%h��o��12�f͞5�cL�&�5tܨ��R���Qq�iMO?�i"�� �����J��D/�~�J��L�i=��e�]�h���e][{܂����3n�@��>��f�+,�y�8���V����YR��L�:ۿ�� "�H�2M�[z�gKP]���G��ZH������D������j��x��u��8Q�]ڬ���G/�����+?٫��[ͥ���Ôg,�����Զ�� �K���XY�r���+�c�:	���z�}S+�	D��^��^�ACI&���]W�>�n��i�ᰀ��r[^p`%s���������6mɺ&�D�K��_�N��"���)Ut���x����S_8&5h���-/��Z������b)��ջ��N5��9�;�8n�ה�!��M�����[,/zNP��
��W�p��S�����4ޞ�A�"^]޸Tɋ�k�	��̺��
�L�;.M}�j+�.�bEPGǀD]Ԉ��I��5���Y�p�꛹�zYFo�`���F5Bd���8����9�������_�QΑ����	w<���P��+`��d~�ڶ���F�����v�vG��Z����J#�������b;���r؃v�[��*%����^<u��=�Wm��X<�}�.śI���������s��B}����[���mm�|Eȴ�Q�h�r�3�(��Ğ-�$w���0:��R��T�;�ʎ,�*"&���q5{�\?��Ix���q�T���Z��8fhVJ,�MS�J�I7`;�s�
y�rnƴ���k�،�\�W�I���,�lrw/�M�Y�Fx��7�o��YA�U!��-&�P�����R-⸵+�s�s��q�L�\zEc���d�d��b.D3`�*u��^��p�|r��]k�綀_j��获� m�o�B�P@դ:�1�·F�z��-�EG�j�� h��2��n$!�_���q	v�e5���r��~p�މ�=�#�.�j?�ǭD��	�V�,��V�`z�O5q���e�֜7\4Mlײ/���� �"/����X�l(��*fT:��r|���d&i&�RJ���t˗a9_Nb|6]��8��cc�]R�%(�~�/�����ڒ&T ���@2�fu��R��� F����M�:�g�δ�3��<4]y�����$D�#���@���:��I
[�¸l��d�o�T�T�x$E���0bqj�����x҆~o4¸y��P��\��*����&r!f,b|�2���H���7	�C"ot���Q/rc>� O�'�}3�x�Q�6�,�Y�7K9:+�c�d �@�ᡑ��+Y�-#�!nX�9��T���&�\vc��F9mo9]��\)W@B�9�;��C��:��,�A$���l�{��Sk[���	Rb�LAx#�3������&M}�}��Y}�9��o��Ǖ��!@�K���_,�a&�u�[f>��)��R���]G����s��_	˃"R�z�,��NѶ�R���k5zȅGB��W�p�@>�YT_1_#!7zF�{���C �`�oI��ߙu����&W���[H�z^�P-���=b?�@��@���ǵ��{V��M�NO�ҿ�{f>;�FY}��aLQC��X��ހ�?ʐ�w{��}wn\F��`(�[5#�?\ w/-fy��L���yjV��>�U����]8�0��]�)5��� A�$J�.�DipA�X���;�>.���K�W� ���T��Dt�8�}�8��>���b���jKO��:���C1���x�pW�=��M����N��X)�\y.�z��V��Tv�.�6��]�!0�r�Q����Kf�����b)��g�K����[�c!������PN�1�� �YN�V��c~Dٔ�ɨ�ʁ�ـ�)�� bG0+E���"��:5��Zq �0��È��O�ـ�H�l����K�a�B�s�L-KQkթ[Ȓ��T��/���T*��+���l�fK����4�m�����ғ�U������Գ�+�.�CwR��0����������	[2���! z�i�\%+��i�'�}s�ͼUPhV�
D�A��n��\a�ʷ=8=u�%��NNڦW6�2�=�~�WѹlL0�?ȴ(Uf -\*�G�Kiu	B�����}5�5�?l� �h�=]���>�N��&�>3�a��������,ȶ�R���>晳��p��	����ص�X ��*���;x�I���h!-�����M��2B���2�1J+d��of�\��y�5��rmrM���6��{������|�􅩁�)y��v�$ In穬D��gu� F�U�|ڗ����S[�&�j�g�I�	���E�q��)��ؔ7]��<�>}��j���Os�O�\��MA ��:�^
G���y���qskW�q�ѯ���d�
k�e�-S<���C����_�k`/k�s{��8e�������PjEˢa; 	K��d�&��<�.L��Yh���d�K�� ?��h#�L٨�~cD�6��1� �yIu�x����?9p��b�Ѭ!X��f�C2�!x�H^�E�6l(������L��^��H������>s��e�&+9�����`�30闕.���z��qz���,E2��
,@vEz?�>�NԚ�1V"z^�N��M69� *Ӧ=Y��=����\U��:��sp\@>~�e�ԧ���s8�n�����VM��_�Ē��&���d��_��{BT}��\ݤ�á4���74J|�%!n/	��$z3`!J	�9��y��w��e(�*�D�k�j�}��%.�H�2g�?
y�Ib9��������it'���I�ir��~�F�[j0FA��H��g��@���P$�.i������ބ�Sr��U䚫����eO��m�1h�&��je1PrH�6�c�6?���0f�!!�`���<��/�騪�!r^�h���1.��3�;yR�K����Fh��6��HF�]��z>;i�v�������+'�k�g5M��\_�W55�C������y�@9Ԁ�S���O�0'3��X#�<�I*8�W_��V��󣃇���3�R�9f�@�g��8���Td�������_��:�X�ө�b�0�"���J8��gΕ��d).u_��Q ���	���2p��H��gY*�}���<vk��%{�!aa�	{ZlT�M����'\��%��2��E��ʮ�/�����2�c���N@�{����"�O��5�~A��w'��	��D�3a�;�
G#Y��S�vZ~���*�u/N��;\�� ׃QX*�p�߄Cu�Bѧ (Zp�>�C$�f'HN����!Tx;�H�&KѴX�&@���(�Uc�sSl`����[^\i6LL�8P���O��BR��n]a�}y@󰶀�s�n�o��0��'1�	�z�t�E<�o ��L\7��?�PQ崿7� �k��,��6?!�#�Z=yWI����;t�2g$	��H���������Q����TZ���� I�%�T��oj�IRO�i�D?,k�v�&�שV�s��]�jk�x$������h��{*��:ޑ�csp�>��,ϡ�@��78S(����<�6?�P9�"��`�W6��i�-9�+�TbP�e��4g�[
�s��O �2PV?��x<��9R��51��q�N���ǚ�^�Ħna���� ��!t����@F2��}uI�0�j��w/��xq���&"����J�;ǎ(2��{I����q6����9��q��6%��j{T�ާ,�LY=��"��&���4����\iO�(�&,/;�����G�j�����N2�|��κ�'Z����OZ��8�?�����M�(��C5���<���3(��nωu:RaIa�����ʟ�2~��F�����\�b
0��m�~���L�	���n9i�Y�}g�yԣl��i��=>,}!��{�a��#ym�F��ê`k�������;�-w����N�1��Y�c8�7�Z~j��
'���,@���MƠ�M�����z��1���81���ssysB챡��HO jN	�g�xk���@��E�9�q��UY���s��g�cYG��]ﾏ5�e���e��Nd�8<K`zY=���׎�l�<:��ٔ��0�R�����8̇�-W\264~�3v���!�1n�@g4��ґ,�'�H<ƶ6��s?�O���w�/�z�y�ԑ�V�,�OV=X��e#���x.ׅ��Xq�L!��v��WQM��9�i��F5���ާ�`kg����n(-�0w�R�[���'�0ϕ��"rǿ�Zt�U�.g��]��5��ff��F ���A��l���eL�W-�<�E����,A���Rl~h��iv=�sg�p���	���/�4����B���>h@d��ãg��;#�"3ܧhg��X*��RK�.?�Yߤ��#fQeE�-\;��%p�G@�< }����"B3��<d�6����u����F�i��BDUUN\/��C�1U�>������w.�b�$��6��Gr���w�Z� h��>�C6s&�xb 6�G�8t0�ڪ(��<�p7��,�,%la�c:��j�=�E�l]�:�o�xϣL���
�~���D�A��0:�I�� Ì� ��&�:lp3��zd[�l�*n��S��I�o�jέ���i��|��-��� �V�s���6!A�&�:5y���Q���:>�(�0S�g��r7��g����Gh�'� q!��<�#a��4K��QQ��P"LF��j�zxx��I�����)�ؗ��/�
�?�C��'�]��U����_0�=�8�C�KQ�^r�A�}�jК8��6j��8T'ٴ��/�T��_�B���ʾ�R��WL
��YsO���]��j�����:�}��v ���}���`���J���k2�z0�U��3�d;a�����I��.�{���(6���W��ZB��Q���]�\^��'�=��ν���U�
�FYP�����(fJd
@��հRb��Z�Dף��16N���6�Z1�QQh��X�[3�޺��lѲ\Ċ[�uyM58�.k�Q$�#���������z:�������,l�H:�\�M� �{�\ �_�M��4�25�#ϱg�I�ރfu�;�bY�r���?�ys�������Ȼ)����j^��q=B��g�?Lf������)��M�J�}5;qϯ/Q���?h���� �מ<�d'"(�x�?��(��+[G����;�����խnf���a�9�*c��=
.��JK����TJ�����u�a�	�axh"�}�~h��� ���, ���ߥi~�������E+��ŨY�G�g{��7Kn��A�tZ�i�K�m������z�>S���,*Cen[熦����t'���|1��$uo]�kjbPG� 磡�u�h8�*�� w��r���l��DD���X q_qM�P�zi�$2�U�Q\�0Q 0�wA�F��,+����5.Bð������<�y)M;,��5w�8n$�������F�I��|"h�i0V����SDW��h�a�c�5��<����Y�H5�Ƀ��a
o�Z���c#��b �8}F'(���:f��a�����*�����#����d�̀_�SEP��_
%DxkMv�_��CG�i��{~�)��� w�	�@���: Z��i3�_>�6E�t�]�^�k��ڢ!A�BkG��Y�vo�p���hf��P��8���W��A5�B:�`]�ͼ��54KR`4$_�2^1~p�P��W�s^�>y�=)OV�|��t)~���q�A�ٛ"����?�C���ؔ�=�f�DZ��;��}ԗ�SM��U�j.�+���mI
�]|!W1��v�RY�=�nn2��X���o'|ᄂ��"g�T�5��X�pҜ��H� v��a�S�E�c��8d����3w�e3	({�8�-�</��k��uҌ�y?��]�Ь���*����z>�"��b�QΗǣ�p� #��_��Y��΂�uR����?��9)��n���V��.��-h⁞�IH��T������x��+��;x���Eѿ-��t��5u��ȥ���ň�5Z^2�ߐ��0���o&W2���� S�[Ym)�/��0�ԙ���Og�M�	+^�4$JZ�^-d�H�l��
��=�cZ��C�;�6�do����+ϒ��>ь����4\��Y&T���k~
��P|�d�������s�k��Z��e<q��x��B2qd��x.{����%ݼ��|����m6�� P2o.��:2�����w��i��>%X	M���W�ەc�R����䲜����=���Η��2��6�����F�cǂ�����r[a�Ȼ3Q�j=P$��r�̈́����IQ���O؋��.�)OF&qy���f�R$j�%zf;]����._�ii��1H�����A���k>A��p}K���
H(}���f7>������鞎�~������;�)?��!N� �'�����7/�_6Ц:�q�ì���tN��_�����sosz�]�%z7��L;R�~�����HlI}{8��2�y�;'^s�_���3�\����Dd�2n�#X?�*5QK�'��`�>zc-u+�k|������2���dzA�a��jyL�,�K}!�N �=P52��~�!�����VJ:��)�8��Uս�7��c}�(��/ xX��F��sZv�;�Ј�,h��,����;AP��<�@${O�e�K�Ʀ�2�͗3���MZ�@�7>����̕��Q����t�}��~�h5[�zh�W��� �!	-p����(��b�����{1X�5��h��r���'#���y&�������²W�S��d���e�9f���{�L-Y��)Z2X��u��V������ՕnM��1��!,�c
�P2$g�}�֡ +N��j�����M��ذ����]�����?��{M=����3�����a�8ů��� ��-I-�e�䅰�_5`��֔�ִ��Y2Am����ݛ*�Q���)m>�c?X/��4r���~��_̭�����g}Dvi�.��F�xa�_����[$��߅�)_v�\��n�rI�#<�R*$�����x��}H�0��z�-��a�KT��XF9b#�I��5�5����A�;��*dģ��K@0)2N��CV�w!�*�|�������c6H{6��,:���l�a��-���D,�9
#[W��>�V�ő�1��u��Z�H�"�ϊ��+�0�N��9Nܙ-�I������5�Li��o���wd{0�|�Akյq~�rL��Sx�R��6t��鑒sp�H�����V�uK���C��Z��4���v'N�AuV�u�����ܨ��P��­c�<�k�=�}T�J�X�>�4�7�y��X�{F�^��k�\Z ^��*��M�1�E�����o�}�u�P,Xt��"~nVboSE�F�n�n�9�����O�����v
�IeQ��ޯ\#tt<�POI��5Z�y���P��2nD��U��L�;GL��b�8P8
W�ixն<�����,��M�s[�� m��@�67����K����&(I���$��
b��Ò�1�H�0e�X�u|�Y@Cܜ�P�A��ע�fS�Rrr�E�������r�i�#���n��F\N��/!�:hͧ���} �L*�1)#�*4��d�D�h@5��$d���G�n��'u��$�!N~(|X�P{�&���������Af灃u��p��4���e�A����y���=��<U�g��E�8_Ը7�Z!I�|ԒLa��ѲA�7\���f|��	��s��.Z��߃�tk,l�s	�xo��c@�A�̈́'44v�fo^�/�,	ü��"��l*9���ͽ�#��tJ�Y��J�!�=�;t��,�#��+�t�4$Ѓ1I��./t �1K��7P�ɳ�yu��!�š(*;�����.hai�h����L���ǋ@�i;�XqEv�9y�|} ��?a
\�����p�`w� �"/�IBüԔ�0�Sp}�l����)Aq�}�J�ɤ�\����i�O����[)"tty+��<ߧ�Bt2�-Z9O��">6̺$�pioM ���iR�k"�����\|�o�L�A�<�*���k��8�3��ω< ���"��mͶg�5ts�/�?|J�b��!z6f<���=��,�h�"�y�5G3�]'����������K���u�k�pH0ȼ�l��n_f���F޳�t�ڃ̯�kH?�e_i��e�iq��z3�>8��ڼ_(/��ݳu�*G�z�v��)y:%at��~��s�=�0��;o�D���}TI�mf��U\Qn���$f���;�rC,@�⛷��δm�jo�U?ί�����ǰV��.�D�mH�~��%U���n��"s�Ā�J~TH�Q㣏���m7�Ł����qrQa!����"aW�`$�Պ�-��L]ݍdnM���-�+�J2c�vg�.?���{ �R<�##�(����'@-o4�Gq'g�v��B��bp�z��\��|��C�:�A�WZ��\��d2�N�G��q�7և��Q'>�������J�a��H٠ֱ�Va:t�^�x*�5�<��Sw͓�k�R� �U#Gku!���eKH���G3o�и����Ҽ�0Hua��O��݅M�!K��hZ�ط;-��;��a���h��R1�#&x�� 	����q�é��P�O���E�6ѧzFX Wo_q�۬��3e'�e�	<=�Ҡ��ۿ�I����?�\�&����{	fl����{�Zv�?l��kT�
p
UF�����@�(��:�j����]�)�����EV>�Vxfd�jR�Ä�Y�)g�g*�V�1�ԁ>��_��{d�蟎<��l��8����ׂ�SNA8�-�](�Z�˕M*���J�wn{~a/Xt�%WUe|�
dd=�� �k]�?��^��mAi�x����d#��qO���_��d�W�=�M�՝JQm5"�D�̑��حj�1N�Y>`ܠK���2Y��:��q-�{��t�l�V��1i��0��D�A�f��P�(VF��˘�0u6" ��6$h7���PE�	��!c$  j☫�FM�����C�S&+[=���~U�F� �;�ñe!>�(ty�
��Fc�`�tO�}��$���AX��G.G `��u~��r�u��(t�!]��C�\A^H�����*9��v�d�����AL\H�jOl *;�JW�׺��4;,����l��>���K�=����v�- �X�֞�>(�?�gZ���"	�J)��K;�;ƀV�O��6�������)KP��!�嶹���{�\<y$���=�O'X�L��	���,��m2�7�X�K��mOg�mZ�]��(5zeB��L�C}pla�_���`�0�?c���^"*����� ��Y�I���l��p�y�#_4&".L�l�
 �5���$?PtD}����<�Kd�+x]ٓp93rO$n���$�4���s��w
r�y�2����﨡Vp!ﻑػ�As��r#O��m�,5��s4B\�y�H&� yܺ����c�� 28�C�����������:ea�7�����x���B�.���Ukԍ�F�ٮ�oЈ k���aw{��� ?2�v�+=@l� ��<&a�*^<.z��Od���8�!Q���fiN��f\u6}�:X����*��K0��fȩ~l��ݐ]M3{·�W�uP�3�1�?�ۘ�f?5��SM�X����ܹ"��,��[j�#y1�G��2G;3c-c���M|�4c���:��E���FC�]��T��S��i{��vɛb�e��=\��@ts��&�y�v�?揚�.��������P��)�{��&߭���ZEm��&��
�1r�B���;`�v���>z|�Y��ןz��>w��q�XE"����;��x_!��:�Þ���8M���"K��Qi��xe����!�ys+s Xw��0�&5ɽ.�Y���IqwĆzJ!��Z��}3�~�M����J�[q�.�!}EU}�����,N�0�_�P�У�T�� ���#�>6�/5�y���Z"�n[�k���O�'ʹ)�^�x%��썍o`-��]�*��0�΃���7�)DL�t,�����˱ϑG⽰�`�ܬ]�|&�5I��"�\��<�8��9�-2B��L���X�Y�P�x�k-�Jy�e ���S� ���(p�r��l#�(>�'06���ª�]�[�=�dQ����*��q�t܂�?��P���+��Ƌ�`���{��'�WDGvT	�n�w���RqC�,,,��>TZ��KCw2������P{����?�q}]�^հ8�+f὜w�(��K�܈��ei� ƍ�\�G���}>��B�,Σ���e��|!�M��R��|]�+�z9#ng�H�\� z)�,�>
�8��|OW	]������5�&R�;�� �����m���U���8;G�� �<#`�)�Q�t7����+�.� `Z�	=�I}��`��� �p������Xk�l`�����Aű�ETuAFv8~)��
��n��$��*
Uϋ�o��X��Z@�}��p��)N����=�ꓞ�L����_������~���3Q��U��օ�����a`&���z�\�?��y�|�֙�T� �fs�qH�s�d��������/Ƥ��jm4�!ڥT��B?o��*GH�J(Aˡ�Xr�Y�ms�A=](i��t(�}pWE���/�N��J<mS�o�6�pW���,�������B��V�G۝�k�}�;A�c/b��n+p$"[��\t;0.NloN?9���wv���B���
C��q����f�>��2�a[�l$�o���7�Eշ8���+wF���M���`�f��u��x�����.�i����{n6'b�5/8T-B��8��Uz��$���[� yymt2���uBw�m~���j��=�=���9cʂ�ŜϏ<=���L�ļ���Hk|��>u��V�^�~�8�.�yn.Խ
�Y_%������ω<7�(����¿I�\mP*���u޹2Y�sѮ�STa*[H㳝Σ��6]����}��/b�}P�K٦c�'|]�Z
��RUf�ヾ	��u[b�4�����Lgߢ2����Q؉ݯ)}�÷$eV�����?�M]�������%APt��_���E*�ih���Nؗ�
��i�X��|xR3� ���	1���K�W�ǭ���lb�����;(��������Ό����6�l�� �r�5��L�9�6����\;N��t"���^����MJ�V@�[i����9i~)t�RÛ��o���D����&V��fG�_�>��N�3��O�\l��Ӗdh٘i|;X�Wo��~[�ej�A��f��d@ �mE�f�#J#��e�Cu�ҞX�~��v�`ow�Eꪂ�s4i��7>�'�\�Qn���\Ӥ ��G���m?����фs^X���}f� ����/9:Z�2�Ɛc+�����h%�Qgx�11�e�@h��ldU�>)�F��ΠgN}n+�c9�#Lt��s�U=z�1�{��	��۱�Ky�e�zBE�~O��3b3A��Ś{a�5������}I�R/�q|�!�<B����.��5[S���.���_D����=;���R��=v��w%��8�3_�������jT���5&A�&�[��pR�&��e�ݜ���tB��_t,��I�	R��ǽ8BS�D����S�i�]�ލ��塱Kک����z���\m��*�4�c����3�bS��X����@���q��JŖ��T���_rt��t$R3C���M37�T�8?���)�͗ǵ�X�EX]]�o������f/�%�S���Y4�z	���ƼW���;���}�Je� ��]������	�q:�|D-+��Ӂ/��{K��Կ	���]ry�y��]��7s��Wt��g{�~�X�-���?�s��<��]â���4e����9�9l{
�ΎQ��+��O�{�p�(����.V�EAذ([B��^�����oe9v�}$���.=�tb��6d�YVvz/��i��o*�G�"�Yǝ(��9?}�%䌊ɢ�]�MN������b�)�Ƭ��'��eRY�B�M��l;�͉H��{�6EJ}��J�.�׈Y8:����2�%+�z��&qP�G���=㹗�I8��T�#��A� ��A�@29�fg�� T݊U���$[�����^9���W���(TR�e�:�
���{����4^��������T�g?�0����Gk+�����[� ����"}���R�X-��L���n�Щ��B��Ƶ�V�2��o�؃e�i���}��H�mwW�:9�D������պ���L�]�=��aӝ����jg]�c�H|\�yd>\�n<����)��X�3��\,�U�*��vA�G��'4��65��B�y5�[n)�^��P�w���I��n��#]u����,�� �DH���)K<�{f=��ٮ��5�s����
B���4�E���R}%-��%��vA2Z$��B����|��eo�#�y1�5eRh���	��0>��uEL��B/+����F�7	D?=�˒M�k|;�(;�LW�O�?&V0�MD�@Q��Z���
w�w��;�u�E�"�/�6! r
5ߪfv��֡�`_�m �kB���a����J�A��o>��3f�TT�Y�PD�S�+є��#�02�\�S�������C&��Ed����l��"-��	�#��A]�D[����b)�!aZ/R,B��O��u���un����1ô�:ܧW�z��� ����Q��8����f����<�fR�O�ɍ������gCF��w�s�kk��"Ow�KhE�ɀ���e:��6F8o�w����r�%�*4Y���es�F��|�"�k�G��k��O��/R|�����A6�>9��@62jO�X�n�q�rw�:# ���ʞ8r�����KÃ���(��K
k#S��¸x[�� �pi$��i�z���{��y�����IKh����X�`�pqZB��T��	9�=�����g���C�zY��������G#ö�u�Jd4J48��dӂ UB��K_PG�Ku�'�\���z ʛ��I�,�1�g��=��Á��!mj�0���v-�KeG]􅇶��Q�
��麟n�JY��v���/VuM�.��.S�2c"�8�(@cfW�>�ρC��/J�J䜭�5��!��ݎ7�Ƚ�C^Q{�z���@K�ݻ>��!�hf�4!HkJ�IW3�1%�6��12	IXl�w���ʆ4���X���	q�,縑�Rh#�y��	A�w��ٚ��64�>쫛��%A%�-Gp�lO^6�e��Ȧ��H���:(�f�6}���?�
g���֕G�';�A����LMȼy�#�����m"U��}���@͂�ݿƩ�Ѩ���MTfB��xL]�7H�����9Q�Ӱ�7�*a
4U��ՠ��8��Z߫�i�u�Z����i��,$&]��}~In�@<p����ʚ�&�����,�4^�i4�P�UADAĠ"�,ͱ7�{4���Xq��}Jf��%���1�8HP<�3'ޟ�B2�F��w�^�d-o%�'��TPw��ԋt	����A���	�Y�2شU��>�v�du��MGNذ.��t#�t���������$?gܡ��1u����!ϥ�x�=$�j*�r,U*�����d�y���5�F&�B�W�ũ2��$aWs��BA�Jb��TSi���7p7��]l���� ��+A���r�nRlܗv��#)$2)0D2�)�-�F�?�]��ȼ<�ǅ�����2ƣ�$%�� ]�g�=]���Bȡ���>�ޞ�Tp?�	Zm���Z���0|^�+��Yi��@ºsR�=��j	gy��Z�8���=_��6���6����pG�SO`�ى��T_A�|^@D���2�W}fǯ2{�H',�ʴ�QE� 'ѐ
5�8s3��i���	�QM>"2��Չ��@�<�U�4jN~Z�ڃ���8�kL8�g�3�Uq���=PU���ՠO!Gbw^K��mO���i1[��#|M@}��j4`r���촵��USb�HY�gEחSjSQ3�:sG���8��-��р�8�� ����]�+�q���5-̄�0$��s)�*�Թ�f���)��ϿN��'T��b�f�˂:~b�h�nC�ѣ��Q���:�A芳8N���"���[�dH�����I�.���D�H�����yAk��`�
J�r2_���^lK���?ac�Rg��_s]*f:���!'RR?����@��W���NBQ�������/R�]�� �.D/�� �XDj��u�� ǉH��&����
^k�]'TOr���rW@�|c�*�a�Ol���es���-S���Mʋ�[[UKnBR��j���j�P����b%KH�����(�^ԏGr�K�M�?�'�`�0l5�H����4w�B��T�p����Gm�9~Ψ�X.�������74Del6zi���-/V��*��X�6y�ف���5P��$,]�>j�YsBioLM@�L���a�}9�_�f�{M��t!�"�2�rJm��>]�F��H�oO?-K:��C��ӶR�ѧHʂ����xY$���:ۂ�Mjc�	��e�}"(t�/>�$�x��%Sr�Gڥ��e�]
b�8��ud�]̮ӗ��'υW(�+���&���c���5�v�Uf0�>�a��γ�p�OpY�nl�,$�h�`�?�^FA,�$f��z�|3���W�㸳������^:��v��{�*+0��@�������W�O�ޗX�#����f�{�Pmt��o��z|�P�q����%�K\ӛO����-�hk|e�v��f��(M	�W'�^L!��H��`f	�q���d���Ȼ�-���g	7LR��.��Dxk�s����<�/T(�������\���r�wώдW*�m3���L��Z�g�X�`��@;w
LW��ym��t�
�����(��W�=`{xzZ�	H���gBAs�/����+N<�^�NO�i��N����W�Y��:�3��ٲ�uO���˃��0�� =K�N6.�ӮP�!C�,F���g����PZ�Pe_�=�S�p(�.��©T]�:���q�*"'�&�<�w��j���?���� A
�H�: G�������~�5͌N�_��"W��c��<�"��S,+� �s����&��BN �3��ߍr�Ba�C���sK6�r$�],Ќ	�u8����/���צ��D��m��'������U @
iH�s���p �����NA[D�摽��,nck=�� &.̠2@^�m&$��@̚��H�����V�eS��"�}y�t!Pb^�&Go'Ϭ�c���ʹ ��ۢQ}5��#>I�6�&d\�^��	�,϶@#��z2��utk#F̦��_�$�6L�vG�_�6rD$W:{���7l|
�&}�ցI4bI��+;�J?����kyW��\K�v#&I�w���_�$rQt���X�3���K¾�i�p����
m;��l�s'�Ξ�k��rim��*b����HJ3'w*w;%!7bd�C�*�@��"^W��%�8D���J�,�����?�vt��9u�go���k�#��Kc�7��$�G���x�.|�:F�S�VcpBB�{HK���}n�1�����v��r�����O��s��u@�31;������[�c�8R@ �+6�.-����;.��MJLJ�^6�w�P'l�9A��_�pW5^����a����}P�0O�@&�Wi|�RQT�Ã��g�:ya���P��gk�rif�����/�-q(d�E�N������9�2��{�Xo��iލ��³���t,�1��W���ͦ��j�%�	��D�8�-+��h��`U�p#a|(�a��zUXҊ�����S�#�g&ܯgƗފ�o�0��L����[���\#���峩��U\	躞���/�(�}�j'J���H�H1S�_�F!?��3��4���F�I�^�8����J2�i�7���y�׿�N
'
Ɩ|C�#��d�[Ш�9�`h��hw�Q��,�r-f��gp�����R֣è=*�P2b����xd�]}��TMj��|n{�©�)4��Y2�'t5ꀦ&��>։*	U�6��vQ_�Ղ*+���w셧�y:��9D%�!I\�8q�摇Mp+p~���Wz�@7��X�9&˞�8��INj@�nꯝ�Z\�������I;��m��U�M#��"�rKC����Y�z`������k�Y�i�*���#?�z���^+m���.���hs��3����|�������G`�(#�_Ȏ�MLN�j��ctp����-ݺW��X�Ў�|���u<��u��G��Z���)HkIv�}�|�����ա6��4�~h��
��/5����j`k�����r�.}QS#"���OQl��QA��`�H�JG���P�A[��V���X,�/.�`)W������c�4�b��Uێ�����HI���2��ɫ�V
!��Oe&&���G��>�60^~��a�P�x�%��?�1"��̎�ΙtB��71����ϵO���{^�d�l�9�_N�����B3��u؀�iTx����x�9|{���w�I;G�+h��l�i�x�+�!�z��o�n����a��NYM�Ӭ��b�M�ao�#P�Ps�LBnN�����*�&aS������i�$K�q+_V�z����B��U@Z�d�b��h[}�h��2{��-QK������G�I���`�]�=�܋����d����]���S�(�k&�L�~UA�:���v�e2���o^'��������GT&[�E����� ;{�Z1��� ��\\��{h�c�;��hqzp[ښ<��j^��+��^�B�&w=@,��x�������R�ژi�{|,sp�NSm�1HL&Bۚ:�̄Z?oo��^OD'��c�����=���0�#����� ���B��-��#�[f6��Z�ѝ��2W��[E����!��O����o¥�
͆�y*V�+/�6v�֘.6p�V�жԄ]յ"��`�>�e�}-W�r���_������v�,�~�:
�Ӓ� C��HMf�_�&�K�G芑�(2�ZnO��� /���X�!�*��tӇ���,"�49o��q�ڼ��*3N܇.X�h�:>R��g]��=��Oz�T�yZ���B�������dO^���If�í'5&��M5��I���+��� ��I���>������{�,�������f5�s{1[�.$�Rj�|�ܾ����_R�oIa}G@f�k�b�B\�#��n�����K��,�H(L������ڝ�Blt�O�ƃ"��D}�M�����/�X[5�.3��^xuB����u�9����ɬ^���MiR7[~�߁D��(b�^�p��y�`��Pk��d���+�Gm"��D����=���l1R%���\�1=Ls��n РL���WԌ1��km��x���ϢI�O`��}縆?j�> S}c#�6�&��>��&ZeoÜ��;Ml�_���{��K΢B����{�f�!�p��b�%�q���z׿W}�_�r4�L����m��}�q�Y{(H����+ΖiC���-ٍh�%�Hve��޲;Y{�S�S#�<��F/.1v2V�Ȱ$ny���� |�bo�z�x�HC�<�}�5L;����C��������?.z�ڱ-vI�i��YK7"x«pϴz]�=��|��S?�(%���[Q�H�f���iy�m���D�g/ HX�	��x.����u�Z��!�|�U�����
z�7�����,z��s}:����!�b�\��Ͻ�����BY��Zyb��Fxlj�h��xۋ
q>~4��V>�Ɋr�WԞj�.�l�:�B�F�x�A�T:�*9fR�Cö�L�@��d�F�89i�^��h�F�0g29��¥���g�߱ű�w�~���>Ã�Q��!�\�,6;���0yL��Qi>�����l~ɰ�>"k&|��/Zb��M�5��7|��-��Pw$�b��2@�WP�o�Ĩ��k`��T��Z���K,C�D�K��L� k��ĈN�p	��_�f��Ypq�!Z�߅H��?��G1�P���SlJu*���S����n7
�L��D=�b91�Vi�:�	tE�����:�������%(Y�E:�Q0��?��O�㕕�nK4��WP�Q���,�����f�+9Hp/���#-n����T�$3I/K�ul ��函[���w�AǘN*t��b&F�Hr�����6Ib��>!�߷t�|]�����eCRG��E��1x�<��K�*�#3�^/8�^O�m@�����
�ي��`�A�W�>,�>��3��)���u(f�q�������6(�=��?��Ưu�q_}E�9��e}Ů�X���B���lE9I������#v�3����rF|���l3�T}?�ѻ�wߏ�ܫ:����w� �dIOi�q����ş�q��?�Z����"OB�{0�����uڸF�F1-�R�z�n�g�1�t'm�S�����b����v�\,�	=2���v���[~��>$��+���<=ۘQ��)�3�v����L@	t?9�]P�����h "��� &�JL��@�r�%
���A�ԢY��?l��ԻuJ�������-h��f���.����~��5�5�ɉ ׍$��:��	ox���9Y���<�-�iH��Zg��5�w��D�:�|uk>�c�TM��:.��x��������W�����E6����Yy;��~���MQY�0	�=�H�;QUlfiٿ�_g~�+'h{����R�E���X�6����h�}�1_'�K:�)/��G4u��^���j%��;z~?}$�����ȳ�����-/9&&	d��Z�!��ıy�*;%��tof���</��n��s��Ni1�h�o�{;'q���I�6���6���`��}�NN���e�$���4������%S��B�
�ƹ�Ч�6M=�U;i4�vJo�.�d�5��%0jc��J5���iT�	�!mz��@�zJ:d,�0�G�$��ւn%gqDp�f��$��l+CR�Rа�B8�ġ(�Ò�-z�ZCʵ�Nx��L\�n�^�
Wԏ[g1m�zA�t0s�WC�v@��7���>�A��֪����h<��\Zܠ� �&��kC��jA�����r��Xޗ����Y_���8��*.`CC��%�ѝR�j3i^\��Uڠ"ĥ�t�Z>^PS�[�2��Y�c�6T�	����X���l��O��I��ۡ/���I�6.�`>+��5�?��_�@C��/mO��b���j���o/��o`����Nݢ�V�FN�C�>���tK_�>{����-6p��2]D�k~���\��g+	���oGȠ�u���F�l	��(�o6�Y�W��4+�����D��(q�����$�����u��K����q�$�eX�d�_������o+�	�ǧ��uu�B<�� _!s����#�����E�L|��?5��F�B����rPd��fe��*�2�~��c\�阮R�����,�\�ɿ��ͣg�ٜ̓Y�m�ڔ	e��A����qk#�i\Йh�?LƉ<���"�>�J���L_�(2+[j6X��d4�0m���'�_�_� ص���jUrɫ��6;Ɔ��6<0@k�J��<��M/l��F$'llP��^c[X]��CTi��O[ �� ���4F��.� �/���^/u����bd�_��à6����8Xt!f������W��?F��rB:X�}_�����U�6�����]��6����N��>��$Y���L�b�\����fK'<V�d���M��_9h*�7g^����7�.��<<?�$�D�MI� 