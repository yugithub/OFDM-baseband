��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n������E�u��#F�R{��:�b;xj���k�8������Ԟ��6���@�T9N_m��K�K֔��~4�YV,3��芦��v� ��?̚��}[C:f��$r_�^����M������كN�ڷ޸S�s�Fߵ�<õ�����s9��]#��o��Y���]�+f%5�n�n��Y�C~8ƍ���|���g&��sD2�r� R*-J���O?A��n#��\�[��T�lv���eA�.���~����f�ٖB�հ�U�����g1���~��@�
��I�T�m[�i�(����1�ћ�dz {\�@�m�*�GB?5�X�a�n%}낭R���a�!�h��Kސ�h���s��AގQ3Z�jH�ǾC�e�""�gg���=NZ�gmG�LDԓ<κ�yu�򼃲e��y��,ۦP�Fj/�������v�(���d�c<y���=���#MH��NbN��� U�Wԁ�����}�����yt"��%L2�����Z��ϰ����4�S���*l�0Q 1�K���MU�7���x�]udb����,���$� �0O�6��z��
�j�HnI����
�!r �XpՌz�t��9��� 	G�T)��1���6_�=�H����yy���OB�K�X�de�mWr�O����5�,b��QbH���؊UzK���W%sk�i0�{j�"�>N�EJ�~�R�&�a�Y�vO����s|�6��%iB!���E��r�D\E5.�w�"?<�~��G]W�t�y�i�� M;E3\Όv*@w0�l뷛A�e/�h����D?rP�9=��t�|v|���XM�cӬ��hE���P�R���Ճs�I�9�����o��C�K9�_'��� 
p���Ŭ���@��M�%�z*A�Y%�pq(0���j��"R�_he�!����a�5����}S�I�[�����h��w	F	9�lG��=Is�Bdz���N�[
E�3��Ȧ� q���#��ֺ�}�Q��^)�7?����Cg����h
@@)���3�君�X�-���88��0�D|qˎG�
`�_wJ�����yA��Hi`ŵ=��N}��qCKm�A'�(}e��I/�l0�0,j�5{�m��&1k04��A��[�,Lhe�M��F0��&9��&r,1]4�6�`�K���"��t���Ϭ�)���^):_S�2;�����)�ջ�G�^�q���g觀ib;�,t��M?:E�7NhBԋ�uz̂q�����
�oV�\�0s�&	qn%b4��"�<C[���C�CS'�o�����v�N����\���rn�LPk>�i�B{ͤ�-��QP���&�f����Ͱ���A���}�"���P�Г��g�H�������c��fדÏ����|�=t��샟X���������A\ݩ'C���1�%�k
e�#���J�v_�{�:F�Tq�G�P�+�0���<.��e��0�J4ʁ�Z��[�;ZN�#64rY�ɓ�8�.� lôk��h�\C&�z1��)'R`�=��U����x�����o��0��� �.�� 7�V����b�KP֮�@�zu#C��})�:�f�t��	1�w�M�+(kw�����'�9�8��Cf�	�=O�@�9Aa�,;�WZv���s��w�*	AB�����(�+v�p���H�$ml���r�p��5�}Ȥr�,��Y�$�<m�
�m`���;nߜc���vф�W!*������g�a�
��}����"%K/2�<���u'�]	��O�[�~���p�΋��Z�|�R��a���aD���Ʉa���\�=it}�b�x�.D���@��8�q�Nt����F�+IE��Wnvp%�o��ka�}��S�2Z��-��u�P8��Tl���lZ]���h�k������p5K��7��xf�����=���k��(�2�8T�?��o^N��L�"j�-�"�ޑ�XP�a��I�_''D0�h4[�&�������e�\� ��!�v$�]c�:��M�������ɤ��3åd�+8<��a�ݠ015����k1��͍�C[�E߈{~FH�f��pW��9.W�63?n�GYa�rS�U�ɜ*�=S��6�����zI��5ŀ��6���ca��Z�wkވ�z]x��=Eg�1���Cb<���,��?��Ɯi�M�2��21k+�Dl���LՓ"Rs��s�=ã��r�q4�ّ��WM�<���Y�K�uO}������r0�j�^9Ս�9c-?���Ii�Np�3
D��?�{����3���e�� c���n�t�\�ڝiv�X�.����=+>M��i�R*���[����XV�K��P��9�
��^/"��v�5�"��q{�T�����^j�����š;ڐ��a>y�Uu3�$�)y��p�x2lg�x�#f�nmo����z���0�ij�0��|�#��R�Ĳ��
�]��S��.=4�g,�j�J\ҟ��lF��D���Fq6��4�˅�CW�
��Ưَ�B�	A�UJtW�"]�z�L*��9r�k�M�QN���x�1�A��X ���e��x~s���G� 㴥���8���
�k���5�0L����Z�ߨА�6
Y�����?��0Mʆ$>G�I�k1�j���(�?�-k��z���."OK)�o2�y��V�VgO�:$�c����}b���4��C�Jo��xp�z�*F,� �W(�?]��U9�~븪Q)����T~�1�J�z�i�<�f��<�B�����aE�(\�$p��k_*�b�(�K��!�cTڡ!��������}��l�/��JFr�};j}����c��$�E������iB�;@��M�"��ٱJ�7�ɅBUo���*�7`xKy�qb���z%Z�&��Z�P;na�����a��Y�l �,� Ɂ�tU��42�������U�-�� iH�H�Rq�15I�(�1�-��\Q?a���*ķ{�9������0V�ip�	\U*®{m�/��z�F���wkS8:W�get�-T�\�(�-�J����������\vC�F�m_9q~�ꕠi���d(:��}��V����X�1�A����j@9�W �[3�`l��n0��E� A�_�蹦�|���(ၣ��v��'�k$�Ud3�{���`J~]:n2ȏ�����l�soT�XՇ*�=�,�C(F�V���G�%���/���ΌW�{#��!Q���_rn��KЪ����ȓ.\���=i�f���\��^L]�#4y��ؾ&����Yr��+?H��Q.�U�H�00�W늷��w�����4� Io��3�蹜���HY9��������1��O���h��+�rEN]���ܱ}Ƈ�s�'��K�0z��n\�M���}�'x�?�N�����x$�.\[X7�+Ԝ'��U�7�Cc <5�!b��a�s5��|�8�ɛ���s�u�C���ו6��U]D�������uD^�H����y�N�\Cu~�!����l����=��y��[��Auۭ��w���i�M�g�G�C�G}��og���b�V�t`)�����x+�Z���IUP�U�׸�@�x�C�ʡr)tm=?����rH����Ӑr/�D*��5t}����2�30i1v����5����Mu#L R7W�y�h��;�w�U�� B`�a*�7�<6	+���H����
�Tq`"')��,���=G_�6����C�b��(�����?�L�z�u����O���B��#��#�c�aFag<�I����d�4Y�p�ɾ�Jɋv(��ǆv"�X�N�K��Zl��:$�P����nS�|UK	$�/������(��9��&�'p<�c�օ�>rdj���p��-(4t�\^7�hȤX��r�e5M���8�� �8>�P�RЕ0b�A���}��b@S������a �Q� ����DIg��u�d�D`?G_��m�V��Z��ͺ>�MDʣ�z��p��~�'�֣����i���l(hV��2}���ȣ'�cn�;3[�$��s{�Cp�e��!���!4���^�ѫT��|����% ��q~%�T�|=�?�01A�\,����`p0<��