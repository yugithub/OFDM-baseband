��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J�-�4ϼA�IŠ��#�U�(�f���+�p-Hv"�-L��wUa
`��.�|1�{��4�ao萴�EC!��>)aV;t ��J�` �c��YNv�W��۶w�"�>��_؏y>Jjuev��#��%�jMՄ����}A�#%8���9F�]�p�)d.�Ӻ&�o��v8|�p}��)o��v��7�, e7R������Ot$����:2������,v�
��F��n�{�t�
lv�-�E�x#�8ዕx����2e *�D@������z�ک��uB�^q�,j	Ϩ�����:xR�iJ�,B�'b�d��K@%�=0�lĵ����|(V_��҂N�E^�9ۃ�F�r���S�a;�k>�!�#��'IzV�A��=pF���
��F1ތC��6��.3��٪���Vtw��M��b^�\:���7�]�ڌo�֒q`�q��S�Ab�l��P?{g��$2�z�ƨQ�t������'�ߺ� sir��NO~�s���ֶtPM�r��l���m��/T2��X8�<y���M<�C���]�����lǯ� m��\��"�c�WA)2�/A��%ÿ��n` �
N�IY23��fbd:���4챢���=�3�M#+���ok���h���'xHw���y�t��}O��b��8�� y"o9��1�Ғ}�ݪ}+:�-D���qE��Յ�EH�X���] �����p���-�x2&5#�����Vਠ2�����i��2����5W�ݱ"���r)��N�:��.��E`����2JO]D�<꫐O|�׶[�j������-�Y���'�학�jAz�,��k�@t����p�D�XC��Z�fNP�@xO�(�;,��GR�����c~����v��F\Ӊ,�����I��Pl�C���V�'Ń���M�t��K���W/VP����i�Z��vis/m?����V�z���l�(x�ei�8C�M���*HsJe�r�>��7�<���͓Xg��؞_ͅ;!y�*�.���� Pm�.X�pI���1����F��E��д��z��AP����vy8N�->f�꾇�z*Y���zQz�T���衊X�ݱE����'y�ӡ���hcoѿ�Γ��eG4\�G����<=�7c�����㨷�۷����Ų�����z����*m9F/۹�X�N�����4� ���ɫ�޳Q�y/����P����?����7���E4'����<߅@�_w��s��vŋ�,���M���m��C#�}��)�onn�.	{��vUmQ�	�D!��w�.� �QV�F~'S�z4g�H�ʗۼ�#5���!��vo�\���';�G$�3aG|otd�*�������j�j�B�H���V����,��"hQwa��64 :m%w�M{��R$�$���خ��w����51���b��t������w�O{�8-WN���7�(���{$�e�/�`Y��{(f5%oLk`�2	�H�U+g�Aտ�����b�h׸]r���~�'ee�R�m5~�[�'~E����V�>-�Ò����^09��T3�a)�3;f5�G�y�q[_�w,y�-D�aA�t����T+��Ƽ�b�?*��	��N��5�ŗ��}�z�:���{;��������"���W��^�%�q�}.F���9� �
S1ݖ�f�ٳ5"i��� a�D� Tbbt/䋫y��l�A,������A$�ֻ��l�FՆd7A3�����h�*jq8�YF�8���_���(q}~B+L��Qj�7�7�aI�/��>����r��ր����Wn,�ѣE��+�QB.��嶘�!�0�o
����܄'q��#��N�^��W�8)��+i��l����:�C��x�x��;��E��� p+�(�W�T��òwL
��@<��0Ֆ����b$� r�f�Oo9X����ޡ�4E��>k�Ä.�ظQOU�.|ԗ�M�u{`|3���_�$�yRʁ�Ғ���MO��>��4�`q?x&�֊ӻ�p~�Pf�_��5��R$�6Wgj�as�s����K���&%��PwuB$M�F�3bA5fEh�x�.���ɖ�������[c�Z�����j���R���0�HE�{���ʇl���I~v��m�7*��l� A?u����M&Ƅ����V�w�� ��K�F�uf]Z�;�w^�(ʥ ��xP�k�u\�[���zFi�*\�g��ԋT�/�}{v���H��꨺oa^M��y�+�v�<���eyL���D*>��.~�8xM���H�2Z��*Sd�6�2#+���t�B7D�+ۃ�U����ᓦ�[J���nڄ�&�<��\Q�)�gV��C�~����	e6<����iB���2(٭��gr��W�"���WA�*�����	�uk�����Z)�h�.�*)�6�]q�;�1�3"���Ul�7|x��[1��Fn����ԍ���V�?�з���u��tgk@�b0�!��	4sƸSQ���Z�ў�CB���]S�@L0x�T�^�7����QK�K����2,<�w$��Ν��.��X:]�A��(<w!�H��ӂ�>Ķ��ߩ�E����å�Ӌ��y��[{Ry᎜�9���������D@x#�w?i�6����[�̷$�s�l�#&���X	�qGI�R}D��[��=���yE�2�Π�j"�W�,�����x�S�鵮���`M$x��>C�E�M�y�u<� ��u9���PX��R\KU�D5��0o��#s�̈o�q���.�i�9e����b@�jT��^�����@Oߗ��|�[�g"|��v�x�慉H�I����{	�D��q��T�Ȕ/6���������{+�����_����lJ�(ML���,J��X"��J�?9���?��VTVc�DLrk(q��bf����7��[1.w�u�~
���ȼ@�|]C���EWY�~F�(��#YT�J��;��[ΐnNW7s�Գ��j)�����X�D�D�3F3?���z�<g�+�R%\��=�n�z0s9���Dx��BHT�q�#lF��µ�L���!z72���� ��dh�#%[@A�jPT�_
2�R��(aT�rq ��5�m��Q���3��~s�iH����;7��g`yW��)�=+?�z|���͉ҏ�8�מN�*��'%!����eb*@,`�NX�SgC�Z"��Ϟ�J�Q��қ�fBB�����Pu�<5�����?v�N�\�&��3�N��S��r�
N��$�j��N`�~�PYn__(�T�����]���F�,1V��4����\�o��
SG��n.��g`��"�1>(Ұ�g�"��������mG��h�0j��1����@g�fp���_Cx%\9�hI^��*ԜM
N۽�MP������Q�k�%TYz�f�L��v�p�(�U%�����JPG��η��aPF������\�/8͝�6�G����j
QW���	���9!/�A3��d7U��Mv̧���ဠ�hU�8]��A�b=��I�ܗ��u���j�U��#�I��Bli�w��;��i0,��C���5���8
����t���
�0M�%���f��-�2�sp���Pl�W2[}���Gs����	2��oh�!~\O$2}A��CΞ�B�A�`־�`��;V��sעP�O�-��p`�Q�r�Y�jl��>�D��sLו�ί(1�}�w���?	#���Nf��o���8��*s��������
�Y��T��HR�F��S w�"�!���Rphmzwr���/��Hə���ۉ�RMp��Ρ�����/���gK����x�%�wԘ��cĻ+�Z4o��/�r	�D�Y��Ug_T ������v+ŗ�X��V^]
�ޟ+���ɇ"p�:(hPq���x>>Б�Y�|����W�x4yuC'ي&����{-�4P�6[�'ث@L��J�ݳ ;Q�ͭ����#�G�@V@W��!h���Wk�5G��$��Xū>�j>(��i�~�]ߦ�|V@LO4�r:g�i�u��;��U �f����m�$�jB�fAi�Ц���k"��������[�A�o2���M���*�:���r�eh�rC���%2L���r��?Ȝ��-P"u[��ږ� xR#G��Б�1Q�e�Ż���ś:�����0R�R����[���� ����~�X]\j�EYKo�&�(x�
���K���w�~���罛�t����dǃ+^U�ʇx�]�P���'ϗ!��|T�t�9�.^�AO��q�s8��%;�~Bͨ�'�j�Y���ݻϲ��l�͸!".�ͱ��~���A���J�={��ߙ�g��t.��@���c�'��p��8,a�!d�0��T�h5��ڦ���8�L����R��}�t(-�%@�9���#ċW¢ M�m�w��V�B{mf�p���#`p)6���sJWH`V�a��ӅADՈu�M&oz��唿�٪Tp