��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ��t-�Y�n�.>�!ɸ�"K�x�EE٠���͹MM�k&�2�uchGE�{��*n�:�
��jIVcQKLC����X���a�>ST��'�<��N��j K�����y������@�f�A}o;
ש$�$uY��T�B�r�s	��i�8����P�x�/jqG�-t���Y���H�D�1(����DV)���M�m?
��f/��G���A���SJJ�����D�������"
>�y���F�����GL�e���iA@7���0ЌKo�qF 0,ҢA�_�;EF�� ���RѨ���n�i�ˣ���AXH@R��Fu�bs����"���9������Bu�U�8�"�>Am��;��������C��_��w�5P[��jYʱk ���d�e0�ɏ�`|���x�ur�V������j��:j�h��QI���9���V��K��?;�\�6�H?H�v	��O�%2����+k'O� $��(i�;��2[�(Ξ�@��8�͆jx�竐��ę+�mH����:ȗ���ۂa����%�:���'\S2<T�I�:�Qg�ӫ�S1���Ol�S|�K��	�)� F[�ې[d?=5��7�R��][��վ �*M�U@��6ST�?�I�4/�>��y������)�����.��F��O���N`���i	à�)�1�;�H���|�0$��^���",6<y^)�	;c�;S�GwQD�"��#����
�B�I����˄;wH�v;��ԑ���eD������á�L����꾴�{�O�j���O	� y�!-��n�e�+�?i���H�3�ّ��[�P�Y7�E �-@��.�@�4��i�"r�p��tB�aE�O§�>!2z�У�u� e"g�5��v�V՟T�8|@���-����&�/���U���Y��ϙ�l_L��%4R��}��7s]��@Y����&<�sAn�U%֗qZ�U�����>���DNT@8��ej̰g����ǁ;�Kez�'�-Y؀%,��3�Pj�=�p�@`�W>}����C���
��Z��|��L-�����+p��������� �;X�wH;8xyf�'�x�8���r/�M�=��j8+̱�8�:f&{^����Y_`�%(���y��Y�����09�%��)��XF؜���@����o��.�Vo-�r�s5��A�Ǣ�a���)F�K;����kX�PO$��x)���R�	��2��z����Q��Z[��{E-��L� ���Z�%y�z��f��-,����4RxԿj���J@��-�pua�
��r���x�p���`G�hY
��R�}�v#��8Ra'��Y,m���6�b��G�.���T[L���aͦ���q��1����e`�;un���A\푑����y�2�-�ӂ�sw��j/N��j��wg"�gXE��A0v���cҐK:s�T��H��e���j�.r��������ݭv4��X�34�<�l���>GO^�ҰWBj�Uo�k�����o"/�������l�9��r��{l�m��gǗ�تΖ��Eu���>�zcd>�:��^�����L��[A2��
�m�@;��pR�A6��Me�e��Up�o/�O�d�xA��l��p`J���3u�8����A@�o�V�v^��j�%L=�]�w(�[��+�۝�J-6��;
�v�a�l�����L����'���=6���L%���vLӹ���c��KN�"je�$q����_�H�jED�w��1p���}
񱪋S���"�r��4���ϺR��j6��a����k.���AG�(���1�-q�D�[5�`Ũ���s�.Yl����\���=�cO'�V!�
{‎~�ܜ��,ɍ����~�7�^�^�RXt�S�o>�٨�S�n 	);�dw��9ybZ���u��U�/tB��K~5�؝?*�����XF���O�4%3��b�JW
UN��k ,!�X$�MV�'����0撯6e�Q�X X�兞��>ى\,����:<�Vq�t����eVj4�9@�X��ޟ=ū��d�A��؈B�$�	A��
��)^��s�����W�	�[͍�|�&j���T@�PW���hز1a���'��PhU�$e%-��G�X�8�fl]޵+=�k=|��J�ֵ2�b
�NEn��4O콻w!�ӳ���C�ZA����D�<���x>�� ������v�S�Z����ueb���;Cð���T�_
������xw\sp3m��)�	k���`��i��KD��1H[����r�	p,owaw�_:�^��Dyi�rDu�+/ˠ�)�<�7���|��G���9$������r�&��@���@����9�^>��g������,�!�g^��ܠ�i
��i�) }Nr$��tB~먷�"� *!.̂��J�:J�5aړ*�EA��Fί��k2�
�r��;�㸤H8�.�����M��N♾)�>�{u�Ty0&u�٫���+��f.�!�/�A���o3�ϋ��p��Xr�0sr��r	�@5HĆοYli�A@��j����S�p��i���&�gO)�)E��a1��`l``kx�QS:��+���%�ݔ�E8I�^�j�l�姸^v�νQ�L�׎���_^(�s"�����Z΃�B맹)x��z��"y�T���M"K�~�L����Q�I�2;D�����PVsn_kx�5`޺�W�DZ�`�2wĵ�kAMcf��O��+���a�?1���*��6�n4@_w�a"�C���"k�_�z�dI����-�_��:�G6���&b��wW'�4�:���f)М5S��<a�;�M��G�������{�E���}\�v�̬�5ٛ�@��:��)w'W�dH7R�!�]<_ή7��
�����?�PMD��X͙{r�T���R��y@��C��c�/�3C:0�x�Q8���$Rd:#�Rx�_/�:0�� +��v!��<B��[�J�޼F�7�'��F~�E���#Yp`MW��[A�!@PQڜ����
���������y=;������Hn���\�V9+n�0�����u�׀Ş�JX��Ӓ��ƛ:#�0�pV�#��/� D/[��z3[��!�p6�&��zD���~���=��e��I;��*���
6Kp�ɭM���R�|��(x�'�
�lG�gU\��1s���:N��_^{�8�bo�Gb��"��:�ӄ�)	�|��2[s�Bk��+4�?���"�b�3"Hp]H�}p�;�!��Gﳫ�.{g�<o�% e�'� ��m��O�&?v�N�lFѯu,����� ��Rr��{��"׊D�G��XkJ������ O�
?��Mk�+Q��[r��#B;Hk��"S��Rڠ4�M�*gO�_���A�������K�`Uh����H������-ǟ�[ѱ�X-�Q�,�ֻ=GQ�)D�)�'B�2�C�g��fr�x�b����;v�n,{j�PD����FY����8S�?����lT�V�!���o�����X��+$�-(� ��+��(���b�l�!X���_��a�Ī!�{&|�Tw�\���a��N�*�ot�I�"��ܦ�����4�ۻſ���h��&}'i� V��F��;�s���L�s
�������r�	����ϙ1K�.gz�>�n���f�~[�,���8��Ȟ��>�$I�~�'z�
NE�7j��%�m���sos��Q8�)*��%�Y<�ȫX�oas���E`r���v�fnw�B�m4J�$��q���	� �\��_o�;��P9��P��LrQ�x.�g����[���E�y^,0X�
��+!j�:4�tu;�s��:�`XJ�)�b@������AT	��;\�����]������$E5.Dۘޕ���'�f_�UH�,!����Wu3��?3[���0��B����*��������?���}�_�;
%�h"�_�m����4�`���(�;>u�s�ʴ��bڵ'켆��ӏ}�$��W wc���x��.Қ�:����!�G�0��O�*�Hk���+:���v�ϼ���D ��`���K�[��*��p{����e�]iԠ!%o)�tM�mb�$��%�V�A��s� })�� ����~Ҍ;]��}#(�I}[��A��="fM��V����h˚�2߲�=v��"�'����a�.2~jtQ�����jJx�!��I���<��L�]ڞp�	S3���H� Vh>d��ʓ�8Ջ�睛~0���&���*A��]� �`<��e����Cy�E��g�\�����C=�N���EU�,����,eq[���+]�Y��(�\p���`v$[-H�2���O���/�B�vya��?C�v���Bx��� D��ЛۂMa�T_!\�����@_��d�02�F�I"�䶌9�,�80�t�ď����@��'Axt���ʌ4N�rU?i���������	E� E=yϪR��IC��E���Iru.�0xN�&6�����PN��xmH��C|U�+0P�_Gi��qUQ���zqU�^�h7Ջ?�xb��B��n�6��o���Ѽ@��>������o�bBv�M���A�[��{���/�2l��]/�7	O�� �S�e��آ�Թ~\[%�s6ft�v:6@�Ճ�U�B��?�a$�x��%�9JB�&'.�d������~�7�PwM�v�f�Pw�)�kiu*#\�f�Vl����%�Ьdz�,8�/ޛ՘f@VC9�T�:����Yeȑ���{�[l�����ͬ�Ջd)��g
��b;�MЂ�\��o`��� ��ҷ�mkA���p�q拃���z���,�m��o�%�M�?����T9KI��"���B�_R 	=r�z�O8�� ����rٛ+혩��3%�f���ՑU��:��N����xJ�K
���Pb�z],�# f0βߋ�G�h���Ǉ���>>8�&���?@xE�EEt�Q["=b�A�F� a�c���e������� ���&�%��s��#"��mt��]���C�)�W#��{B>�T`�O.v4P��M���)3|_M��o�}�Q	I�z�Թi�Z�C��%S҈��Z���91�"���!̤	_H�����O�S�3�5Ś�����'�$�d$�Gw��y�E˸/1��(�k~ZAVFg��m����#F3�[\��
���G��\#�l�p�,Dn�>�К{o�����Ч���v�-hTn�A���;�!L���:�
B��U����;�1�i�m����� �N
�U���>d$MU��n|yQ��t�-Q��Y�g��W�򫇓SgO׍�.��h]Fc�aT��9�-�B��3H���r��e�dmH�>y�w�N~.Gd{�iǴ��z��+7&�f�p�׈
�C�Doq� >pwV0!��?��"B7��G.���$7��,a�ae��O��egN�j�	�rE��4���l�#P
�I0�ӎ��(��o��\�i_������g��t�d���1w2���(W�G^ȵ1���3F���r��������:a&H%��V��������[�a���C���P4t ��J'-����n�H�I��ޛ�
1��ڄ@�O�X�3��~!��e�![ֳV�h}�6�]*5ڛ((q`���)�H��eAU�!���a*���dw����K� �6,�N�.�s�.u���s��+K����N2l�u6!z��%MDBٺ	�=��ҳ����;�3=�f���6�|@�E�*lb��U�R~�~	�%]g:��s�=m�Њ�GԊ%U<��@B��%nn����aų�W��(��f͙�A�Z$I�tUP�ϟ��C�<�f�'���d"s�D �EB)�s��g\�ת^�\.��2G{���S��0mL}	�o��CD\����򌀳?���6\8۠�,)(��<K1�����d�E~�*h'�����un�qN�Vl�$׊��>:����+k?,�ŷ����ڵ�XR�WδQs��LU�$; ���7�c��<!�zo9S(��Ҝ��LtUR��i�G�
��<p����6u嵣�ă�2!臀P���-3	F�ުo�'�X`�eh+��?%��m��Y�ޞ��Ss���r��s��(�k)-Up�L$��������-���A�P&N�d�[
��w�U�O ��m�@vY��-'��@yxM�����DI��%.ɟ�-]�"_��'�o$~4�rq�Dr��:��G��g�9��(�؃�EC$
�x�~"pVi�m��o5��j:*�*E
U�}��/��q��*]�楝�F��⭌�g�>��r�Β{��#�;�6@�?�Mx��s��]D����L�k�����5T{yM�).�)Y���`��X)��AK���:�c&�|�Oω��~k�։z�y㇗T4je�MK�gt��8N��:�!9߹��2���,H�R�9�0��b�_�����6W��b/<d_�nhY`�kA�A~ޔˣ��ԛ��b��пO��@�&��9��(���E7$�ġ�� �<�Sp&inl�~��l�9�l�ܤz\�Z*�E;��:\�vlK)��nT ��	���eX���WC5���M������^$��:����ӹ�7�,�b