��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ��6�'o��3��l�+Ƨ��un�<�y tk$���&�.Q g
(�K���O`���Պ����}k��6+m��G���)������B��L���؞u�]�>=��d�9r�'��9�<�T�,=�n���<�Ty�|(淗S�b��*���ލC�+ؗw�سT�'qH���m���(q���_�?��̊	�ܲ�Ī�Y��w�hd�
�����N�X���]Y��U���C��_o�v͑�l��k���?iԃ;��: H�ne��T��45X�(��.�����
G�2űE|1&�Δ��;Q��̚�o~T�?U�'y�䢬uA�������X�ޱ�ƭ6aM�˟yvzu�=�}��$ ��x�Yѷ4�? �ɭأ�P��&s'�\@�U���k1jaͮ�s2d��+������d��+���
���r�Vخ3 ����X���=��9qv?4*`ն�Ė����A�b?*�=T�D�@
�ZG�#a�ƕۋV���I2����H�2-�j�Y�bX\���)'�8��r	j+H3��^"��z(r�-�_l�<��Ag��+��C����H�Ђd����=j�1��s��I���nX��F8evj�^����)��)W@%���V�Gt�������0��o~����������='���'��hT��[�?�gi�l����:�o]ie�VY2�4X6�8�
��N�p���hȵ��)��K��׺P]��@����,�Rfe���4&~�ф��e������nM��fzH��R��Ҟ"fG�;�O����>�S�M4���u�9�P�d�2G�z�&&m�o�MG芸d���Q�i��[�	D� (�]��1P���7��T�Ʀ@�#�nM��l�u��3�r[W0�8gX#��n&��-��2���`����HA�y|%�j��UVW�8�aXP���ϔd��o��k8��\�c��.�m�(���[��)�2x-G.�r��S�w��HR���Ƅ!�]���gjm��ݍ� �h.;+��p 꺹�A"���vG�O�UBS�L5�a�"K�;X.v�>�h��2����Tl���(�JX��qh!-xcC�l�m$��N:]N`cD܍j0����eC^�����5�w*�K���:��pU��NfS�I�V�������M�Ȉ��"o���$�&� ��*��270/g߽��a�W�>0��e=K�E��B��XV��;�������m�D���0<�P���S��!�m��p��Dw��{$�-jP�?e[��t�~��8�畾Sq%!2�����Q�3�YK׶�s(/>^���w��0�ܩ�Yò�4�E�A
򌻂o.$(����1l��ZE���%́�C���J���,�@���xV��/�X��Bx�T��������5%��d�2�hMݤ]�������"j\��1�R���}��=��h,}	�G�dO���2�G�.�*A��'g��?���"��/?$�{��CS���pӒ���Tȟ������Ց���!����/<��aWK=/���E[G[L%�ϳ۝�o�F�7���}N֔���z/Zcz�(�0,�X��+\l��)���h�ˏS�|/�?�$�n�;t:�,������j_'�0EӋ(�`z�}�����M�U���:��p�I��L��X�EQ�������!����P�"R ��̘��� %�s�V�b�@�B�]�3q�!�����ɝm��t}ef�\���[EB�q�N;�[:#�v�������p�߹0�Ո3#�鸄(�M�J�l ��e!H h��+au�Ȥm�A���վ�[�@����|-g�A`R�>P��QW�l,<dZ�5���$�az%����'�fK��W��Y#n��fX���b�ڄS
�DׄD�m�!��UlU������@dX.��=�Wv�,>�o��e�!C��c��v��`8c���|�^�|&a��t��b���V�gm��61�h�dYQ��/�F���b_��>��u1�&�Y#e�����x�_t�I1"� �v��.z�'���}��!D�i�c�&����Ug5V�$1�~�T�W�|r��=ْ8�(@�UwT݈&�]�"�r��'H�KG,�;4y�]j�Yơ�N�U�4�9�Ӹ�Py@>�I�P�a�ŭ��;��(�h�uKn����#�����HR�Qd6���*;�g	�BA����S�C�Ԇ��&�����q�f�7x�M).����K�~6qͪ�4K�MD+v��v鍷��'�l$�b��3ߪ~�z(���l��(�������F#}��x�5�P=DG�C��2��ܜPmV�͒;6����m��V �R<'�Os��[6�@�LV��l�uP!�&�̼Ԑ��Mz��Ft�Ҷ"A98?%������!7�ɟ5Z����b���<���c60Q)�2����z���,��;�V�G�:�Ba��������Ǫ�`�#T�����]i{;�_� �W�M�~��"׆e�5���1���."�*t��ӂȱ5I�:|8R�L�\C\���vZ<�?���G̈A�~���=�R���B �k�W�E,�v��� D�)����kI�6A�Ǥ�y�$�~�@��u	��<P�s���!���e�F�;W�^ɡ�H-M����'���i��G��e�e�l�fCua�:��T�A!E�x!7&��_@@[j4�M�|�	�T%S8Ϩ�	=�U�+>U�d���S/WS�+��*�����w���Op��G��.��^r�y,]��23@4Xȿ�U�қv�q�]��c��>��{R��ۼ��;�	+X&��N̋���Z1KG+��#�d����.�3/l�U�@�Mj��S % �
��N�r�a.Г�'��vm90�D��5��G�v��g���A8p�q���dX-lB���$������ג
�����V\p�������IRn|%�D+���F~���`!�]p�N4Ч��x�����;R��t�հ��*�uz�qP���թ,{�ĵ�K�<GwR�ƚI�N ��<{8�Ra����h���QV��������B�k��D�#^���y���O�(��6
��[j��H�(��v��*]3��#I���#~�%3��ʸO���P�lm]��_�W�o��#��؃�K �Uڈ�z�u�bE��vo���~�y�c�����$aH�1����� �H��v�����Zb��]Uv#Ȝ�k~�¥��HR�UKs�T�#f�eA���ӛT��yf_|s������ժNCg�4͖{��ͱ�F-��y��U��ְ�s&�An���ZB��n��4F2u]��3�˟ãE��T�E� �J*�OB��DJ�o GO\#�R���P3��pڂ�������2����G���}����nM�Ѵ^����3�ᔸ�
<�=�}��k�L���#w?'D�%�����:6��Ҟ��DIl
�Y)���a�Wwhƿ�W���da!فV���͝@>T����S/2�K��,.���rV=#)�1�ۣ�o*�d7�~��nQ.�v��F�ߤ��S�#	���:x��fZ����T���o!��I^��G�� ܾ�x��r��\N��|�XR�T�s��!8���>b��#KNۇ�h��Ɩ�CN�Q��r\^�V4E��5��e��܏�+�#X���8y?�➒�@ Dgf=r9�Vt����a�T =�SB�r���гO�H'�x�����v��E�`��]�&/��󀵹I��}n�M���{��#������cJ�Z`e�8�&m��]hu.u�����]FN�����[_�O��q��~}[�l_��`���[�fD-'J�V@Z/^&2}��$u�E�T�'�C�a�(�H�G��"�ﶯ*N��q�X�� �4�p�s�z��DP:��ZL��bi�O�T��)0�A�ި������,:q�4O�o+�U�}��G�u� �_� ���4!�+)��k��Hr+U�A��mB��}V����� xW, ��?�*�����U�>��������Bv#:D<
� O#;Q�`�G5�ie���J�M[��qϩ��׻��T<k)@������P�?�4d��{�1�����R��z�D��8�\�J#'��+ԟ���=�iQ){�| ^M���A>`����?--B*y�f��i_yg�	�1�큶��F��K��ܓ���$�lXV�̷���t��﯈��nĪ0��Ow���*�XV^n��}�Y|zv��FC���P/&�o+�XX�%$��Y��L�����gS��؃T���\�8�x�"u��ɬ��s�r�s':�i]��F;,��#��A���E���� �N��q�8��FX\���*!~�M���w��)�����]ܜ���%��U($P���&��r���.21%x�Dd�-�vl�׻�+HW`���>i6�C�R�g$���0-��_�"g�R�V5p��kxh(�����md�G*���W2��Ï��-�xį�|�q2�}HОȋE!��"1D_�P��z�@�����^�O���������?�j�$v�,��D�8��k��$�����E��!���\�(�y2���BRZ$XLQ�g8��	�%��r9�.F�<��>�� o	���{57O�t�&Q�c|:�.��u��ɩ��"��Ls�� 9�Ӣ�b�ymm�yM��1�&�%��.ǅ�yy_R�0�6
\�?9O�3=٨��x(|�mCp˜?�{�=������O��!;R.�,՝�q���UOe�Kh��X����è#�*�l��j��2�����E��ŵi"+{L��Z�KfT�Pu�q�uO��B9qW1�S?F<O�L�@g�pIs[�f���x?�Q|�`Ne]K׼p�;s����H)/3�c�I5��]qJ.�����%�jN\�ľOH@ 7>��C)