��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#�����~H�����pl�Um�v:��L��Q����;�~��?U�b����1�w���`� �2����:S���Bq��6w*��v����m��<�,E�H����,�b�M��1>k�^��&�SV%�n��b77� ��������m?��8��O�07�����v����-��Z�h�-"�f����v�Lk��em.������~A+@$���V�����z�K�Ex�;Q�2���Ij0�P~�ZR[�J�>��As6�a�!9�D0��c7�w�䔋G���ITwߦ�8k��i\˧�Ǚ��3|�İ^?��g!��
&�GCW��'W=+4=i�;(Eq��;�1!�jE�O�UX:k�9�M���L�Y sƑ�~%�{�t�6�]CVz�N�G�3*­TF��^�J+ ���=k4��m�W�Լt�ݑO!�]�"��seq�ޢ��	Z�k���XI�2�=�<���[mGpC^��˶�ҩ[&��V@aw�9��(����5n�f,��}c��Q~2y�����gP�-��y��0C)�-Q �4�UEt1�fl¢3ma>�:c�/��c��#��uc�	�F�<��%㰄�#�Cu��y���u�{p�j�m� �'��3�A��&�$(ɲ.���)��_�Ϧ���ޯ���_}R �p�Fy&O��^�Hè���lуb�1�8[���CҩX*w���5��M����z�_ �5�"4�J��z`y���㇨9<�����ꜵ��j� �= U��J����*E��P�4���qX�~��L+-;�m>u3��[�R춾o�3u|��2��Cܸ���.�	F43T�gYf�>�9�U��Al�i;9J�o�����Y��^��}ڮ�7�X�T�	���X���m������\zI��5w�r����b��t���^۳�>e-M6�i0�35��:�SR*��_EVI��С)���+N��(v4v�3��<�h�Xs�O�����#��Ү��(^#�/�hv֊�pX^wM/`�s����hq�v�����QE��i5���?����MMY�W[S�"�O��r+,\��GWp��
X�EL�t���d�R
X�'���3�E�}����|��I��z��"�9��H�F�[l	�bE��3i:�[��r_���e�᳻f��{���,-�}x�!��\*'��t��4L��@Ȟ�����ou�ǽ�LN!�O�?j3��O�l���`[���}��j��S����#��=�m���3��C���L�\����U2
n��: �������p����
�!ݗ`�Ԋڞ��e��+/E(�U������/*��#��i�.���A�C6[\p�j���&:D��~�t�R�.b�B7mqp�M�D�1�kw��ZQ�	�F94DgJ��q�	F����7\�oݴ;q�\o�\����d24��F��n:��9V�v��ja�^���6��q����O����n�F|��Ldk�d�>>���6���0'~��)�v���Q��K�-��I�nw`��D|qZ}�\��+3�����ea��X��C&�&�϶H�T�W���/��B������Ѐ�kM�~���2D�}�zm��b0�z N�^n�]$*��+��[l��	t�`���ѻڝ=�0D�����l���c���� �h$���e)G��(]R˱�얙�_����8?�x�$��;�F�YA7jU�x�*�堶1z��L�j��j?9��.�ն�̓ȾZx<O��Q�B&ʲ�[^L�#��U層��a=X	ɃD�pf��X�W��>���ǚq��L�w��{��^
�oՉ�a���<�,Lz*E����Շ�c֨�TS�J��9���FO�T1�l��Z`���� 3��IJh�eYEu� �A����͆�R>&+uDc�{�$oY�0i�����B�3mm"f�3gqE1V���s_s(:�O�n��X�;tG�»$��	:y�$"�iQ��x�$qb~@W�Q��!�E�RJ���q.ø�i �b�� �:,�T<W��C�N�Z��U'��̀m�����#l�.~���y?L�a�L%<���S|�+�^����
h�Q���4Y-��^`��	Y*L��w����8�������S�J��:!F�D���r����� ��80,}�ĥ�Uy=Pp?��q�x�x�x\�2Ҷ<�GȞ
���F�T�kAKG/7za��>$� a��k���
\E����Y��@	�|�#(�0/�d�x�#8jp��*bs}���uͣ�}�~r�*q{Y�F�©�y�&�5b�:j<_W�������b?p����ۣ�
���k�O������䄓�i�7��V�TʎZF���ц�Y�d�K�$k���鰜1x�x0�}��9����~��/�K�#Ȝ���(����z=���LԻx�6�U�&%�v��p>U�G�<��ԅ�0��p�����h�����G�PRR 6�{�Y��0�2;js����b�M�����غ�fe�aa�t�� a2R(��A$�+���h��N>�Ri�C$Lţ�]�6�P6C�)_���S�iZ���	�6�)ӴîԘ�e����oϚ��[�p���ֺ��.�v3K+%�Y"�| =H�r�FU��_d�x��ڙ\Ɛ�r��;h��=�,��dWf��KA?�]��Ȇ�:�%g�Pz�����_ՙ��ACAx�zG��=�9�ԳY�㊘<�Ԝ6tv�&��-����h>f�2���;�����2�S�>Fӄ��@-�a�oA�7,�.���;X�` ?�৒JuW2�:
xVXX��Í���cL���I���hV���T[f���?/վ�$B?��ѷXXI��2x�yJ
: ��R��H q��8�c�$>e~�ܲ��%F咜�gN�Uy+��*b��n��-�oKҘUQ�	{����{.�@p؎����N� W�Sϵ ��L"�-����VEc3��H��r��+���C?.Al����H����!)g���R�vskj�"�j���>��D�?����<ȶ���R�e�j����nJ�=g
%a#S<8v�Q�=��h9j��p��[Pv��:����Who��V(�ny���{��p�=	<Q��6rq&�������C��>e�~?׬�6e7�ձz��O3(m��y�;y͓�!�X	f'l�Ԩ
�յ�Ew�C��Xur�p@a�F�վɪ�q�sYF�@��X��g�w����6����	�\Dou����mݼt7k��"f�Ff=�jK��NN?�K���4қP)$�:p~h����݌�l#�榦��\��"/ɘ�)���`ö?CT*�\�O�v�~td�ul���N�H�cJ!���+f�����M���ԣW`������Hζ���
�X��@�����"��Ѻ�X:��̑9~ΦÊ�ád�|,��8��4�^0c���bH�B����b���($��.�ȯ���=A���U)�8���O�զ��m��'ޝwZ]��ax8��.Y���d��i�E�j���H (�3o���.0R�������0Uʀ�SH�b�o׵�Sๅc}��+��������5�3~��.��r<=���s�V�0m.]�_F��t7��7��[~���u�Y@!'E�jqOP�kW��6��RUX�D��Gyf�� q�5�<�װ���A�;���`1�<�ܧ?kh~]�)И�҄�2��f'�RL��"���z�9�	�B˞��gƏld��"c<:�㍖�UdO0m!�'4F������lsu߭]h�Op=)��l�i� ���_�AG�v��4��?|�˂�p	��/�$^��UC�����b�q��N������$Ή�ua���(�����e��������\��i�F�J{����O5a�6�0ñ�F"��r�O�A��Z*/0�����z=��R�b����0��\ZJ9�
��=s`�Y�)���d��@\'6�T��!\� �8 rAu���0���\���|�u���������0pBQ���I�B��(0�:�:�%�斈��'��@l�r�RҐ��u%4����^t���,p�򴫃G$9����ad|Pbfm)�Pя��q G�3:��]�3���ĉ(	}�̌8O�{'˓|K�"�����0/��0�1[{�$���HGG�F��KV�c&4, ��B�5�q��!�z���6��U�Ņ7��&���LA�d(���(G����p��Û��.=0$+�P ��.��#	�����m�]w��]�j�~�F���0&~5	8Yf/1�����.'�[1&�֥�&�#�J)<�ERmoXt�\=-�H��6Y>�-����@���W��	�	�R�Կ��
�f���N���}%z�H{��wXX=b�g��/��B�>.w#A� &����X�Gn1�Jė�	 ��+[�AA,�D�=��©�����WV쓟/'���L�*{ٛ}�8IM�)�_N���v���Ȓ̛`�ĸ˱c{5)OD* @�v�-z,ބ���_q!ٛ�b�ԗ��eO�@:���A��&)D�0P�o���#~^ˇ\]��J���q�Ɋ5
�����"q��`l�gB7ry:l���s����Yf�u `[S�WR����o��ŕ�	)F^�{��烁�������`����vI0���WV}��/Ym���\�T�R���a_z�O���;��-Blɢ=t4o=�F���t�d��G�0�
s�H���X��!��OU����?��5yt1�^�5�;*�����H�R�l�����[���Y)��hJ�����V�dŁ��l�茝kb�}�f���i�
�MU�9�Ao)�����rQY�V|�TE�Ћ�S1g"��ܨ��<�&�#�W�_�$mxwg!9?�w�\�M��ßH���L(E[�!�x(cJvn�������'<��zI;�<�yp����ìֹ넙Un�Lq��gF��.hyF�ʂ�m2�T�=���4�v�X��Pz�K�T�⎁}o�2zFgڐn$�e��q�5�On��Y횃��0�Yi�<����i  �]}߹Aj#��;GC5����,5�Mp nZs� !�^ɧ� x(��r��<Z���8�G��2�Ӌ�IR�6�"��`~���!��!8��>g�g��k����?����]����S���C��kV�9�~A���y�R�� 3�s^�S:�ȹ�z��7T�D��JCo�;�nY�4q�7v@�^nn\hkr=�N<��,2�)�[f@��Q�g�F��DYTh@s��g���z��m����*şk���a�Ӧ�@�~��zNw��3����|��W��E��������g��t}�s�i�����U��oE�� a�"�"@"�d���VD �k�iQ�$M��ƹ`�cw�����������~��(�C�lI�i��O� Џ&�/�|X���� �����E*7�~}b!_q���
[�QV�;;dڑ�φt�>n�56bn@� �x��'�>��`��4RC��`�hn0?\�"0~� FJ ��u?qJ*��)��{)�ՑI�9Mzz}P���JCi�����Ґ���O��N���W���<+���8��eaH&Y�I�.��>��l�=,�B�|5Va��t�����RB4�����ɦ�!�Bʧ�ʹ���q�ƥl}�v���s����0��> �2�;l^��l%4��������~�<�4RU2�C�3膆��V���7�|3�5.��\�s����K ��Y�=u`�`��<��,+uU��>� W�33����ύt�����{��Hb=go�V��%c���	�B�@)��$v�-�����OG�Z�?�lHɮ�e�pI:����G����iLͶМMz���4mI��+�E�g�i�R���Z��tk��J�s�.��uߥ �}�� Ix�˳K��.���<�����Ql��R�Һ�"au֐&�k,ō��2_($y�����Bj��i����&bv�:
����3�
5��"��s���D�J��V�M��Q��R�T��=ׁ9�l�ƻ���'#��3�M9�4�� j��t*�9�n�'p�֢C�QK�8n}��D�"\�����bL���|�(*QJ<��0k�ۓՋ��/�Ⱥ����p����V!kv1Z����Cj��{[�O�V��(�H�&�Z"I|5���"��� ,�Y�,�>��{f��1�uH(l����Y`i#[n�9��%�C�ś�\`0ƚ�Z��A�Ok��A��b+�F߸.@l��u�N���٧�l�N�6���5�ߨ�N`ax���ki�6V�ӏ��$��IY�/�x.>2|l�1�<'���<�E�egf�k���6)��W�66����J;}p�b�l��8���YM��(Ԕb,�l�,�6��Z�0.�$�U�,8�ր��(�z��J��yk� ��v��[1�*�2J� 
d���5��6�u�4��6%s�ZX�����)`{D-$r��^�*�)J5��~��6�\^
�ڤ�Zn^詄�&��9��g�
�y�?+식v�l+� �Zb#IGHsK:b�S{*ҏ�#��}%�	���\�Em�c�%M���|7���l�'���Bg�M"$���wZ#���+��Mav>4@�����#���h�3�x�:�HT��bG����.��6�F�����'b�e�S��h�E{*Ɩ?�`�^�ɿDM��q�+�}�G��R9B$0Ց���t
�e��p�����:�b)��~��|T�epET��C"�gs��6��Q�/8���7��&����ăY���4V�uU4���s�)�)'�v���:o"p��[�̕j�W´�po�W,�؟��92M�<%�U����Ƹ�y���R�u��-�Ԋl]����� J���2S!x;�#Ś�
!}��1H�m�}�3� i���t%6�<�ь�6m)��j�����j���;����g��$�/�%��9`-F�b�LQa�t-��@��τ0�6q��E�t	����I��L`�:�LVd#���tY9 >>'(VA"���P:����:b&��'�+c�r ��zs���y0<��3��i�(�lt�IV i�5�bKm��,z��uD��4=gL!�n��μ
qh�3���{��ɼ��9]o�_�m��4�d�M�(��qk�����pCFb�vh��O�K�I��+��WJ�-P6�=h��O�0.U$K�/�J� ��इ�)�6�w��T��dJ3	ҹ&���V���2�[h��z�׾�j��95�V�L�vE鴺�^��0���"?D���g�uǲ�W�f7��&��'��ϖ�l�B��x{���ٞ�ѩ��I�(V�����aj3�)��x�)-=�@ӌ�P�ܬ��'Ѽقc�U@�`u�Ƣ�4�D�/ݲ�7vܴ|�:9��n��=��L+'�Q�W�wM1��!�jđ w�7�Y$�ḑV�g���H�V�*��sd�V.nɧ�J�ka|����y������r�wV�����/���{�^�ِ��*&��a�^��e��g��������Nz*�)���� r6w���Aз~�/E`��W�tÝ,lʦ�#���S�ǅ��� 4~Vp�}���R[~/��i:���b���'{�"1�_���ݳ>��E���Q�,���F�LlH�rƭ���Ĺc��T�{A��I��\.w4��'E�x��Ut�^�U�gy����3�^ᖩ�ڭ��D�����,{�'=+)a��ͱ��҆Z$J=xkK#g�)�Yt�+ҧ��>�`�a���*�����F6����N�<.'�	+���>���(�^���+�X���>L'�I�\$ް]5r��S-�{Ǡ&[�L����"4�_0L˕tY�-W�M�7
��Pްb����w�^��:�r��t�tZn��3�Zf��6/���1��d�����s�E��h�R+iB��8��ȎD@��K7�	�T$�n ٙu\����W��P:�T�]B���cӨ��G&{Z��	��<�B$���c�uR�|��s�6���v\����%�!�����0�\�G0�6��6(ߩQE1۾X���@ĹՇ�Ϩ��<�����Oܳk�l�Z���k4;c�-�1{&5[����Ro8���E?�Wz��2��y��/����9���[N�/:f�.V5
TUȾ�(e�b��*�h�����FW�Y�n�
r��?�ɯ��V'�;{�l�	v}ډ��?��fAQ3� κ��)k'=e%ƥ������;5ɰ�/���}jG��y��\Ą�\fC�J�y�g�EI|�Q|�z�n���T:A̈����i/�VB��`���X��z8�+�UR�*{U^3��n+~L�-�Gى���PP��C!��Es��Ng�qUoX�J��>*�_�A��6 o]�Z���۟>���j�Tة�I���<�tu��1��!�L�\���'�;��x6�G�9��pހ��j������qԮV�d�W�F%�7c���>;��|�m)��pq��܂���;��BU��_�f���o�硿W��F'=�$6{z�b��]ٝ
�s��Hp����Ms#`���_yPv|�����8�lmA�T�o��S�"�D)5���e��=��������Շ��7��t����k��E��������F�[5������$o'K�L1��H�ݖ��k|`[X�0�];~��أB.�洊�1��_`w)��X�c�i�@mD�n�mb���ŊON%��m��9јQ��0g���a�d�μ��t���ط�6�1doy���xX2�ưl�v�	�foI
�wr���+"�M���_�&� ~7;�Q�C����X@��@c�n⠙��Viz�_���4��=�U��Ι���Rj��E�
66�D�&ۺZPD@����S�Eqǩ�\�1X�C��pd�G@X��@�JҦ�`uDaf��c��}l�r��Oŵ�M;�`-�L!]d�ᷛ��,b\�����A�87��x�\������z��\/O:dm��嗢i?��OP��Qp�����3������qܦy~2���W�A���t�l��7 �.N��I���F0�߷���I������`|�o,�8#��y����UDL��)�B�	��Ş���%6�rJoĆF)������G����,bv� �@x���D�}Va�';+r��v@�E��7�m<�ÿ��}����;�6H{H )Т���1"$��*�ĉ;�������/ŀ���S
V���'��Fp_�~�J6�dS�&BcB0t2�_�2�߹�ڴg���U
�ae�ܱ��81B���r��(���B�=��Jt��6Ϛ��S�T3�y�er;ef���\
��o�#�p��ы�j�R���%��[i}�K��o�Y���oa��p�z�x�tJ{�x�e�f qQ�Tp�]���7~���wX^����}��s �P�q=B=���kp���6I�2
5��H�A��666�`B@+{�|X�f�b�G����}���� ���Dm5?5<R9F�U�����"2�y�O�����������U�����5�G9���V������]��7N�ki�P�=���V���IP���u��֟\��M,D{x�9�����5��9�.a;����7�?ϰ�W
b9�t�[5
�~��Z&dI =�n����9K���/��L�]�%���&��a�*���1�8x��nVS�%A�7��Ƣ��N��[��������zR��S�P㷭/�>}�(���_��ڦ�G�l�7}!����1g��{r����Kh���a�Qfs��h�|����򡃳�b�] +�>���*�Ž�z��6L�����Q�ז]tU\ߦ��3ҁ���MF��Q�Z���z��q��B_�8��.�{��U.��Bu�H�K���j|�#�In�|X ���H���@F&���X�8�.�
�ޡӿm�4�D�ٱ�&?=��j��!q�D[��n���%m+oE��_ �
�EŲ�j�3&���@|��v��ɏ��QF��_�=���-�i�1 ��1�\r��A��T��`L8<���Wq��Q�템8�E��h�SS,��X'�����@���f�wR�a
�����������A\\%o?�=Sd���z<%1���3I�V�w��g�V/��r�'�qrY���L������WUYs��!Wh(D;%L�F�P�`���2�3�pck�o�4"����k;�e�a0�i+?J��E 줺
��+�pe��5�]jV�n�K���6eʮ�˄n�ؿ!
�R�����`+W8/�3�XU�T�#��<K���;�j$_o�HWR�㎫�>�A1����hz=xl)�\�;���������ݽ���b������8����x�K�e�<D�C����d�1��p�Ef��T�=�0�(���D�y���VC�e�b��ψ��M�SYy)*6`�����-[��]��g���fw�a����ZWMM8��]��'s��y'��L �;�*݉��J9��g���8
J��rz��� c¢��x[xk����GU	E��:i���r�g�Sk����15��f;��2:Wx����T3@��V�dV'���s��=X���;�ۤ\����kD�����4-����\�����y����m�#[q��her]c��w�v�%���|AZBO$�Q��>%<�NRpA菤�ކ(����	1S�f��nn�g�v�����=��2�%�#>b��Gܨ�X.�������Lt�.�o!�v���F��,�-BH	�p{b	I����xJ��ۦ�<�0	��-�������Ȧ�%C��B�}�0�� �li�Z���nzY/�e���.1�߿0D�������?d��sT���=�C���0.�a��pRͽ��ˁ�7ȫ���(-;��r�0��b��%��\Œ$;���}�8_�̀�֯y.e�
�~��>ރ�GE����Lz��=?��:�N��t�`l��!Q�i�<�Q�%��X�I3u���q?�BrK�㽭[��S�5��O5IR���^/eq�M���9:�,zm'��'[��r��6z0���J�Ls��¯���d�:ĻW�-��k8$�
۬���������G����iv�B����ML+]�D���Ayr-K�$�*s���q-�x�L �f��ـp�|�Ã�{#�u��䐴� �'�u����eu��&�fw}�3�����J-�qk��nv��Y@u!c�S�)%��d���ߐ`T�䨔É����F)+7�N2�!�����'�S�|��؇�YLE��P�L�ͤ�@���s-ƹ ~h�|Q5�y�B���g�٥��$�#4iL��J5��/�����р����g��T�3 �j!D~	 w؇;���}M�(��r�9�CM$�����yƸ{_?���j� ��Q�lr �$Q�'v�@�DCDii-���8)�]��Ji�X�g��s����[��Co&_=�a}���R B:��Qo���D��)��4�G&����Q#[Ԥ���ͤ�L�aА�����9+n9���#I��[ۦ�� ���i�P@��7�F-��mN���L�&�F�	����:Q����������8�FA>��Z��`�A��x�]rڊVNjJTR�[��I�t����v���:����x_�<d&��Ӷ�p!��<�ٖA�=�4�R�����9+���xN�i�T �h8u�3�6�m�q����$5z���+�9y�Җ��X���ޠ���S�.��'u��Ҕ���Z�W=1�e�̝/Y���]�T�y@��8�>%�"q?�)|֊��"\|Y��%��Ǜ'��yZ��}+�h���nW��^���{�a(dS��>+�ab�p�SD��zL�Qot;�3�|&���Go�n�� %AQЛ
���