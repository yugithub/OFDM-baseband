��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#�����a�qbZ�dS��dW�����&�jӅ�Y�j=���H������]�����X��S��=��rZǳy�y9[V��9 ��B)�����8������#���ٶq�]�����"�����I��p>Fs�C��w9�A}�9�Y��.c� &���~�0y�ېSս�x��.V��<�TV{	.��/,����K�,��@���
�����Ѭ�,E�BQ��9} O⫝�D�}{����C�o;x�9n�p0u/���W�u�HqjɃ�o��X�6�7}˖A��!�ܓٿ2:��k���N�"zywB}p���2]�I< �J��,���/����c�$�)�KuNZ�Ţ4
\�8+���$'G 5&c}o�c�e�`���E���
���į�7�9�� �@�F����G`��R�eS���j�4�s\=�B0U��J���#t�b=U��W�����S�����崓�:0	-�FFHq%O/��^�g����t\���Ȕ����t�>m����C�M(�Mo?�~+8wLI��`t|#<!�����i}��+%��,J�(>�J����J�C�|_"��珡��K��>F޴t[����2���>�ZM����H~%0R3�e)H=����`;�u�\	���z��XJ����8k�2�Ђ�6�i�9��k�©ӨN@� ��](��?c�#�hJ�e�9��J�Ӑf�I�m7��V�7�I�����ʰ&�T���Zh��ι�:f�¤��fL�i~�|)��&Aw�����:�K3�)x1��
�")g���r,��$̭�����ů�"��>�����K����K���alXqE
��9��H����u�n��f�����/u"yZ�Џg7F��FT��0�#s��M����W��=Ƹ9y�
�����i`c��A�+ޭ�s��o�t
��A�
�!�8���*h7iތfc>iyf4S��A	tݥ���U1v�?�[lT0@��e]�E�8�cྕ��8��G�l'7) �n�-Ř��K�0�i�`���{r�N|�M \$�,��ŷvPL��"6�u�Z/E~�9�[�}zRM):/f]60k�TtU4��~��w�R����S��=ot�8�ێ�"��Ì"^��,)�Ɛ��@ MYr�v{D����w~_����ዉ+)� �m"�%dk�U�T��:�Q�i*X�xb���ś���x�ڷƭq���ޒ�����Wݡ��q⥤n#Cvd`ɜ#ȫ�]Fy�/�0�Q��g��'�Ũy�zW����1���S���zo�>۩T�n6OީѴ=��[Rt<��@��|sm� �H6A���Q�G�\c)?F!mНY�
������l�#����g�}i�2$wQF�Q|g�!a���8�zQuy�?t��U}}4�����6���#��+�Y	ok=����) �l6m&wm0�bp:R�O��{��g{�?�Wv��6��@}�K��2Y�7�L���a�I�f�R��~/�V%�fuk<T}?���c��W&�r/`���X�i')�i�m���Ҋ_҃��.�a�?�N⑐}q��B�9ӭ��Q�U�5����vR��c��@���� .ĝۓw�+cè��U>�hz2[X�d
�j�I2���M���Wm�������ĵ���Lk~#HɼA�i�X{�B2�fy��f�ð_��]B�:��Iw�;y�ś��j~��l.Q�2�b��&@<��_���h���!�ڝ))g�U���E�6��0%X�E�@�}��u#�����N��
2�5O�&��|�L`5��g��it�>�����2ڴyǥ3i�,�-o�}�P�X$��-��S|P��E��;����f�oT�x�u�n�H���N	�w�F�D�~B���[y�!�7ns�(hј��|��=�r�*;X3P�F�x���4�uɷI��l��xT$�A\�N�,-ծ7�r֧����nA&6/0~�A)P�H�\0����Q���5�Z|��}(�WI�BL��5x0��RgD��X�Ӹ}�0��M����/O�G\Eɒr��\*~SS@�)�z��b��;3�JV��`+���OR�{���҄.|5E�j�H߶�GI&	�BG
��1M�&<�\��H��S#E�^����޴/)����uF��� dx;W���s��\�M5� M�<�@��*H�CY�&.z1�ح��J��M��e��\?��*U�1��ˋ�4�G#�Ȕ>�#�ߦ����.�]�P㌾�������z��b�䷗KL���VdF����L7�~O蚇�I��_���s�Q�1
g/)�[M��^If \>z���z�L"4���*(e�8��C�MYD5
�j�Nj��z+L 0�bL)�~{+�2X_[O����D�/�eR������<��a�XEf��2�q�A�������Jq{����]A�����D��]����4��:���.�a5�3���dl����:K8��8�n���f=qa2k��Ez?刯�1�J⦱��B�nj�W�./&<
��`,�k����ݫ)r�ۑ~�
