��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6>�M56�M����br�x�Ш�ء�J�
���~8+�`yAFC�#?�di���>�á��e�P)���m�Q����߹B@�|4�M�ۢ�4�5sV����\;��
��O��Yj�"ƾ$z=-������E	KZL�,Kc�A3T��b	`{[)�|բ;�"#w���*���#a�ǆ��K��E�Ml�5��~d�L�زWn2�A��aYo��O�!�d��|l����ީ/��k�^�aF��7���;���<��� �O`>����+�YNN�(�aY}� ^����١��7�����F ��.�徆�WZ'~��x�:Έ��.���#?��m�T��"}2�����	��y~Q^�m\��w�F���z���m=#j�( �<T)2�w_�>�����]��I�S�%�^��Փ�Fh�eڧǆc�8C�af���{�#	έ�vv�h�Y�Ww/���f�oq����F�Ot.��,S;�P3G��V�ej͎l��1�5��ܡ�֔�
��|����c�T�V�z�h$jOy�܉3Kd����6@���쨜,A ��y	�����ؖ�m>��8q>�
���GgG��ct�kr��|அpNq^�_�� ';�z�|z.@m�	%-Ё�\	��]4�S�����c(+ǻ%WD�A�iq\��)-�-M�%@8}`Z8��`/N�`ms���j��H��hW��'��U��d���@����|����P����]9�C�j�����]�^�X/tGíK1��ȋ~�B�,J����l[���?�6}���[a-CO��=���4�̡3`a��"80S�a	P���y2��P��g���d�v��lZ��=�D�X�M$�֍ÏO��!0A��zp��yi�8Դ!��AnMX�A�%N�>���*_ 9%���Dn��$w��?s�o>��?y���C�_^7�hX���(��X���Ep�#kӻ,ס����?��RBcʅ�5�(?_�(sZ��sr����d8r�R����Z<\?6�bk�ݕβ��>J��=���ML8n/���fϸ��ùri�Ul����*�&��f=��:[ͻ���������r3sC��ۖ�����ڊ,��9��K@�M؍y�F^*���WV��V�C�1��n�]�uư�6��y�P`ȥq�QEh�+���ް{��v<�B�w��`_��2U��m��$��N0e�j"T�v�V5m�)7�T]��C�O_��InB�vɢA���a�}���IS!9|pzJ���|�W��
����p�_,�v�'��;�Uz[��uڂ ��:�%�R>�b�8�@��3dN�
>a孔(��p�j^�\r���nZ��݋��D�W�-�jm^k;�R���?��buMmҕզ�s��� ��������Ѱ)���_	y)b4�xSz�9}p���'j#��w1 ���D����(�?K��07����^�A��wD�y�g�>�Ǆ�>�U�^�7�cy�;MҘ^��r�S]���O�f�7w_�T���Փ4�����ѕ�ۿ���P��+�<�"L$B6������J���]
L�W��XB2�����|��2a����g�D�9I�e���u�Z0�G%��S�X]B��)��v����6^���oÂTp;��{�J��U~���]����狼c_�Q�@dMlee�j4׷Ι�fЖ�+�W��;��������{ñ�h�π�,���.�n.D5��\g�ӻ�(�̮n���Xw��~�ȃ47:�N�����Y+�W�>��-�J�}���B��W����U.����9�>;U��r6��;�Ǽ�C}/vܦ�\G�Z������!�HQ�v��3bF}:4u��4?>�S%�G}2;��|$u���l����B����D���c��K� T�l o�wt�7�@rG1 ��c�\�.+�@���ùa��Y7'A�{C�w����?�]5�Gzx�����?�sE�h���;y����{��y���#*�s?"��kjfw�}�gk#�[�bY��ql���2��ŻX�mg����>O���f��*w��+ו칊:J�6X��L�ٯw43���JZz2��.���@c��(ICj	�-NK>��\P3�Fq�$�(�j�p�?�����T����<�Wua�s���ex�����ǁ�Åy��
���5'����}�����Bcj�@���Q5eXerG6�e�?���öQ�7��6�FG��W˨Â�=>��K�0�a޸&����O���$�Hl��Þ���v��,���G,����H7��?[�ۅnX+�8�mBR�Q~�d@*��6ߝ?�K�T"sα
[���|X|��E�����b�a���C�KZ���9>m	y�R�zD1;�߲��2�6�er����0��vt���f���.�r��\{�9y@�~�@�ұFh,�&�����rboOq{$x^��-{��R�"@��D�]/nBLw�-����3���� ����鹛M7g�y`)g#�a���$��}RH�|�� �w�LnG����������0r(C���蝄H�zi|E�7Θ ��ϑ�Tf�c`��qu����0zH[F*������BD�:��[e�:YsՅmspX/�U��ܺ.���eLh�H�����/�4:��b�~w�$���6[�0�^�,�݇=5g�Q�8Q�|'�rq=Y�2ˍ��:�Y��B�a���^/6Қr�Ν�%��ǆ�׾�^n����h�.}������1��l\3dM+eU8�KG�uQ
���^9�3hύ+d����h�ckL�ü�7�l��:��'/l��y�Kh����}�7�a��ɓa�Tt�����ݴ[����d�V:���Pg�k��5��A!	WN��18VcM�E_h3Y��1�jI��,��DJ
�
R9�`�.o�Vz�g[����L-{�q�Ȯ�����[NL4����rF���tUˏ�.j��s�f+D��b^3T[�ȯx"��	D��#� 4&�:�M��4Q������{�]P��q�Ǭ;�I-m����`��h�Og_
�l��F�e��yԩ�Ԗ�<�,f ���.U�^��O����p73&/��5͇��⅕���ZW�6�n��	���5�RJ�J�X��G��p���{��P�JD��f�<�Q��&���z�b�*E�Fc��	U
����P�V��1W5��~/C�E~��0ĩW8�'{�<��^,���)�b�{DV(?��H��L@=�Қd�k��JQ�R��f�c��X�paX�}F�Ԥrq�&��|HwRL��{�Wė�����"=�v�k�q�D��l�ax=�8Ĭ�cIc��9w�p4�Α,VzV����N����٭
C'x�s�I��ed�b���wʋ�G۳3b�vl#�&d���Dq_��{t�T"8��Li���D4t1R�*�ٯ�ռQx1kj��!$1o�j7��"����j�h���kWyT��8�=�\,v�c�N�4B����IS���$��F&��z��>w�Bd�2�wH�}�����H�A���>x���� #�ɺ�U���X���k�d{��͎�;}�t$tZ�8���v��8.�< z!q���>^*�­���ȫ�D"�{�ļ�"�̿��|\?C�:��1��������_���­���E�$�"��

.���32��^V��D��B�Do���6�s'�Z��9kx��D�	����1/�"�aHq23��gB���,���L����L=\ƾ
����?X�9�`7��B��E%���M�]����Eyh�5*e����w����{󔇷�m��f��2i����5gf2�#]��=zq� �V�Y���k}���2��Y�|���q,���V��?G�����%x8l %��"N�����\(�vEt`�'�ob�����""��+;�+�N��\~"�K����PR6���hwQ�:�p`��z�:��0��RU�5��ȕ�E�}NC׌��vT�Z^��R���8Ƣ	�f��B�� �=\��=ʱmw{J��"�1 ��i$��Ʊ��-��<�6k�j�!^�jI%
���a��b1��8��UT�@�d�j���U��"��g:@��Aɇƒ�6�����[���0D�\?�B�d�~"e�\�٣�b*��ʮU���,��� �Nq7 &2�$
~Č%aV��z�'x�"h��9U'�/�!tٚ0g�=�Ud�n)=i��]�i�T)Z�Z��H���E���=7���=�Cp\�'�!��2��^����c�~�hM�~v/Ă��� �S�{J7���N ��E�eM�2��:e�I��� u���*lw�+P����Z+UJB$���4U��R���mZ7��=zn\.��{&�A��4C2B�9�T9xx��)U����c`E|U�x�y��}F�ϗ�'xP���:�cΐ���ٜ͵���*{���u�P_/޻h��T�+�v�Iz���WX��&^Ϲ@����7�����ȟn�����q='!�(2I-�`�D���]k|�z};�<��N.8L���F�	q;��c�:m�y��E�/f8J5�����2��są�dG_`+���)A���9��%N>�S��z��)��Q��tB�*8Y��g"���`�X�
)��N����KJ��S���&/L,\ｳ8�'�"$��m2zM���l�>�FdK7x�UN�f�u
~[s 9�&*[5f3���C�q�+'��7!'e�u��o�W��48=)I�3(��<j8<����,e�^S�rw7s�M�p�]�:�`�G~dY���m E�������
<_/M
��3b�-�5v��>�݃1�?�D���$�ZN�w�"�%V`o0;��D]z��.�E��AB>�GC�%���s�ƍ���7��j� ���R
��_F1R1�8v��ނ�����������H�����́c��&u�p3��	�oC���A���RL�T2��	��*K��ڬ0���O��.���p^�h#�� !���!jg�!`.Ж͢��Ԍji[�#t \����=u�w�D���3�n(0l@��v�0�����g����H8!t	!#�vx�y���$�'�VB�&6.��6喂�ǉM��>$��f�:=l-���-��L�!���Oh�|�^;2&e�I("W��>C�JA�hW9y�+*�*�J��V�'�)ϊ\�
�E�/��$5�#�՘����f�� Vl�W�:S�~��q�Jt����M���i\a���n����׆u�P�"L��I���wzY�7Z��8'k�I�+�_�϶���X=�S,K4����@$zE���Х0ه^Dj����6d�'b��ɽ�����R����`��m�r�]Jу�.�@D���]x�˴?�:WN�-#��MԵv	��I����>��bʑX��m�ْL��Np�R���7�$����i����Kܙ�B�Io���_��S�7�Tё"��r�'��8*�8MK7�k���s&���{�yI���*�ܨ�_x�� _&��R���B��	''�h����Q����\�[f-t�z뉠��,^qN/⏅���u����	��w�
彈X0��HGBVn���G)�i��`K7������3$�6��ɦ���۬�9)��FwE!��Zͪl<{W�B���6m9�RP��_S��zE2�����3�V#�F��R0��d\JJGdRB�9�ӝ7�2��;���nlA/L�,�>Bd���#�M�qJږ+��+|ڙ��{�͙�L�Z�i�/��D���{�H��{���]wZ'�mO���:�gܙ8>�I$Y-�33�b�}�"��EM�� >h�L�*�a��r�))�X��"�:�_���b�J2B\�����r�\��#ַx#]�R���y�\-��=+$2s� ���I���Dw-�r�bu��8���Us�哓�P�/(j�&�Sb���BSb�%�p��� N����߈#@�W.3�3���KؾYv����j! |��0����g�&@\�W��_rҗ�hV�b�H�������&R��ux��2��lj���P��2���cx"d�O�l�1kL��'e�������8���[�D�d7 e(x��4g3�ΠxB�E]#f�s�=�
��m9���nz�ߌ4{��wD�^���!;J��f�`���Z�NA�����	��F,ZYԀdI��t�à����~S��!>����P�mN�f�܎�]�M@Ƣ��ܽ �_�&�ó��h~����{t`��@7NK 1��Q)ebI:A����l��#��2wh�*+Љn�7뻜ŘG��fF]}?�84秾YJ�����X�2����"�a�.��Sؓ���ؑ�tԣ��5S}ݺ���������*��F��dtzO����S��=N�_�+Q:�����{H8��Wepp�S.V� �]+�֋3�0�cʺ"8&~x�oMN6�O$�q����N��;�_&��<�.�Gu���,�q���=�����Pkˮ$z�Ƶ�,x��U�|�؅�����/`�/Y����jSa�L*��QyLBU�}�RK3Ե���4�`�qþ9�IwV���VK���u��b½CjїФ
�}�ALՌ����ހ$D�̓Xϯr$��w�=^�)��X��a.]K`�z�3���H$�z��ԲH�}�|����^(U������l8:���!64��L�y1��|y�e���J$�`�G�������6��bT��H�U�a69�麿W�ƨ�I�i�^�aJ�� ��\��!߳=��j�Q�u}S�h����-���ѣ`�u�����<kR;K|���E�%���'�̈́nӣ����0<����T�k��8�ȸ��Ȃ�:$I�̇�,�hA�ekf��5�4t9-��ϊ��L�Z�i3��;���`�/�Zv����0a�c��D����j�W��6�*=�!R�ob�m_�(ἅ�X��������W26	���=gO��o�s��T�noy�-�h��م�T��UH�{0T�/V����)�0�W��'�Ӷ��@w��g�n/;�K$z�A��CyE��-� ��}(>Ō�U 1��#��A��$C�������3w&p��"�Y3�0��Yl���
��|�n]��.�G<�?������Xe(q�����`޽��:��ݻ�/^c�{!�