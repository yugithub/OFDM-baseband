��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�X,��W��l!��g��Wxe�Q�,Õ�LF�rP����(pO��L(9q��W��:�n�Zj��"�bޥݤ��L�k�c�)+�Z^���k��v����$�+eP	������	����å^�8���GYu|f�]��o�0�/X֡�'����-��9�V�Uf��"�n�A~2��~+���΋������TZ�
]�t&�nQ����r�D��N(~.�#�v�&� Z*jt2܋�̵�D��|@4�1Z�XG�[���I�6W��S;idE��8"3\e���v�T"%C6:����R�8P�1��$�e�]���٭c��S&?%�n����ɨ��,�䬁� ~��@�SI q%��[��e�';d���i���W��YhqC��U��'�C�.���������D��?a˗z?4�����;�,��R����C�mftv�9�,��3�����%�Yȩ���6n�(a,ǯ�wJ�_S����i������7_�!`fy&�^������Mw ɔ�$�������pGy���G���N��[<�t��>�1&�f�z�q/����󴣡$��hRɽ$���4[����2�Azv+�	y������H{y��C�*�e'�+J�!��h.��^o �xA�EhDH���cN��������09�h�V��/� ���r��p�f��!30j	�8��Z>�Td��t����~o-�!U }�.!P�jٳ[�A��A�� �h~��j��-=FЭs���$�L�.˭����WE-q�w�\>�2�|6���J��x���p\Z�۶�X�.^�4{�ٺk����I#��(�K�i�������do��`H��{OLԤfF&g�H��[��BQ��j:���~�T)=L���ߡ]���y��-��׌Q\	�{(d�c�.�����&�Q�\��?L2��7�����	���o�Fb(F/|�m�6�}Pe���O���y�Ǭ�pRA�u �
^m�x�Ue�u+֝&�y:��{(����D8!L�#��I�6ÚJ��k��^͠7�������N*`3��d��b&;]��$\'�gl��$M�JS�k[����9m�g��;}�����	����i���s��.�S�Z:��M�0q�ۄ��	�ZQ%�*�	����X����:)a�7��t���yT'�����nq ������(��
59x��C�Ͻ;������tOPvK6w����5\:YN�D��n�����`^`�G2���1.�D*�Η�e��ə�������X�ZaR�Xe�̼����o&�X"�:D*6�^,M`.��Q�=�Y��چD��fή�*|& �'�����ܰ>�8�ӂ���s���<��({�B%�<���������X��@�����Ij����5iaҷ�+QN�6R��%�Fq�?��,�[+���.�lI�-���@�Tc�U��1+_x2= ������Y�\#�Gh�+?r���s	�U�Z>��4�?�����L����z�]�G2��xLZ	�>���w�F�"�'�˔
���#������R��v90�}���6?��(�O.R'�4����d�ELVJ�{E_����t��OM��<|���;8l�E|��ā�Q�P� %�]ҹW���04����� +��j�h&:�]"�\��kv�
��D>����`�"��b��(��s�VzD�4��eB,�TM^w�u�2k
�7+����jL�D��r�/��L��n�KW?�Z�C�޳1��i�9ޏ.X�3ͺN����#�V�;�J��_��.��W}�_Ĳ�N
���m�fG��`@��T�!�I��5���a}$�g�K7HS>���6��H�}�������.4�\���̒[[����^���z�Jku�M�d��콇�ƭ����5B��E�z�e�ˋ�IX��C?�$��2�α��t���&�?3��A�of�c+� )���j�_2P6~�Ϧ"���AP1��Z��R�fVqyv���4��ؐ�>,sHRc��W}��!��|���(�.�b�϶�r�K��z����� s�K����i����"�p�0�37�E�VWMעi=	.�@���l���G�̗�)�b�����Wq�C�MQ���|��nϳo��. }���k�+�pK�e`�t�:�UZ*iEL�:�>��0G
-s����}h��vGW���K����Ћ���S��T��Z�J/�J򬇯�]�s�vS򑢴}A�-BP_c��T�Tk����C�V�2�'�j_��!�z�C}[� �1<�?447xZoڌ���GZ� ��	*O��QK�'5�d��Ϝ~����Ƕr8��f����2���d�$qAqi(���`��q�AQ*�usvf�]��D:ú���F6�w�hz�:���t`~F��*�۞_&�M[��n����?�t��~�޽N:��]>f��w��V���d,��۸�N���$>�¸f�@��0��é��&�		�'����\X��cz���������	�b<�÷B'=�_�V���pǅ�ȵ��3���|�Ĝ�e���uÈ'�+[�u��pH�.��L{P_�}	����u�E�7��.���^N�>��#��¾��$��������^ tBD������h�E�~Ҹ�$�+�޷v#_j�B{��g���A{ԇ�Qq��3�I7�S',����wDퟢk�<t�ܻ��S��f���g����ٮG� ���U��/��x����7+�I�=�aMƟPr�!��pP�%�7�!�~m��M��SǙ#5$�;|� @m���������/��7�d��,�m���C~�f홁4�އ����f��%��eL�I�����ۇ:)��Q���ˎli���R��ZI�_O�N���R��vc��K���(���R��������#�`�5�����I6V����c�H��e0%�)��*{���f!0��ҏb���VW�J9@�+�hS�M�&���,r��5M��+*�!E��vc�T3&h�Ǳ�N")za���KؚC~f�v��@:o��%����<b�����Z�!�Ȳ�����O����T�4م�3��2�a�6zDm���f	�6���]���^%��(���;<�(|���^������	XZS�K��lCRSp`hw�LL����4\�&m�/A4{��/���&�W%a�)�`��]i*�T�q$��O�+s��g���l���U��ټKo�,'K۱�!���a
I����vL��?=ى�#�F��ufN����{~���r	�o驖.!�,#%�� �JA���4��5�۳w�?r'��-�6%K�� �6O��J��rWU��
�_|PbL�����F�b~T:�Sm���F\F]�c!ݧ�b�c�J�^}U�.��2_ձ��s���3? s�KX�lN"�iv;/Ϸ[{�4��t�_��'��ȏ~�:Mo�(��Z��f9� ������f���ʈ��[�� ���X�����ן�O�$�i��Gl]qv.�|=�\ =�E̪P��ʜʌʋ����bE۫��XM(�}fng7
M� /p�х�
�]����!�v"�����;A��A��1�a���[��i�۠J�p�$�in�1�E�<X7�CH3s�w�/��#����?pSZqhSA�w�{`���{�]j��WoF3�Z��s���d�OU�f��$�N��+M-NGv����7Ì.=���NL������э�	p��a^J)���J�O��O_��w�������/k��[{�*YO�/eY^���1���G�z�X�2��ڢ=�y�����\}F��v�p�N�miQ��~`�Q$X&7��$���M��rP���Uj>"��;f�E�(�U�t��B�%D�blFa"�zd��
Q�G��Ϻ�$��~��
 >9�Р���Ӏ�ao�G�$�X��T��%�v�}�3��gt��Dɝ�}�$L�S+�J0�}�H\�ǢL��w{��w�@�Y�Z D�����z�fhT�R��IS�uf������(��|���D����\�����S�f�ܵ���)ÔU�wN�i��h���W�i*Ƅy�xY�4 ��5�e15T�WY;����᧍����D��.*� <aW��� o�	��d��6�%X��`gN^�xw�V�n
�Mt���
bV,l�ben�K,Ȯ�j��Sg����HO��q@�^D�SWt���G���ҷ�_��|�`
�ݎBI��:����l��J���C�,ԮNBLn��̊�!����B��+vK\ϯ�����"9���oz�#�)���� ^�����k9ɘU�V�*���sQt�@���֌���]n�����P�ݬ�WX�� �+n����#�_ �!�=�
Oj���F��-WF&i]�1���{�r*?P-Pl6h��~�j>�T	�Z��tF�Z�LhgϦ�jS^>����4ՌO��H7��T�Ps5%�e��k
uR��?�w?�n������O����]�Q��Ǎ�n.iRC�BUv�]m5c�OU5���13W�#
T*A���r%����o�
;η��P1y`���/��x�x��RK$h��<�K�u��S�z�Zz�j�7����t�a$2m�T�ПW��<� ڪ�Jʙr�a�?3ٟ�_�Myw��l�0��HR��*T����>���4l�����sZd�������\FH/��I�f)���t#�NW���BY����#���!��`��B��R`n�?�4���Nz��̖���'��Y~dg{X���2V��ž�%
��^Q���/j�7�s�Z`41�Ƣ���>S��B�G�a����q�ҥ��#�3|�'xg�Kj�cS���i0&��B��N	�Dq�B�	����%9��-߹n_�Pĺ5p�d̜�P�M�ܮh;wR�� ��Y��,;��˛�!H��v�k�ȩpU���B��z'G7pf�5ث�/Ԓ�1���P��'K�f
�����ʬ�pxGrlo6���T�JO�!�bn�lkDI~w}|Ǧ,��,�5QΏ7i��<2�����i��I���Z��I�,I�8��~o��ս`��&�C P�-|f�_�.w�
SU�XЋ�'�����A�`�Y8{V��/L����cdPz- .ZW���Э���+�!��E�9�J��c��׿&,i;߮Ǝ��G�l�C*b���$�@A��B(�G��!�{Flr��?PZ���d��rw��/	�D�V�Fd|��I:�(g
��νB�敏�7��=Jb�+`�+I�8#��Q���dqI|d��<SD ѕTň��� %3m��*�.�� 
U%U�_fJ�t^�W���6�/(n��7.9=NG ��љ����4\awdM�Hh)����No<�89q�S;"�	�K���)��0��΋�lz8=�$r4�n ��å�h�.�=�ӈ?ͨxʩ�s��v�w�C"�}�������ɵ���-ɱ�f{j����`m�a�M.�Cy�b��aY�&���RD��,
JZt����^�@�wU��x�,~��S���UaM�����+=A[�>�����I �@ƣ�Y ��j�ŵ����aQQ��F�� �
�r��ʌoQ��c��������W������ m���qz"���l�q�Z�4�A�>��C("a�X���J=(�M%f����]^OU �������(� �g�Nx$��7-\"��Qq��כ���2rhfN7�ˍ����4K�ᵣWe}�;��3�����~E�;Z�F`�$_+��N�6R�TN۬���'y?�:-������f]�p滐/?���_[�o\����V:`���F�ʵ�*���g 1+߂ ��.>�孌�=�`[��$���	S6`�?rN��I�H0=*m�����G�E�e���^�	������N�<�-L K�G�^��ytuS}��9��/�[��}�p+��YAt�)-̄�p	���*(�����
��?����O`M9EK��g�!pz]uɅsV����E`Q�1/��55���1�78;�̬w�ӟ���v�i�Hs~����k�p�Ӵ�9��D���`ч�93v �Ƀ�;"��{U5��/p4aW���+�MZ�^�c��ˍ�E��1WC���f�CI#p��PP�,6s`��<�y��@0xU�-7́�j
�BV����c�w9̬-']Mx)SOK_3Ig(+����OO�R�	(��2��c��h�������:őE/�O��k�>݀��|�'J��f��yցD�C:��Ëy�]��H	�t�KwU�θ�xw��Ѯ`$����&XE[�^}��.Kn�"Ē����r����+P�SB>W��P 7<��L���΍�考�?�'=#��X���bF>@	��u-6w���mͰ��� ��`\0�[��+H�Y�\*a����~���]�kZ�0�Ъ�:�Ï���[I�n�&j2�o�],���[ʙV���{I4��f1�u�$�q��,_۩+R��@�l��R]��~�4����ݓ30ʌ	ޞ�ݑ��sK�i��������r�MSQ[���59���p�Ή6���w��� ���@�Ƶ��;��>�Y�%�`�v�=�H3ϴ���\�lw��ޤ������r_��^�k|��Y��=�A�0v�9�З����o�����aP[�'F�;�T�y�,uFq��8,��,W�V%ᙤrP������h={�AٯNKa<�g=>�R���St@�
�W N�4�\C��X"
�,]	����x-Q�ZT�9�0��!��$˂�L��fv?���K#6�_$v�YU��gB���b����\H[.�	OG��H�A�_ ~�.�d���RL^��z�S��R��a��&�?���,���>��0�y�z� ��t�P�?/�Z��f��@Ƈ���,�%��o߲� �?�����F:-��h�f���t�k6������3 ����m�z��������ڂ �4�\�ɂ���� �bv���h6������SCS��dԬ��-�@G4���B�_k��N�V�膇�Ս6\kJZ;�V�N:� �3'q�?��6x���(����?�Ӳ ��^VA�O�����b�m-��J؍�}��b|R�. ��s�1n�:�,Hgœ<�ǳ��hQV:�w�m���sh�S�)6�埦�PI���v��=�i�j��;@ɦ��V�H���N3��h�G(�5��ޛ�(���X��3p(��_�������K�S꛳���;�-`��l2�n���)<x�����KUj]��|�^�KR�e}'\���2}������]�ƃP��-z, ��@k��r��r|}�r�F2��qz���̲�� P�:��n��oSݱH�7 E�*_� �D%"�,���C[���j0o�i1�=����c�M�>1�åH�$����>�_0�-�����E�Wv��0�������=�[Ȱ/���UO�y����n��#�m�
�`��!R�(b:�$��ZO�毾�*)�vaa���9��[���]_��B�FD������<R���/��H��kAZ�F�=��T)p�/��&k�먈���c�a�xh��D$��	��&�����vf����W��K2�S9�ϻb�Ǉ�ߨpRތ&��կ����
Ѱy;W7��%�-got�Et߃x����H�-�e=J�!K�fg�>���;�=�B3Hg��g�{z^9 �+c5��J�[+��wi�?r��GqԥВ�|,��TMt��e�T�5��v�6U�Ɯ�)�wy���SO�Й�v��{y^]��-U�-L��)�~�S�����/Jkk�����gpA�H�+���ް@����[?�?I���0��h6���M�@.��g�9���>ۮw&�:@�ͅ[8h;	�o����	e�)�`)�!��-��'u���քӇ�j�"��v��2�����"^����\K�|�9�T^�[��b^V�ی�h�Lv����K-"\yW}�u�3���LV�o�±�ľ�_�\����D">B�_T���\�  �7�\�Q#5܇��O���h�c�m��?���x���#TB�ؘkT�X������8��������D%�_8�j���l^���.�j�m��X������6s�� �����@.�����T��SA;4�=��%�.;H!�_dJ)h��2'C��
��G{�2�!��"���f�E|������� i�hw0Lz*�D<��d� >1���
�������ي���.��ks*D���A������W���/����L�醯s�uV��>^�^ި�����C��X_����=�/<tk� IJ��:2�|'�
���j�Z�NVIE�$�b�cG�&�{m�\�&����f���E�'��Lx�̬U�s��������lMK�����4�V���O��)�|��ǡҧ���(�E��>�o/�����ҷ\�*TM��I��{�H�Yf����	.K��x0�����E�4tQ�d
U�)���HD��d�-�PK~c�HV}]�kG��^0��v�yj� ��QZ��;)�K�]^�Ӵ�mu�fʹ����~n�S�ݲ�M�A�p��ʼo�K�(0N�qxe'��șU
����PlM6���f��&��ܳ�ýBF������͒�6l�|��:Q-}�3Zxf1�S��I�����o��'���M�lA�]��k?�Ꜽ���z�`ъ���"P�@�,�����^!�n��7n�xu�k5� �L��W0s��2�sS*�Q�2�o��xF4g���o�~�7�0N]∞X_