��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#�����~H�����pl�Um�v:��L��Q����;�~��?U�b����1�w���`� �2����:S���Bq��6w*��v����m��<�,E�H����,�b�M��1>k�^��&�SV%�n��b77� ��������m?��8��O�07�����v����-��Z�h�-"�f����v�Lk��em.������~A+@$���V�����z�K�Ex�;Q�2���Ij0�P~�ZR[�J�>��As6�a�!9�D0��c7�w�䔋G���ITwߦ�8k��i\˧�Ǚ��3|�İ^?��g!��
&�GCW��'W=+4=i�;(Eq��;�1!�jE�O�UX:k�9�M���L�Y sƑ�~%�{ݽz�}�poô{��n�Y��%g��Dm��^Mifߴ+�������P<�l�W���o=�WƔ�}��8�@��?�`f�n��j�P��.a���] �/ �Ӊ �P��)����'�&�h'VcЏva���2��b�f���z�h�%��G�B�����ؐS3��6p��"��Y�)��
�nP� 5�9��N!e�`��1�C�5�A�:�أ�YS>�j�3����1��eL��� �{�9���wT�C�(�B:34!� '�iڃ�7��#��b�.��Wt�C��S(�������!04�.��a#�@�3�!Zd���p�{���N�qy���΃g��Sۚ�����qUZ>`�b��I�d���Kp|�#���?�z,��6
W,/P���R|�����o8�������J���V��7x;#WK��c�r��(��(1���k�ߎ�Hk�Iš<&�
��JU��^���re����9���6�(���3"�c�O��&���"8-��)��=`aL�A ��&)���,�+���u1 ��
X$X셻łT��<ᨡ5˹�3�Ŀ�V[�s+�N�i������,[�c���@+��Ѐ������Fꭵ���+h�l�1�d?�����O�-yV�����/:�N�A��4��8����@�<kp��l��\�	��\����!@�/�ߞP�8W��I�wG��Z+���-��Se�:���5�V���B�D��"�Po�%������W����-k��
�n��q
9QdL ��KK�zd�X�~�������>YG`�Z+�]����F�t�fv�\�9g�uo�Bp�J�V!�q�H�YPBܮ<XRejO�/Sr�$`O��;|�Kn�课�5$�(O�d�h(���)Sx�ThU�e�!��H�~D�ܘ�q�˪'�LI�y[�q�z>�Sѝʄ�&,��;�Ej/�P{x=���b�X�$3X_Tī�y�c��O���#S�\%-*D����C�:+�TW�X,��v��D�?^�T����O	?3�u�]~2�Z��dP�x{ʴ�H}(����C/`�X"��U�%�d�k�~���$����  ��g�����ܢ�P�ő�b�թ�������`n�ww��)|�����A.�.qz���:yב�#ىA
r[[�M�0�kݖ�f���6L:��r�pYy��Ey��כs���y䐔�RV�J³h��9A�.����n�ٝ��j� �c���^�7:+b���Cg�Z7��* 3n���M�y T�@1���(���_�|��K �53�ҋ`��.-ġW�3�����.O��z�ey@n�R�CΚE��
<�\���/f���Š�
���8�{*��f��+�@��s��/�+k1|�ݹ��(����1��z� 	����ji�%��}����G��aH.��
�G���/|T��4ag+�8�z��#ĳ�5�w���f�#�:0K]<T-��V��|��ک��M�ů_!�;�̪D��L��˦���%;��"���"�!��ԓC�Ń��3�b�ʄ��[i�w�GX��Y7L֕5��_T��9�Λ��9�<r/2J�S��lJ��}�K��.-F`���Òlm��[-t�1���
�ƪ��t7q�u_`  C��g]�FQ�>��X���������fF5�N����1�J-6X�>��[P����i?������'k���j��ZY��fVR2�"��ٿM�N �o��O%i*'j��c�����u�I��f�Bq�+�ʯ�/��+�Y���,klC'B��ɬ�N�;��[��YB���@Xal��6�h�k��6(_����k#�{�5a��FM��{oE09��W�1C�l�����YF�|L$d�X��!�� ���\9f�}-���ȹ+���礰��:K0�l��C�8���)p��CLPm���V��mN��_��
��;���������<��ĥJM��[U���KOv�WM ���4�|~�ׂbv�s�r� �#f���H���:eT�#�Ú�x�"E^���*כ��̤h�!P�(��Ɉ�Z�-���JOR(m/���8`X��L�*���}RF�z�������4H�seZ��WB���Lu���+�(��7��S��U����{<!$�x4xޓ�72܄l���sgF��B�3�,)�ed������pc4�%l����r��Sc���S�\�D�ި��݂��������N��oëk�*�TI��Z_t�k��ir���1��D�3�~��i/\�/_jrMOqA���������O���i���;L~D�����I��E!�ϓ4�e �PN�a�V�Y�8���W� �êKd�؄mw,=�#>&��gͭC���#k�Ӗ����M�<��M�!C�i��G�]�XF�w�ќ�_-&8�9s%s��� 
0�g�b�{�1�7k�r���ι���H��ln)}d\��<��Os�	e�Ы͵3�
��?zr�5�$�/�U=y�`�;�\�Z]vq��܀(�Q�|˃�-Or(̰���>� 	v�/#�Yh��M���j, ӪU�tc�V矊5*B� L���xi6�k_sw��Y�%�N.-n{ßl�� i�n&os��X���l�:�ǘye�W���g�c��4|N�	O�ƻ:�3YgX�������g�l�J\�'��Y���c�_��i,�6�f���̌�1���"��U<�����A#��;�v�:�\���u�dJ}c)�����E��?*�M���_h�n��AZ��6�|�.cX��W�R0����tpvG"�z�Fb��o����|Yw�x�?�thJ�!a�C�����,��].
�/i�Oеˡ��T�'�HR�P�K�9]T��`�I�+�V���'C�sGd�ϑ����k&T0�=#e��*���N₂�j.�e岶��t��ƃ�hl��D�Qj3ī�������2�}�`:QB?ϗOް5��6QAU�7)p�5+�)L}���S�IT��`��h����!�?�F��+_i#��y��t��d���pR��w������d��;G��aA��x�c{�FYM��oE�E/P����X���rN�����დX�����U�D���%�:���Sp	팘5;�Ϫ�Q:� �~9#k�@i�$��F�/�|sC�QJ~���U���ݨG�?��|Zt��RL�ƫA���A��U\�t.}wΞ�v~�oe�BTI�3���M;������b�5���q��{�&W��NY�(ۼ�|����f�yT6�Fw�c��d��s������q7|.��P���e�	��+���S�����Ĩ�Q� $=(1v��?��Mݐa�F��<�r�y�*�U$��,�k�8��bN*�vv��Cd��B��	���#6+Nѥ6T��tn���8�����QG��:%����������]��b�e�2�|��n����VXr-��͉�h�o4�$ƃ� �Z0���h���'�Wt祈���s]���v�'$%(��ruC�����@=?iD�d���e��
��j�͚lJB����XUY+Y�m9e��J�(�Q)�����m�N�z���#nH�?&x ,�ㅩGe�T�+P\���3G#s`�h��b#g���V5!~A+������~�����d�H�ۆTI�a�e�8�{|�2t��6�4q�I�,���g�/����zf��\�+�E���p�#ִ_�K��	�C����݇"�K�\������%Bų�	],'����`���J����mu;Ob�bJ���E�\?��ו� ���rÉ-V�^�_�+���i���>�9�����TM���ٹ�?1�ԁ�P8��32S;��j�2#��&,�ۂ��J�5�A�r�įk;���A+r�Nū�bi��ͶF/s�Jǘ^�����[��T,�+X�qj]2�)�7��Rt2+��������?��>!_�k���7YB+��W�OG��6�Ѝ�i�_���F�dB{���������������9���'$Rb��F�>:�d�3�g�ρ@���X�j]F;LvJ=���Y�����#\K��*���_[0qŪ���\�������:�e��)��=�e_U$��,��XM(}��4�Rq�vG1\�K��ὤح��F�z�k�5+E icE��L�Q��]>9��L{Nr���P1ђ��%�olx=�����W�
��+(�f?�R�0>��Z����*�x��2�g�P�i���iHU�$��,�/�E�I?SBL�bP�.�;������+ ��T7򮟒_��VV�I��-~�F�u�dc��Q�|��0Q��>g���/�T~5ε����Gm��x3g�yʆ��������>E>����n@״\�gs���&��x�tA=�B�`���	qzVP�.9�vmNFYiEq����V�X5�G��a��a�.C�ͭ�1<P�qC�T��L�m(2�����:�@�ݰf纼&��X̖�G��Y�3t�5��7�a����W�jD�	��x,ېW.������^\h���v����9#�#�����;�o���Ux�O�+�V%w�*��Z���R��X��凨�Ygu���E[Q�����d��>�Tx�6iS.�S�ƴ�*�[ɚS0��7��(YW3:�R!����*��7N"�p(�7$�Ħ�A�>�`@Z���Ҳ����5;}��x��6��a�����`B����f���qv�)�����LGR���<خ�,/Q��t��NX��Cl��ٻJP��>(�c�햻���B�.�&3���Q��S���n�0���b(��N3/4��4R_�s�W#"���3g���ד¡� C�BI1!?���-�M��~N��D
UwY��| ��$ILV�W� L#t��ă��E�
�)A�@�5Q�+�;�Z���M�m�{L@��L~�S&��������hb�d:�� �s��Cz�aJsG���츤�B���y����e�zM�T���d:�����h�j�wh �a�&�Ah��I�KP�9��?^��*��ʶN{
"�%'n�v\�;�-�^N���g��=�T�B5���� .����/gFQԿ�L��a}�&��Vm������<N�J��~W�'�1X(�&v���8��3t=�@he7�+�}���u$��Re���fOՐ�>��5�J��y�g��߳y0\�%���r-�ˋ��W��W�\#i
�he��t���X�a!�YCu͗�6�\��W^K�=�eJ&Ѳo���0'�@���X	�HVP[Lh?��h���m��Q>^]�	4����w����v)�)�uK:��E�>���ٸ����*�}��]�D�M-��69�	�p�e��b=Z9-��u;�og�+aF\�����Wi��7�a��^73��M`�a�T2����9�ҴV7|����B�Qu�G^�44��ۂ�n�������-RtԌ4>��)�}+��f��ʪ�z��}I�[M&)���,z-_Ϊ6<-<�/G����(�T_"[����#��nݦ�E��a-�	�r�IJ�*'���ΰ�N�_��H��O���Z;�)%�	# �`y�����5�8Q�루~�~�7$�S�H+���G��cqz� �������2Q�WF�a�����ZbA�b�'�S�;e<`��B}x>}���dJ�~h�H���Ƙ����&�]	�epW���W
-�!�2/wj�ՙ�MλB��qj�	��Լ�J���O�3�S����N�����ge��y.o�=��	��l!���M�V��V��<�%	/c:j@���������YqY�NFJ+�
ڷ�[٭����P;,���!d���X��{�AP�
��*UEq��Z�B�Z;	m�䳘7�	=���ɢF�Dhl�� ���#��� ���n��08�|w]*DSL$I���.��L?C/�
��K�+~ZA2-T3h��ƻ1 n��3�8$���������Ϟ���K�d�H��T,M\������q�;�D�ׅ� �z�a��8���'��5�iɍ�I߿ɠ`�����T�#' �>��ܻ��<J�ަ�.���i�n�Ȩ挾��l4W�G�W ���^��	���kx�b��l�~��Q�$�m�~Bd�FܷQ�Og�l�h�A�~&8�����	���`���4�^�x��:��t� km����n�u��e��,_����=��#�o���/� `���ѥ��(Y?�C���k��o�`��z��G�{u
][+˝Ʒo����lW����O���m�T�۳��1yX�(}O��dd�!�Q��`Yt8��f}��t�=��?2�E��M%���c��;��b�\@{���i�w\qIC�Q�a��#!t��<��`b­,�y����5~�H�ڻ���'�)dl��s8-��j&��L=�8C�)�[�G��+�Ms�ω���r;]��1?l��ڂ[˱b�,:͜k*��
H)��ط8_��)^D|�?���+��C�K�K��P֒1�X!�����{����蜢_��U?Z�W���ҧZqr�#w\�̈́ߢ_�H/������ ������@5�������dQ�-���G�u��L�7d�Mö���+�LV���"�[���d: 	��4l��B�6����2	=vV�.�q��'���.*��(����,���O.��^�ܭ�5��;�v���t��]@զ�{���@.���F�� �e��^tn���fn�#��Z�q�E��7��D���y��qt����	;�L���9����#��}kl#e��)
֭3AoTPK:�4�\�03-}�X"Q�Ů_�	^D��	!�g�x4�#1EJ��7^����m�y�n�|��r~��e�Q~�G�q��0f�
&�_��)���y.��W��c�f�oq:���Kl�W��E�,?�.�kQ������P�a�P��>���O�)|�I&-�n{��ߺ��y���Y��!?���#=i���$���ra?F�C����w���AAN�=�s��֪3�
��Eز���"B���ǷjP����,�n8��;�A���Ye�km �p��P�Н��ƒ / Eb�*������?	�;��d�2��̋<�����R�5��1	*����$5�wj#� -�u�ؔ"��=��#8�sA��3%4SDh��y-�DY�^��E$�Q��E��|�ð�����ih�>�x��ob�Y�4���ԝ��p�8Z�@
b ���1!�ű,do;i��!����_��)�W�WN�	��8�3Dh" B�s��X\E���_�!|��lX���!dz,J�D�]��Nxv<��7���)�(Go�[�~��I����r�^b{F�Z"G�4��80N;���c���7g�Z����+�����>��{��400x���Rr���I���}�����$M)o^t����æ�xTr�`E��	��� 5����+�x֚��F&a����˶"��*\��������HI<m~�ե�gI�CH���2dp�S���8�_�"y�y�� �;�U����u��L�x��R�|m�\���'���+ۜ�-�Q(��^��El=?ag�8�s�_�e&�v�#I�����S�xI���}a_�֦4p^�!Y�
=����%%�8�<����l���F��稧K��P�eZ|�Go\+���{���v�X��	�k�b�5�Qk�ȔO�G�	N?u�w��Ce�P��FD�O/ZbN9����Gcn�[����k���pȕ3jR��/m�h���21�:��~Ԣ.�n����O4-�����)8���N8�&�'6�/"]�&Ejm>Q�ch~0ĺ ��Ά��:�`�!ɺY�x�3{e��!<g�9��ؾb�������.��]�R�vɘ��W�#�������%��0�u@�~��W��.��(u\�pK�AZ/.��c.��Ř~����Jr>��#�7[�)��f�2�$R~|]�w���{�#�='�����7w��@�4`˛�(oQ�uyc�*x��eYd�Byֽ2�"Ԓ�FӸ���F]�_�=�@��?jEK���t��c���;���(M:}����u�¥p{M�J�ģ/oA]����;�׺�}Ė�����.D	L]P����s�es�.2�c�ϧJ������!vA"djeh�I��dX�$�;�2�+?�Dlj����	ar!y � �2/��C $�2��ǈ�4u����}쁵\�o@�ǵa�����:�&� !Т��b�KU�)�:c��՜ScZ�vr��֧�OF���e��nl��l%z�G��Q�������7
!�-�p���=x��
M{N�`D�Y���[�t3fQ*�c��W�8��s���w	��H�o�����#e�����oA1���"a��k�x�h����h#ȍ�땒N���e�y�M��+��f-us���H�iB~a営;��W�\��u2�{��}I��3���3_1��l�;�=*"c�G�Qkm�0S.�n׆���7�7BX������4�5������"n�k�DoX�D�S��!�LRKꮅ}ކ唃��Y��O�Dok�K�	����C�ߣ�ɶ��v�0zΡ+���r��=��*�>�L&�P�>±I�9�u�G�<*k�)���b�(��v��?���q,�(N�ٺS��u�w��8�l!�ANz��#��f�}��=z9��:9J+,OR1&�q��@Dlg9$ָm3z�'E�E9+|ԟE�"�ܼ���J����d8c��zy)7�h<|�SE���u�1��3f���d��q�ucY�亇y�����N?7�ɣ~,z{��N��p.�ׯ�Q0]Q݁�>���h�t���i�EI�C�'��� �E`�aPÅS�Z�|�pf�[��qɜ���B�|mp�TJ2+�#5qmZ����d]K����iB���fe�۵��T�3��:8M�g�0`�_�*R�@7�Ps�Ap�ı�-C�3�P�nX�i{��sZ�<��u��F���{*�涼ӓ���x~��}_�}�t)� ˽��S��rǵy�g��F���8S(Qy�y��t�s�4:�J4̲����e�7?��5-[;�6mqMY�TPpY�q3�����^�~��b��T��*n���-�IJ��B�Z�q���8�뤅K��;K�Fo��'�R�q9����� ���J]#�Ղ�@���������?� �q���}Sw�}�9��*X�
.��Ȃr���wW�0SU<�a<�g��� �/A�<�4�iG����I����Tz�8{A���G�'p��w��t$d&5�\T>o5�3�4�
���+}?�rY��x���rTz�i�b�M�n�`	q;�:dJ.�L}2񅻭)]�5�6	xJ�aHq�ri�� 2��V�P$�DpU��v@6��e�5}p��#�\svў�6���C��qn�Fx:D5���9��Nb��.!�����CD�i�:E�b_]uA�y��cUr��k�QP�#���2�/��O��_�Im��1�BNy_�쬚��m�L&��G��ԬB�⊖��Wh����7$ۆd�/�m�E���e �����{ЌQTy�K
�-O��=#S���,"��w��w��*��8��<�ͲD����chb�c:zȶ�i���T�+��0B�:繁u���0��c�`�>�;�@���w	3f���c�_�~"z�ͩ���iK+h9��i�=�O\}�v����ߧ�D������|%�KT54W�o_��w+���fP�
M�^u	��g���^,q5\\�6�J�y�<[/5Fqw9�s�_�sq�����3�@�4�ȫB!�6�o��.�)��[�Y�RW�xg�ˤZ���?ȸ$�Έ���Ulb&r^����V@�y�ŷ�ۿ��r�gYj���n�%��V=�F Z��f�l�wG�g�%R�J���^���:�٪�t�Ma�`�
��%bd��=G�9֚x����{����i��nt���vW@���@v'� &�Af\����Ob
ږ�W.0������/���Ӭ4�����7�4h `Tch�7��1̶�c���9��@�&&s�GE������_�Ҏ=# � �	,�����lJ�_X�ۭ⬕��J�\4�Aa��,ZP���3�Ae���R����N�1�Z�R��� ��E���Y�C�:�8^t�����o��B�Xm[�����#�w��	���̨�!��Wf���c.�?a8,�H8�@�
�(�o��?�'��W������X%�� �5\'�������]��0���bv\� �zAVاu�L��p��o�D��o᭑F�Ę��M�c��~˯��%|	9<}����%�"�qϺ�Gz��2�"zm!�(�1mD�f/�c�%����D.獛p"�-��8�1B!r��#������D�
����t�`5�F�g�,D���5MR�(v��fsF9p��\� ��p�b"�A��l�m"�P��;�pF)ülV�9,��u��1AA7�#TF�	�p�48�r�S]S=hb���6]A2�P-�>=�>�r#�W�Վ��;A����㔘4K��U��F��BĪ��L�Xbts]�8'�+25_��7v��ۃ��{o�)}�,z��0/4����p��
@1hy��;7�L�j�ُ�]��b^�S�-Nѿa$}k����F��Х����}0r����&?q5��$r��]:e���	R�+�[^t�f�4S���֐
Ax��w�����W��*�?q�10M;u$�Φt!���E�E�a�k�������)�+G��r���۝3e�|C@�s�4�1�:{�	�����w�)�$��a98x������`��Hw�>�]�X*�Iʶ��ES�4@�L��Ȗ�O��)8o��P�
�w�jҭ&�X��Pmp�H�����2��ȏH��D�%EP�#��S��A�˧��z�eU����R���3�<��k��8�T�T�4�[�6���p��t 5S�:�_+�u�8d��Z��C���˒�����"vֱ�&���?�8lD�>��-i�_��F�^d�%��э�yLv��BA��&̚E~���*�Po�o��o��I+�����f���m�2�r����#x&�<<ZrC%񧰹9Z��ꣂ����S�h����a���s� 6>D�ʬ����}۷w<&�e��iU���"��\�d��We�K����J�D�Mz�/�&R��.$�v4D���T I�*���b��g�",R��*?J�߫�ZC/ȢG�8�!sjt�z,�'�d{0]r�;�^[� P�D��'v9¹�߈�����#���^G��0����Ā��l�a��;�i�)�ؗ��	�e�z�CӞ�x5���H@���Z{�Y��Ҡ��]7(}�V�(�<�_�B��8īỺ�f��I���^IU�=�A+H`\�7[��b��	>�l��Ӛ�g[�� kJ������'����0��s�܄�c�e���0_�Ю:������p�d�$���B�9��)v�1��_�ؽ��&*`���藣f���h��ޡM�fvClYk+���rH��6x+O
+�hnXJ�(删���rU+L�6L�E�
���B��>����b�v�#DU��<�}�h`;���ܥe�rLPx�cإYF�<p����ﳅ8e����`'�I���b�Q�F,Kb#���E�Ŕ8�����#�e���7�٦�f%	�iU������G�s-W�z���e&jr�-�'��*�d�/���d�?YO?{��
�fo}���֒��(.u�A�0�&#H�Kx��w��Ծ�i�@����V�S5�NE���`R$��4B����/9^������*�yܐ���w�RxE�3�+6��S !zF'� �`�|�����g{;]�QI��}�������Y��p2�[���_��H��;�
�dG����v~ߪ�`�١woC�r�ظ�gJ�T��:5�YvQ�<G�k�ȓi���rlpF�����uW�~�8;�R��Zc{~	���'�/�1)�?ίRI�QO}���^G�� �o�ޅMo;/�qƎ��F-���ſtmk���.Fw�z8,Bͮ���|S�� �	��0i�� m�ˋ��yJl�~�f�O�����F6^���R�r�_������c��F�+��4I<�^]�3����\���F,�q�N8x���̦�^���JΧRT�嶀Қ�H<W�M����\�޺h&+6BL��Y����f����c��|N	�P���d���|���<���@���klh�O�c�tM�F��@�a�H�,��	H�+w9U��K�"�Lh�������b��^eg�oN��S��.��ܞ[�of�!=�WA
ϙ��(\�%��y;�ݼж�=O��F�?q�Sb��=߳�h�ݿ8�׋T��a��
�A�JϾ���Pl�s1��q�!1pϟ�A�-��4�>xTq�qw(ԙrk+���O@�w4o�B=�IE+W�(��q�):N����c|A��}]�Z��c>t� Pc~@��Ⓤ�!��G0�Yڃg?�>�ݻ9��ph�T��Dg<-��O2tgT4��S�L�� �8��s�B�����G(DyO�m{�j��X���R��w?���{Fb?SqN���y�� �I�enV���\��~� �kl���Rǐ���I$����)��_�h>�3������'�ų�I�r�U\��h��Ϊ����HN(?�u(���Q�'{�d�� oՋ9c� \�v�
�6�EH��(����y�[w�k��Q��ڳ!�0���(΍����@�N����QZ �Uȓa���aL$N���Uq�<���e�	��C�����?e����0�2����3�$|^�ª�r}l}���R�fN�\��Sq�_ ��}Y
G���څVXE-���Z���`�һ=hPw�Q�ݪ��Ik�F;-eؔh.!F�l��V����&M�Kb����.�Ѷ�R�L�r΃�F��gc|"�Ap""[�e��+�0~NZ�%h#1̅�U3l���o�9C6����Pe�%CHQ7����rZJ�"�=�;�\ͧJ�G|�gn_�����.!�fu�\l���)�2�ʣ=B.��C.��BX@�c�������a�g�rS�bbT�5�u2⋑�)l��H�*K�,*��pYhot�9tb������|̘ iX�Z/�E&���5	p��19i8������n���f9IPU:�jW4���c?���5,IK���Vzb[7�P�Qӣ� pKӯ�AD��F[��|-V�1J�X����a�;�5 [�=�\|:��
Z�F!X�'�g$_����F���=��W"�ܖB��牵/�ʰr��>Wk���]u̱4ų�p��g�e������]ylHC�μ/�2P4�	K�5=��(��vU޸�H��[(3� ����eɛօ�2�dS�l��V5y�u��[�F�#�&�6�1Q?��B�B�V��^�in�¯ o;SF��4fJ�h-���>m9D��y��'�ɵN����kݞG�ڗ�e(v�Ts��Z�X���n�r��cW�K�yG=�dW�i��A��~�*�`�,�����KH�ѯ��d7���=��եC��a�k�Ѯ
���Ma��ө<U2o}�&�f��P��=j�G��{u�!��o�U-��F����#�y�'p�qz_X���i*r7��]�=x��=��o�?�(B����gN�����F��ndp��X�[�Q�5�����n��̙�_t�L�y��f	&{��	�"�}�hD�◚:�-|���N8x` c�.�NO)=(յ�A��S�`+Wg|�1�y��݀"���:��f��
D����b;�j�K>��'���F�e�OF-���@��4a�A�W�R��ݿd��#���i3g�j����3�	�"g&�lO�A�2Վ�N�D���Yҋd���<f����*o�!�	Y��Mc��&?��6�����_i�:'�m�]��s�_N>3��1�hy�:������e+C��p���Z�3!$#����-͂s�|���M��l�qH�Y�d�?�f�ޢ�\�F#e�&vq�1�"/�xi�B n�l8'�|V9��j��td(�ǺA̕)H>�ʉk�tR��ssmxiՁUV�Z��]W���������t��1f�9�Ii�K�D��98D�}�&�|N��Ň�����<D��-3P��#<�5��j&0l�(�{��� �٥\�y&���3d}'��/4�����_�3�|�j���ӎ�t��_�|cQ"B�g.,�@ɾM�w2k��*r|��Ÿ�N�ƫ߈,��ub�A��R�����+	��AS0�bi_sT�e��ʞ��ǿ�����[�B�u��3/^��H�!r�ڄ��##i�R<s�;q��G�_&ݲHoע,%�Ȭm��������q���#Ɇ��A��,�n(?��*�D�-A+��y��%4D݌�Ŀ��R�fI���=fZl�	J�"�:7A�"(���v��(����6�^��a�h�e$�iÜ��ҕ��}���P��gmk �K����[2TlN������5�puS����l~fɹ���Ϡ�5W�I˫�
%�8^i��7¶�O�<���}��j�|a��2�yU��@��ʥ�:"�f�q�-�*D�M_���c �02,_�z4p p�����/u�n�7���$Sepm��x[��3�V04�*�D���E���M�3}퍛4�l{x-w�3n��Da\/J��\�*H~s�3[��mu���޵T��ɳQQ����I!�
͍|���B��vڈ�W���J�t�F��M'_���|J��9�t&.�;�9'���o�]�F�%)�<�g�Y�S������:D��M���S8@m�\�l�����f4���
�k ����AP�
�Hg _�;�%�jC̴���� eT�cU��#���K�$�;?fx0︮5�J��T�c-$�]fi~f����⡾R�Q��Y���^��gW���`�'i�p���8��5'`���Ȳ��5���m~D�Y�����Mh��j��]u����L*�$�cf����+��S��Ԇ�wq�fQ4�YT�����x������� 5G��mO���,�ǰ�y�L%2 o�ߊ���)��u�t�^�s �38��#��Q��9c����� �����]j�.���sK�7����S"�gX��{F�f���>�8��J�����&B���-s����C��O�;�i�Ń����?H���K�*�P8E]H�*j�S�4s퉜s{��-/�x�W��h�~���C1���E��'oo��ÄRȇ�K#�V�f�*j����~�����pu��IH����Q�ߤk���[�\����2||崦a�����d��#^q��%�1ƨ�U�T\���ݝ̵�h${s��sc	O�&�����I��k\�S�ƨ�<����^�&�a]�_�����]��7 ��oD�˃u+X���"}�M2qcչ�F�$����m8%y���8�!{M߿h�^N�:b��_�2�F�'��H�C<b��T�.w��
��L+�d
��sj���?���*|���ˀ����ʅ�����S�lC�9�m�n�㟭�&�7-	��������9���^j�%R^�]z7��8.�bgr���t��tcq����%i���D��1d7y-�w�8�w�9�	��T�sX���>4{i�Xda�nn��=U����p�؅�cޛ����8�y�i�w�L(��<O���:1"_��T�����A��zyI�4G�'��\�yAG\�(/W��'n�K����.�D��F ��g$���D�p��N��_-7Wk�P=k8ى�f�H�9)�A}*�s��:�4���M�-"ư	�b��)�_@�ÊSh�%����5/��p=�+i�b�� ��c�v�D��^���:�O���g�����aRi('k�c�����;�����'hЂj���/��G3����^���������5;�Xmx�O6�6P�~c9o��羑p��1�E�p�����+���"[�d�@��c��X���V��֩�f��o:<zf��24�@)����B1�d6��(�)[Bg�i@R_Q�f���@I�[py�����m\��aV�����FI�}=+<������<��Fr��[a���M����>~�.���wFa��?���� ?|���/i���<~�Zk�4&Ɲ���ӱ���mwO��������d2��)xʞ��uM,�W&Uh=6�k�8$������q���u��y���o�qݽ��Hu�<�h��lu�o�6B���:�O./ڒ)p��܃�*���bt":\�p�;2���sٛ )�`�X]fhc��H}_�IZ����-��Y�����usp�ؠ��b[A����17&]U=�A�0Q�N�
o����/��a���$_U{:�7阣�C451y}��rc�f�,Ǭ��N�=�61��1�{�����+��n��ͧ����
I�^\6L���*r��?i��Z�Hu:=�=v���U��T.�p�F���3�nO��y���ҙ�;��R�{0��[��`!�5@�9U�vu�9ZK�$��;�Z�g*+͠�7qb!}輻R�p��^ڋ,-ݴ�*^m�u3��2Q�*Њ�Lp��^x��6�|���Xʟh�<��/�!=Ȣ���H�<����i0�@Œ�SqDG�u���xJ�H:���4r ���F1�lw1ud��Q����v�N��¢�}6��(4����af�HZ�׳��q��ruba�e��7i{dI��ɿ�˰�����7�]�Ahs��4|��,��ܗ�J��N�q,�76�� �֫%��]�Ϣ͛��Hg}_Ӑ��+��� ��$�IN ��KyH���֛B�Cc8��B`g�����qV��^;��8�ZHU�i��p�G��5K����Q�}�v� rsɈ;L�%}�by�x�YI�G���]M��i!�
V�Yǲt��x���H�h��o_s�S��9�D�j�-��m��\�o%?�=7�F�%5��l�gP�L�:�_�>�hI�3�f��K���Ќ�HC$u��c`#����󪵠Y�I�����qr����zf����q��El���CՕf|�4�KFx����3~��d�{޹V3}�ŭ�haL]p}�k�M�l���F�FGC�����B�_�V��>I�b���|Ն����xVΩ���*�̔��qJ&�=<�j GϮ;A����Uh�1R!�Z���{9F7oV^<`A�`K�>U���71���KT#ɇ�)�uWfdq��ׅ��*u�h�̮����?���<RMJ1	9���j��"uq���1_�*����%�-�[·��F9]�ן(:�0My�|�sB�*T�p�ơ�ahy	����9)!F#�W����~b"����q��)8J9�	�%]��Ro����|A"{�M�Q��+����2p�d��)���ofe���EЭ�C��X���B/��8ޝtK���b��7C�Oj�jG��o�N���-�K~�4�g��r�M�$/Vή �̘����Ojfz�+�6	��p��+uN�qqcJ�m����|k�d���
�t�S���A��=�������A�U��o�cZ)��@ᕀʭ �����~~�*c��<t������&%�j2�����>j���e���;OL��O^�9�WaI��%��u	.F�P�Bݨ(��Ȧ�dK{�<?	w��a1|������=��~�j9�mkŎ��Q�b���s$%S�[���O����v�-�xKmi�F�VHx�'��lS��(Ck).�Ȍѻ?����!���<,��G�Dx�A�t���֕��n:A&&)Bqe�m�0��Cj��41t�6�������~��\��K���p�¼�ma:^���4û3z?��/���*9�����h��n��- >��E.�'��gg3��85���ȍ�*p����	1����t�D����I
Q�m���&�W`�<����H�>J�=8g>�{b�����QJ�<j��4}m���o|f�o1�3i��G�%��#c�\ԼӸp��'����u����"����-���.Bc��q���}o6�5�h����1���z�*V%z{���^�p�a�
D���eڐl�io����7���ُ��]�,��K&N�Ѣ@bi��7m����0���������ad�Q��9�*0�a\ar���T}MQ5�nÔ
�$��g%�R�4/^-�O���M����<!��٨�|��d�pi�j���A��ݡ4� �d\���m�`YN�	?��UV�&�GK�u�/-��Gu���?u����\�2}��)3����C�B/��g�E�U!�dUPޣ;O�14@�pAh��!����ß+�Ω���i�⭔t_�h�L���=�:�vF�j��	(���}~��)�3p����(���+�x��,����qRXc��K���ÐU�mt�Qki;Ƣ��c�ഺ6��eh��F���o��^�U�	LQ���������d�V"�+���d�:r���c>��[E�����|��L\���������6�a��0��p�����U*o����"����X_P���q M�ps�m`φ+M�.�����Ouco?���pDV�{����Sg*J!��v��p݊�K�B֘���k�j��b�C�RS��q�J#��3O���Rx#���[uP4n1^!G�Z��u�v�YwkP���l�[A�	U3��n�o�ګ�!|p�ٞ:i����-�U E�q���:|��됝vq��ܨ��� �VW�t�TJ�͹�Q��3+�{�ư����sPX��0�4�JX2��n������K8x�J����8Rs[͗�1k(��Gс��g��Q���Օ]�DT=j!^=;��%XM�/��>��ë���.1�Y����ol���K�wSl�G_VX"�H�ޗ#��H�����V���*�H"��N�VF�U���܆�r�13Q��翅 g����Mf���4Ѐd��?�*����u��\<�A�V:�EIBi>��LB �� �و��s����С��eӜ����	Tx�#��Bg���;?�Y&�p�Hn�<�݀y9Je��pа,F%�<���k�����
6	H���-%P	�m����^u���A.��J㻑k?����Z�0ػ��=:�Մ��7��/G,����C*��-�f XE�)]�J�L���o�.V3z�pS�w�\�nݛ���y�h��:�>��{T3���8
�խ"����6?+�
�X��鐓�w��r�N�Sr!jV(������g�h��NZ���b���=C ������G��g�5��R��7m���;��|9��KZj����_�Oah����%�N�����SE���Ce����RI�J���Rr�0�����Q�S'J+Lds޸w��w�^2�[�s�̞�.��cļ3�����9%�
�yȷWъP�_���1� ��R�xA���o���w׈[������n��C����Tc���Iw@!D�0�Оz�C�Q�~l�֓k�V�--R���'��Tʾ��F�����u�*�e��nyܘb�ff������幁0���N̍��$�=+u�hB�RI$<C��ޡ쏽��۳�\�fѩO���ꪲ�O��qG��n^Q�T:�#�_�L1�9r��!E ��O��T^��%=O�QD۬��{x|pX�-��}B�
�{L�>K���sg%��ϧ��U�)��I��/������V��HL"�,�q�/�5�ϐ��@Z���5�C���oM�1wQK���<�R{n.��x�<��O��LU�֌?s�g<����u�Њ��7�'hM�ٶހ�t��F��g��[�*/qX"9|��P|$D�%�1�iQ>/U��'����&�%qxs©����t�ಠԐJ�����ϩe��eJ ЎC��X�c�%}1a�c�ǁ!�����=/��Zb� ?��|��Ysp� ��uv���XJ�����I� zP �yU�bu>*؜���
�����*�s	v���*(�ԟ�l�K�TIl�j�n6��H��Y��W�g4nO��]?���H���rDo[��Cf؞R|����X~���0�qq�������aU�$�_�8�6�ء�5Rɴ�Ư��1ܔ�d&��fa��V�*aW�FX>��"1Q,N]�˄�MCUڂ}U�S�!��9�۔��r$_�L4�o��D�t��+�P}):��8�՘�?GX��v��;D�������m4r�	�@w4�x���ʒ	��t����gځ�����Ay�뿐�1�����A)�I�/���O�;ut�r�/=��ʒ*,����14h3�D�����#���u,D	�)� �����<�������j̚W�1
wS�f��s<rH�!X�l����nا�	H��r�������"�55 Գ6!��2�8��,�r�o֕�,�Y)�L��6��S96�X(�O���TY\�n�t�M��r>�t�_?����9݀A2EW�"���ʀ�Z#bϜ3��@�޷����UeW���o̙�� h�i�=C[<�̋�@E4Kazg�87���r3u���F�.�&�:?\��X��h�:� �a�'�?+���t�5��j@�vV%�.d ��0M ht?Wj=p��KJp"��h�A(�\@�U\>^��Su�� ��'F8,����.}X�Y�x �Q��*X&���#�䤎e/�Y]�-y,����ʾ�)�z(׺i��ꌸ�Ɩ
����c��/X�}P��l%��,�?v�4p;�[b 3�e>2݀��&˂�T"�˺�I�EЫѲ�W�:؂����%Uڇ��N+�%�J�*R��XO����^����GM�~j���Ҥ*��$߲�/�`�����`}��a�oج�ҟ���|��0�Sbbu�� ī�:h�-�l\}7-Q�&�[�(?�.� ���ti�̳��"��t����`"O��4�B�P�7[E}5|$r�;�&�t='��f��9�PWp
�(���+�|q�qC�����:n�r�7��<��p��M�o5�"�s�>{$��q ��"����ݘ���S��"�W���J�$�r�A~s*b6$sT��3%9D��Y�F�Ņ�U�E��:���	���J��kHu\5��(����M��5<�.�^SK`����X�}���ԣI}�и��Ѿ�*Ȩ�K���p���T^u�z�7�7�w���:f�G�5^�es.Œ�p�-�����j{+�r�?�_��ڻ{�|}�
�#�u�8V�k����ţ��#0�di�;�A�e�d%X�ʩY2� �s���<`Q� ����6;|�B��f����DJ����lng�<�Q3֌�N���c���	�?J �i,�]>�/Csg������P㚼����>�����v����F
jFl����k~F~�7���BA�0Q���0�K�:�L/U�3�׺��]�&���SD���$��MЭ���H�~)�wq3������J���-����7۬<)iA.oT�<X*aܻ5��iңZ�M��#��m�F�u9'�=�!O��&�zZK�;����c*��J%��0O7�����\�J�@��x�L��3��;��܆�ݤuگ�	{
�)�	ZV
��E)/g��i��ο��_��cN�����5�eQf����c@fɓ��lޢ^ͦ!
J[�Nh�"E��鰙� nm㘖��Lg�����L6����ݤƑ�"���-䁝yϹk*���������yY.��{iG�M�[�3�{�����"00S��:MU8,���A+>D��P�'�z��=!���P�N��p����>~0�x�q�K/2򗽙�6�����>7�gJ陉be�Շ�}�H�-9�2��1-E�g�w�8����N��~���)|�s�Z��Aܧ�S��s6��u�
RN@�9Z�:�qZ�;�;>Ǿ��3�孞M�w��2�x&!XE4yQ(���;tR�
v�T����K�����t��5cZt���
�A|���2�*22of�=�O�1������)"���A�>���	�n>̷G�um@E�}�>#�8��?%���P-ӣFS���r���<E����o���N;��ku>¤���Ugg2�8u{�Ԧy���?�w�G+!y�;{����˄�͆,X0����<���{�,����@B�c�Vv&|�-�|�������h^W�0���z2`�� ��f���n
UDD{�F]��[��w4��Aa�bA��;�Vq��D~�
�u�?��:d;�G�������-%-aPն3C����=5��W LC���P�?��}H��-��t	BV;��vw6¤i{e��}>�%,mc,������:dQ��xSw=FmO�V�ǘ֖���1~f��H��ܣ�v�hh��.�ex�Y����7ט�O�`�s�(,v�oCp\�Zn�_�ζ��a-���-�٘���N��&��:ZR���CiE"�$hq��QE<E|�@�]��Q8�ӎa��S�h�u\��3f��ya�rGN]����Vs�I�؁�|���"嘐.��W�K�l�����"����ş_�=����ٲ��bv<o@ây"���N�R�P�n��d- |b*:"�����eg��gۤ�����횒� �������S`�ܒ:���C7`"�s���Խ��KԷ7��a�����#�; �<���Ύ��ݹ�����-j�Xɭ�J:LȻ1!t��d�8r���Ͷ������ːU��YG���S2r#=(��G}k�I���!�p܍�0C��Qe�ti�T[�W���%AQ��Ш�Z�������h��G�f�����m�`�w`W��6�]��\���IL��8b�M��C����s�.��+�L�w���g��@���[�r�t霣Y��v�(D�r�����)WS��NW�љ@��R5z��'�> �.:U}�-�H��~&��%#XcĠY/L�!DeD��iM�!v�	�-ތ��@A;��3썟�>�X���3�kv��l�cN&��D&qaPn".E,�B#�>�r*��\�C����� M��"�͊�e/��Gr�rԕ�kB�/��>�-ߝ�,ft����K�9�M0�j$����1?�N�� ���:�d��M�@���x"s�e�䴝�.~i�\��4�7ͽ���h8��f&�^j��`�9ْUi��m�t��04D���u""���:�z/tâ�W]��Ps��\�%ȷX,��Bh�ʭfw�f�>X������`��8�дF�&Hg�l��d�'
]Q�$`,��
*�#�D��s�	n��餲N���R��:e��O|�<�����G?k�8T�+ ��ܩȼ�
�Hh�p���o�`ɉ���M�1�)�P�ox&�G� �m��(+"��?���~�%{�;��1�%��Or9@}���J�;��,�Vr=Z��t4�i��Z�Ѓj{��1)�.������n�%j�_2���
���L�P͙�����ٍ��� ��	e�|g��x����@6�)F��j����y�O#���U��Mc^����Q�;���ۊR�/��'%�{w-6�Z�d�Dr�q���V;>��HR���m�A���e��W&��� ��!���5QZ9亞���<)Dhw��}Y^�v	����,^�ڙغ4�mѵ�S��� ��^�)}p�*�z,dД]`�e�i�[�;�O��c@"�0�E��D�3�xg:��y�l<���BT��˥a^�Ɵۇ�]<޲�1��e��Ğy��ۈ��}=-�"+nz'K��s��/.P��[	�j9:;*�ҙ|�i�v8�@֓L�z��Kl�-��GW�5(���9�ִ����ш��y�8I!�q��� b�&�4�6�"�:t�`}��K��h����ݳ#c����YP"c~:����1��O�ma3U3�6gSӆ�=]�k���6H����m� aI���E�A��>��8����8[E=a\����#&��e��'�'�\*w��,Ə��a=w-�.-ޏ��}����K���~���#0Lܪ������J����5�I2sK$z��;^G��|S�>dB�.\ʫB+J;9I%��4���8��o���'}�M���������eS�鴆5���q5�Z3�Q��ƓXM=��am����Yva�����WH�t_��4�JݼYWT6��JI�*�[���[t[�����w�:��2U�_�$�Ϧ��lP䚑� E���E�2�uL<�Y�~E��>{���]m<7;�/!���	�2�V�����G59����@���?bXW�ԐZ= xBh�"/�'�I�:������U%�<Z�ヅ�.�i�/��X���ߎ���
3�� �e�bsm$8������
v�I��}�>�v��srT�ha��9w������KmH<i;��cx��6X�+�Y.O@�6|&��:�s���-�:`A%��q[�r��4�)�@��2+%x���	R�ab��5:_ǉ85��WR�Ł���3`G8��
�[��8��͋�M�"� �1�BBհ�����4T.��x��;s_�Ru�A>Obgy�JZy�P-F���A�I�mK���[�Rc�[L����Բ�����֧��`��v��c��V��=�v3���D��s5�	��^|,�X�.�
�"��ݪ��\5���
�	/�:��^l̲g2��TV>N�_�+�OQ�p���^ac-%kt_��y7�+C��	�\���gX��0̓|��W�%<:>���2�7J)f\�c)�� L $Z��z�i��_5h`#�m�0�����8i��k ����}��(��t�����by�	�W���nd_h��E\0�$"gM��KVZ]~�dP�/1�5��U-,і�ɥs��oo	�
�E%4�5E��5��=���/f���lـ�LA������K,,06�2�n�Kp䏭��;�Y�.~$��z,��	��ߚK�b���EO����4|��Z����'
XpPS�F�<!�Z�k�'�)��"� ɖ=�����H��C�醜~�m�F ���3]�
�|/����7�����&��M_�e�<'(�m�>h>��A�R(e�_|����OV\8�G� ��+hUߌI�e.wD��D��O�7��w����!�������sVzv�������޾� \|t7k��1�f.W{{v�xk�e�Z���BQ��|D��^�!R5"�T���#�]�~�kG�{wƠ�jGd����ik�p@�=E�l,l��و��9�IH��}�t��l%��� �Ó�QXڠ����7�C��w)�q:,�R�'�T��%wi}MLJ�'���"(/s�"��qA��jے*���_�DA���qOY��IO�J��ǥ�=����U=,�F� A�^��uJ���R�h�4{&���~��C��AB(;:D���\̄����1�j�7�.�@]r��j^�x2�߹`��e�۴Z'��A�D[�p�k9�Af���d����b
G�ӎ7��>��a{��C�n���:&;S���r�<�����G���?�/LmP��* �L��>v{�Ϋg�Q��8�����Jp����|��f.9Ƭ a>y�g�Z��0�09��`Q�x?���a��8���S�mt}�t�]��.d]^@ЊZF��؏'m�t�
}�YHmx�Qr(x�����9uO[�qͯ�;V�AW�kltk�'�G����d7��xp��lM2'������$	"�� ��
ntru_7&*���&� ��3,%)��nl|���;���>��B�)�.@i]�Wdw�� ~��R	uw����y$�/�+�`��!�}29�s�׮�r�H�4.�����ٰI�N�{Djz;�lel�'-�������ʽ���$R $dLƿ� �6 ���%���b��,M�}=wX�����1 ��u�y���H ��E����0��J�;֯O��]� X�{-��)�"�ץ��H'���3Bt
z��}��~� ���=Őݷ���.w��rk�� ���M��A�*U1qN�,G6�8�Os����d��,s9�|���!��κD2�8�� ���[suԒY����H)��:�6���?�	�����r���/�`&���k�g�8�|��vt*/�E!Ń	t���x-����l�^9\�IK^'y41�/a�Fd�.����W��C���[�c��U����60&�����n��̢"9���`At�eJ�[^�wV6:��w�����rJ]��<���ˣ���Sh�b޺֌���o 4�s�3&��Ō��=�X�T����؇�5��+R���]�t�LPpEvn��õ���?�eF 5W��C�ϘP6���`�c%���̄svgRPԀ���&՚��En�3�!},v�ij�E�61�Xe�)�7I�1��-'8� �}A���p5bc��$�d[�j$���xc��/_�d�ܣ�7۫ۜ�jbdA���e����Y��Z�dN	w�6�(R�vݚ|�Լ'� ��yr#��p��q�� 
6�4a���\�kb�����Dd��(R�U��yl���P<��U�1�0��«M�۠�SŅn��-���g^�(���
���1h� �p�Q�ʰ�A���%@B_؆�w����8�OOE퉫��D��Z��jG|.���E������.�:�p���3�{�R�D��h6F �ĺ���)�A%�͍��^�9F8c����_g�r7Xw 4�r��)#�n����IE݆O��1��]tϔμ$<�ˀ)�ρT��"����\k��C`f��%��/��~xG�j���\[�leo�i9�c��x�Je�5HS���+��I�y���D��Dj�GBx/�KC�����f��@J�/v�q�X�&�EW���LOIѣ̫����]|ɮ����U=��2L�V����m�^�1��nĈ:A����4�Y$5?ڮ�Ɖo���Q����]�vN\�t���X��	���s�ς&қg�%ѽl>[��G���a�֡�^�h��ݤ�CʔJh/u�@�����%�W���� ]����Ud������ˋ��g<�O��ZǴN�:�>�"�������\�J��H�V�f��G��j�_�bרY�~� �[��ܐ�g��X_�En�%\��W�ɖ��G�E�9��Gj}���î_[��V�	Ya�l�b^�}=B��.�7m��^��	L�S0Ԅa:�zc"I����R6 uGoL�q!��n��j�ہ5�?tκi�r̔[�������E��`�vdW�����<&p2y7��[�[
�����o� ���' ���xI���sI��sz=[a��Q�M&�U�?b��4�P��Ǜ_i�g=Q���^�UpC�Fv��s�,P2�2]�*�4mg�z��sܞ����Yh��B2v�򏗷���1[=Ķ
�$�ObĆ���/2Y8L����`:�����삥������sg>��e{$�]��0F�̎��])�*�aOp�U����+t��-�ꄛ�n�7��P�����U	$Cy�˖S��+S�p�S��[�$�||�t��9��/��'-�%l����x�5>�2��Q��H�`K1�H��5��5��k1�X�	w�B`��J�����`#��#�͙)���ʏD�{-\\�iq�=u�R�ye�.��3M���xm��l�U�T��,���@ag��7>�"ūK�i:��PÍ�A=ؾx�p�R%��>C�j'_Z1<+D��lĽ~�tjD)*�Y�F��A���=�����u�C3�����t��]�?�J�~��N���/�|�N]��c{�D!6wK[we������ק:G�;�đL��.���ԋI�`zq�qO=�j�����	p"y3rx¶�{��ы�?���DTQ�����*�w8��^a�����;��*j��O`���E�P��SQYY��A���14���?\�i�j##��EΆ�\G���S�.GYv��E%o�&��!��y˶�{�jP8Q_��u�_�ƻ�#�CjٶV�7(i�FW~�X��8�����\9���}$��E�B�)��Bt(M�3��P�.0�B��������ӥK�M
m:{�c�'�8�Y�DI,rf��4��&�b�7z�uJ4���շ�pd��Ǔ�~6g7l5'S�,5&����t\K���qw�sj��V�|-�� 
�O�v�$ݶ;K`6���o��x9�R����p�I��@睪Ĝ'�%�-o�/#e�gf~��Πk����(�����'�y^�0L��w	�M	�p�*5���ŞX�Dc �/ȣ�>�9$v�8`t�6!�g8�����`���[�c��n�g�ȩ�r�-�I��Vդ(ہ��w�-�^�v���[rGm���c�	�Ob�!���+�x~5�׹޶Z������O7��� =�k�Z]Ŋ����׻���B�'��58�;�[� w�B9I� X�2)�l���8�ߏ�XjA��:�y̧����Q�^�ּ�%3�*\^���/6W��p����>B12��z�9�J��H��x��{A�ݕ��Ci�C��pn�����:�ۡԬC;�˩a��B���j�E&�P��(�qdXZ@�+��;r���
PZ�.�q��Ŕ9J�cY�	�Y��.���b�
�)N���Q)
I��_�ƞ5h�U)l`h͋N�s:_c5����Z�|e�;L%0H3���]�vg��$�[��bE(I��B�tX�{0g���G^�Dt�1i	�OKȁž �yf��@�L�#�Y��\��He�Ak��>_ө�7I� �൳�L(�H�ǥ�)V>������b*<���i���&�JC��b�k����ׄ��ȕױ�wO�K�2�Ireo �g�9�SN*���M�wZ�~I���52�4Lk1�
@Ac:����󆺝�`^�qel��Љ��lо$���:�b(}����{Ee�����Wx�řӳ��R$#�9i��+��^1v惡"�Nk�󐩌��>>2����3k�v��%�Nˤ��U���+?-a>?�7~~+�"I:W-ύ"�­Ԙ[Q��,ռ4�ق?�H�9QX@w��a*�&���P�rb��ˆ��ܙ�ҋ4��e�Ϭ���z2~^�aq>��^sz�J^��tP^�4 G�/
"ޡ�۫���nF��i?�=�rP���op3�VQ�_���7�/0�����p廄.����R"��kYa��k�,�c�������y���ֵ��E��6����fHt����:� (Np�)Q�0$Iw����sZ��L�<��W��,��Et~�A��EW�V����o�*�~N�=�`���6���GHR��P��Bν�M�>��>H�1�Q�w�.�����P�kX� ��� m�:����x�?��~PЋǂ�޶��N�� � ���F��i��.���PF��*"�cDQ��`�%d���:����4�^��]}�}I��E��y�,؉��b��Y�Y_�ɺHx�ѱ�$b����;�MΛ���2�7{6�<����L�������I�%�1 0��t���7�y��/����C<�MY�eN�{U����(�P�f*���6
��1��!�>ʓ�Qt�D�4�8�I-�ZS��o�eM*�N���\A�ԑ�{�@�U���/0���/�T͟×*xנc��/GۣY'���>$Pw[ 5�0q���[$��_��?{�+���oi������nAGS:t$�%�E�5\����g���!����d �������'�n��PS��CG}�F凌E(�z �;�������O<	�����&�+�:�#���6$R�HUq�m��E����%z7Vq���d�=�L|sn���1O���L���i����4��SG�ȕ���5�g&�0 ���s���w�}krPՑі�{"p��Du?�x�6�����]���þa�"� j�����^��A��c�"�s#5�O�.�*���N��v|��_z)z���}{k����:X�H�5>�)���U	�m~������}Q�|�c��U^�p�
��	�"k�&���غ�!E�Z���\�2(����v���w�EU<�j��=A��	�[e�_�p�)J�ߟ$\���zO:�",<�nZy���$�v�'��f�`�W+�q���Ҩ�@v��g3�;(��L�p�!����.��Q����0�ĭ�yٗ�ߗ��}�m��ꈋ�U�I�^�}Q֔PWB�������٣�u�Ft�<UY?�T���@���m������.�i�~����R�j���nt��(���ua\�^�լ8O�S&'��O�OR�2��=�0a��Dzh��M��6�Q��#�6����+�~j��̯A0�J���K�?�l?A�� ��z�FH���;��8%V���\�*������O|+&��c9�<궊�{�|�� �D��.�8�mN*}�cVV�����1Pc4p���U�}�J)b�
nkU�ڷ�)����ި[���v�o]���S���Fx�1(��`Q���R2���H�ˤ����E��}���ĬdA�1���e��#�i}2�(h����v�`+U�4,�v9řӷ��.����3����ُ}+�+O�YD�6�{�&�e�k1�w���Hz�eЇ�^�N݈��yBL�<��,7�>�,X�<q��4���
���D�v
�U��#6O��`���uE�����Af�$�`�?`�6,�Q���M�]�T^���t4�N�z�AY.޽!/R!UmZ�PMS����L�.+��yPJ�K��̡1~J�t�4_�casK9�Ue�ܻ�u��mS��ڠ�)C���!p�J��Z����L�Ovc� "��ѓH���Z�����J����ʇp�䰶P)�zo�X����%�k���j ��;d���_�v�f�(/�������� ��_���/P�g,���?��O�w�X6�%���:�w��%�c�|�=�c�v�ě�ڰO?n:��%�=#�h��o�u3Cn��ϛg �QP4Dmc8�*�'�P�䉨r�O%���w�듧��;�J�Z]Ϗ��wSs���P��>:nJ�2�����0�h��~�0w-9!�a
W�sZ��/e���C{}W}�{��r����Us�9D��n��:>]=�X6�G"�ug�m�)�U�6��ׄb<����$+Kk��1�q'�!�'���N��N�>�kℬ)�!(S$\�Z�(
�����p)���4r0���	m0#l284�g���x��ٸO��m�.�;�b��<q�Cg/�w��6�5s.~Z�zv(tM��m�z c<>�ܿ/�\�2_�㣽�ͨLv<|n����L�	}Ǎ�0�L������1լ��\"1�Op�Z	�lJ���K��!���b���A�x|�ړ�������Q��q��ZȤSZ4]�0J{;L��s�+��ytNnpm�)�Q7�9�� 7�d3��e��%BB9�6�3���\A�fJwti�<&\�aG,�W��1��iSn����W�q��������ʰ��t��W��9�@mc��6W�e^��T�S�|���Ul<�$��<]4r�:<9ec���O��o��I"ۯa���ʣ��t��K���'6n���׷{I��b�yӽ�Yc�XX��`�2Ԅo�d<�=@�גm/�50����KQ�s�l�w���~i�}
��m˳@P�W\i�l��$T�s��*�A�lu�?0v
���D�k�hv�-��h�߀���'��M�������M�������/wK3J�tc����6��;$.Y�#ee�`�.��Wiq>-��D�7�T��V����N��2�(H;�J��ć��O��K'��V X�ƚ7�����(�����׷����$�����s/�zq�h�6l�{�w�}f�$i�T�B���ւ����[�i����,K�O_A�ػ��%y_�6OȢ����Axa�.��'ؾ���+���7[	Ј��IY�'�K#cr�n�d4kp�!�l�i$���v��_�y6��V�p3�8 .����~��'(�}�D�H�%����C�h�Y:Q]y_�`�,T��K�
�n{�rt��P)����r��p�xъ���cv��{>�*�Ǯ�����]<K�G��]P�E�(���E�-L@�|
���'�EWQy���V�����
�LՄܓ��r�t�ʖ��V�Ӻ���4-�}��9��醧��	L�\�IK܌�X�$ 5{�s:z�j���d�jn|�[I��0�#����;��b���@S�����y�o���h�Ry5��Ȟo	󷭎��a��_ɡ�؛rw��m�X���x;��������{�x�d�v}��r �ryV?%ff�lq�%Gar� ��E�s�v�;�O��[�1�� ��	Zx~�);�@)��D�6g[Q0n�#U��L!B����!�_;��		�?%�����8!�|Vd�����T^3����e�y��2�J�FMY$�P=��o�;Fm��h}{u�;CyT�(4�.{d�η^a��P�����=ֿhpnW-?ް}P:�C1o���l��O;���]��K�k#}Յ�"��&a�6�KN�pS��_�o���2�n�R�Q�a$ ��%��(���-�C,M��2�vS��
����7ЌG�T�j��C���ma7A\�.��(67�ܦo����X?T��ŉ� {���#���@�r���5+Ѻ|� d�d���
���t33��d{��Ll3H�ޘfI��$Ȯie�|Y�@ݱ�;Z��������b"��9���yŠ8����#��vvg)��X��Т?�;`ӎ )!S,�ҋRq~`}P1�ʡRBT�C�l�/�0�niB���t3�装�����Z�+!&-�z�v�
��1R�{r	Xx��[�R��K>0���E��k��.e��.��^�����
�U�uhX)�7��8�JH^ّ_μ&i��u�Nf����{�@4��A��I�=[2$�{��t��� -�D8�6}l��wv�	_~-��.��D���\]J؞4i1K	�����s�8ov����a��|�u��ǋ�a�"��q��^F!�S2>�'�Sר.5�l��] �*=y�DI;V�:�>r)���uN��t����J�|]lM��f�&�' ~L��}j��([�m�����`��y	b�e0B�*�6IL�ۭH�V�����R��5��5N@��I���S
"���s�� c����20� .
i��9גnK=]��*���+}�z��^/���${�\�t1�8��f�.�W�V�?�L�Ã����Q����}�N/ptP�|]�/��!��*��D���")����ӱG0Z�k�k{Z��d�՞!��p9��w#��A�z����3��aM\Z��ʕK4ƄAԠ�U$6��v>f�5!�\�ճ��I� d`T�L��>b��G<W,��bD.�5)��p��ƻ��=��Q�#��]�c�-EՖ|61Sg 04����B����gT�&�q"���]41�C���r���7�(�g���׻�#��v�(z9��R+Bem��o���j���s��g�{P�7���<B�]�~1&���9Y&�������к�]���1~0�)Q����VN�%4�LLǟ�����m�e	�DyЕɳ� �`eFaϒ�R/����E9�_���n}N�n�"r��ʆ���S
K3���ۣ�X6Nk��f�����Y�x�~����kKOr;�]Q;KF�m�fk�Ç���\�3�cg ���Y��#�5u>�m+|7ԚD%�0�y�i�fĩy�53ؠ(�?� �Ȥ���<���(9W�,�w�C��=bs5�̈�U������J�Dt����=i�Ԡ�E�&��T��M{�F�0�����[w��=Y#kT1g2�,s-���O��s�!�W8Z��F�L"{^�y���<�:�a�����^`ՠ��e���sΉ�_tgO!�.	�t�@�;=H��GWJ( ����=�e�T!�us���L7�a�E-�y�����i�'�D�D<t�/�Z�b�1�~{��Y��bD6�`!�|��U�0c�Q����5�W�aH����,���3䕐hwN졶����G*D?(�b\�;7F����~*���%h���Z��ڦ�V��g�l��"6��f�&#�kV�=���0P��+�V�@��FȰ?>|.��l��(���L��/�6�g��P^����k��.P�� +س�$X�z��1�<5췋b�38D�W�ܘ� A ��.���>����x���Ѻ�~!p�����i)(�C��5��u'
 ��^u�=3'�ٌ��e�x�$x��>��:4����u
A$r]�WBN���É�h�lK�C�2Bx��>b�H�;>'�ӕ:z
<�NU�������J�<��ʺv���	$����X@P���ߦ�G*s��B�܉��G��Q�)*��J�|�N$�;�88&w��>3�KI{Xy�q�u�6���Dќ�Ld�Oc��޻&���W��>_��XB��A�2KA�[��yz7���� C�b�2�����Q�n��t@h�+���,Vs��fRd��BZn�=�ތ֥�v�u��9,�ȗVQt�Wa��ݬ�䚊�+�"��ٚV�';ѿ�w��>��&�$�=��
��B�7����E��hx����%t�+0�%��?:_�@�$�B�����p�#���p:�Xꊽ��ѷ�縚PK����#2��x�fc��������j�zM��� ˤ#�k�.�9@M����W}K��eP��ϵ��CTT9��~.
`g9��e�4]��	!�jqGs���u(֤T�;�ϭ�����%Ya�����!G�,q�3�t�C�N��q����/�p���89cP��X��XS�JɁ���*�K6����q.��b�醩H\���fz���T+_�y5�b�����F��h�M����G��%^�Λ�t��W�$�W8�(i�!q�&fr��|�9h����U�y�jϹR�Z+��Gζ� �י���? ��������i_�+��JϹkr6�3�v��5�@\�=�����C�2�$T��.#�z-ձ	��v���d�qS�堹�ķ6�%��E�N�ܒ�cN؏&<�wU��[+w�ܳ@ T���������Ԁx��
T9��V������?�c�� ��6 Y��Byi�pA~f^��@O��F�/���]�1m����IW'��wĴ֛ۮ���
g���5��1��>a��=�����~3([ȓ�����p�B���mk�P����0�^P��H��%�,΂�#���c�W���~E��������L�&�ٓ))b5u�7�J�O��d�BA���Hd#ɲ)�
0��ԟk�����(ʨ#}���*�rԯ×0{f�>�~]C�6��
M��ؼ�$��g��N�R����}Q�'��j���q9�*n����S493�����+�(Ȝ�Q���\	�C;��	tuq
��ab�5D��2#)�/_2��Qs�	E��H����8�.vs��&��AvQ�u�Ok#K�If`^�U٠&�@_#E�)i��o����O�`7jp�q�����"��v��!�2 *# kQ@7��$��(�����5�53  ������%�$;F�"�Y璭eCl1�ˀv$@����OT�	i�°9�P�=����OBƯAw�����֜ϫ��T|�f��@�њe�����9�F<!<X֬���?���V(��������j��vr�^�,�,g�S< ��..���X��>��[�Y�>ǧ`��KK�Rdh^�&��073moG\#��\$�=�M���p�¼�^��PTM��Ƹ����ڶ��:v�ۖ��]����5&��-�k�4L�2���b"�d�-6r��f���`-M����2���n�#qp%Ӗ������~o��=xf��wS��Ls�5ꗧi�)'���0�&��<��;�`c��?��W@.�2Q�r�=)�b-�7I@����%�r�bN���ƨ�5�z3����da�Xb|'�"�XHXnL���' ���;J�߭N��giS�m�n�?�A���N���T|Ac�n<���"��eػ�{x�54f�
e���&�ˬC�пmC5�c�Ib�g�9R�pvn��[�&�,��SM�U`KȢ2dQ�!۝U��6ci���p���iԀw���+�Ђ�+� mq�~� m�7�ر>�FJt���W&���c�=[͈6�Z�5:vJ���i���;;54,$�o<���x9l���`M����2\��H%@��޳�гl�#�>K4�G��;9�pl�x�ϐ��r��x9�-@����.B4�,����d�a�:v��Dݏz�<N\���<*� \�ɧ��	(�|���Ȥ�>�����ՠ�q_���n�(4��l�4�u�����
�qqy��9/�s��f�����^���cîV�$�F�d���ݐ���E��J����_.���E�-���{��#b�LH��Ͱ��)�d��@�(����8uɬ}
��=*Q����ݒ�_���ŻL��;�Rr���-݀�=r^=����/�B^�9�2�����ڣK%t���Y[��pRu�"�܁�'��%���'b}�Re�v�����6}�����7���TnVGn��n�Z?k��3��|�J�eJ�� s�~�7Q�wc���C�C���W���&I��s�=�Dzt�H�8�2�<����.j���}�@bXfd;X�v���[�s����Җ#�\qd�$M�`2�aNJ��|�$���WGP�;��"����� ������yLA��J�hܣ���U6oF�Й8'�+֚���V"{�D �$l�A��J�Gdv�j�?3؆_���
p��E�"ܥ6��SMS���?��.A(���M���2t7��:�$�^5�F4>��-�Y����ю>�����c>�J}�;��݀yL�!�������ƞ{�,� ��g0����_4�DH�`���gZK�Ɩ���)�&uY��O���l�C��n�BU�����*$���tJ��.D+�?��Jk�Q�@}м�|x�f���n�K��⃻�1��v7�����6R�(qP	���*U@y4T"��Ą�i�ڳFy�1l�N���?>�ƒ�;�R�ߩWq)��nBk��`� o��\���4₭.6-�)%��B@E�/V'��!�=�����N��Ffi����x�}��AJ��h�h#��B����Τa��o����Z�c\��k?��q�<_I�����r�m��.��w;�����B��a<@ʏ��7���I�!���+�d=թ��鐘����v �����@��W��~k�n�(�`e3\�yo2A$0ܕ/���������Cb�'tG+�ۿw��I���ޓ� P�"�p��A)�3�Q�_>>
t�ij��8q��P$��Z}6&Aq�m������=YBzgXY�2C�q#��R��#����Ѩj���-��+6n��&�=�wv��ƍ��6{������?�8����G�Mب%��J��6�&�+��i�~��ȩ{�厕�Iѣ���o�W�2���@����_CA߬pS7L�|N��3N��Qb�g;� ivR=5I.&�� B�����[�:�a�8z����\�.���!�|lO)���yN��=�x��B	�=iC(�}_�� ,�G.�����Z�v�>�Q��꿣�ܶ�/O�;�g��LL�$̇�'�?����|��p��铝y�J.�6�H� �����]��F=;K��|��K!��k�a�������~P>��H���~�k�#��˺�|1�]����刞�>����&ȶy�[�hO�ɪ�~z)�x?�d�%Y+�:��ؽ���}�pYtH������ϟc���%n�����Fb�C�[ԑ���pe �c����a��c��C�^yC(��'"|�kH������A��ML_��'W�+�y��֘򔵶��vG�è�j�<⚍P�)����\�n 4�z���0����R6�"��4�Α(�{�X�����z�(�P5�Э���/dP���&�RI�8AF/�sےA��Q`t�܎?3���N+�^4�?kj�6�bN@@�N��AB��z����.S���g�R1{Q'�%2�)� 
i0cĵ�i����%v��*�h�H�%c���$<��;?��#;U�Z��D���~�u�MtQ�
�Em&p���GW�OV���s��4��ǵV����_"; �H�e3G(�P�a�WNE���)q�DbUT�V��~��SH�N�$鋗�g?a&�2��""�v
����~_��C���=�?� �����O
��2�r���g�y��B�F��r�� J��E�Q�R86e���̪�bZU*�S��)'�%#��u|Ѐ��^.v_�+7�ۍ�p..�9������־�)����'���f�X�R�U�R3n
 ~[��}��DF}������=��ձ�Q�G�M6�a��$^'M!N�>¬G��Ɍm����T�5�z�<[��"V� ��=ţ��`"=.jYf�䭞�kں_��7�z�a��3�ɝ�jW-K�� ~���J��әݷ�8bc[g����nS�є���(v�V]����Mϭ:I����C+�}�pO&B�8I�9oU�ᄲ�)����yM�E��S�.�EBz:�����������]M^u>��p��I�D�+|[���>%�Ɯ�2́�/�ڔ(���lX�i;
J�U�	��f��t)9RC�V��LWM}bTC�UY-�lfd�\���<t
;9u�gD��zP�^UF=�Su���Zw�Ex�:�hJ�Ҝ�S�J��~�c��~b.*N�A�R����w�SW�����B�l��y�W��9�N�Gي�jM@�**�/5�9��;��k�LLUܓ�)�:���ݖ�\]�g+�E�Pvd0���Ͻ�vj��+Q�(�z/�т�o���G���ˬ��'�ڏB���KQ��@6�En����f�Zm�h�Vi b��6�$�`� �&�#�偆7�]�w4�6��7��o��<��!����?�nv�e?2�x%�;�n
�7�����XQ=;kcd2g�\���y��;!�'�!4��1�UPU��д��V�� ੁ[�cW�k�bz#�:#�s�����SEmx	%���c���t��(�F"����r w16�!"l���%D�1��Ee(�
�ZQ�!���fR�Bn������Ť,1*c77�4/�W��4=>eޏ"�R�����9zC\D!͊�Յ�P!�ģ��w9�:E��g��=RP�1�&��R��L]Jhֻ^��5�*0I�~r�N9¼5�9Dx'w]�^��Js��"�L��Zz�y$6�
|�މ�y�E�c�����_����U�"klU���vL���������;F�CU��/�gpEt1l�x�?v���i\��"<�3�^�̧%��Xa%p/���7�EQ��7�kr������#^Q��8d��w)���6�ȡz��^qsڍS�g֐BS9�G֙�.�C{���&f�6B�)E��[
�)�[�*ޔG[l�)8������I��<4���z�C���s�Νs��`Q_��
��?����쇊.dy�S	��?Y+>,�nV�f͛˟�@�_�e�R�� �	�����SY��u���.E����L9+��B��2�>E���m:��"�W�\@�0�lF����C�=O֏���9g��ѷrUP����ō��A�94l��}R�]������:��?�႖*������{�WГ��� ���=��t��Z1���R���ƥ�^�ڝ�7E���5���&6��bM�*J�[�\�,�Yڍ�<�H,�n�[�V�!#�\7˯�i�e��ְ��j)f��ޔ�p�82*o��PZ��p��{ e�eJ6����ͻ~p5��W�0�S�dP��[V`�ס��TAC����>��/�	!���y��ǰ�(SWTm�4{!?L��ɚ�J��]>e�>9���:y�qps�u�T\��;��S�e��"�-�_i�r��� ��UMj���=p3zɇhă]�����#-�TK;�a�h����Y����Pf�%�z�^'�l�ÝW���U�q[� g��&HȬ�7�e��{M҂?�Kk���X��y��)����5�X�|�����.����=}9V��z��F��:H=-�M�))�ކ�V�z�V��Fr\7ۡ� H�OM8�����!$���_�g���.j�\
K��tX���V�J_��j7��g��tl
���/�����:�=�U7�a���{���>��-�@M�l7C�䙞� G&a-��~�j��د��!Y��W@^sL��Ƃc�6�ڣ���5��/�l,NO���?���K�a^}3̫s�i
p<ܙaǽ�Vw3J�d�K"�B�
О)�՘��;M��si=�q�&��BL�e�H�f�������(l�ap� H�b�t1�.]������`gE_2��;���)��7���3���\e*&�E1(^�#Ns���*�� ���(NT��3�%?�m=�(��f���kӼq�W��8)�'t.�ˮz����<����׋��Mg���L���U���f8�Xն��K�W�x��ƌl��N�s�|̓%�z�څ�� /�&��� �����R��ٯM�C��r�<p�k��W��+7��� ��8�%0>,�>>K�8-���R=)"S���̆�D��]�[}�th���2ݞ������#M�� ��g�r��u��0�)��PHH�=�}*IL�_H&;��j��o�4]3]Ѣ��Y�0�a+$�r�s/������%�;�#����Р|��/ݤ{��-�ú���{{6`c�_Dχ�޼�߉?'��9�������zCk4�Q!V�d��/�A��>?��&�"ݟP�q���y	5X�q�B�?Fṟ�bT9K�^��k�r�sZ�u���|�$���戗5Kd�$#3j��ٓ�\J�,;�b�����K�D�%Ž�.�9lU*�8?�[�3�������B�%MKa�p�W�6"^���
��[��6�d��H$�[#��[�%J����kRЉݤ�yp�x�RM�~���0:�5�>7�SГ�e��E��bRiӮ�x� �o��KLh�_�~G�^�kஓ)h�����nar����x|@M�M3��~+x|p�����l��1�V�RܪLa�\1�5)'!����~tژ���D�b�3����R��j� )��B�0�B+/���I��/��D�d��b�Ѩa���(2�Լ��Wl��չ��p��Iw�c��Sz\�M�k-�~��Ye�D�e�k:���)7+6[ڗ���{�c6�6���R��<��9I���!އ��v�䄘u>�3�EH��d>���H�yy�ԋ�ԭyH���PJw�n�d>�u_!-�=�h�ǩ�ϗ-0�xA͊YmqR��2� [h���҆���C�Z���:�1�ר#!�m�/��I���˻8����	m��ţ�+�C"_l�U$�QZ]-F6�^�(j��qޕ�T�N)�PH�_��$�����'�>��f�1
�_����'�8��W_+���/���R��<y��C�R�u���6`[�v�D_�g} ��u1�j�ъ~��01y�B̖�&�;^f�.Z�<��G� ��[����7��5��,�����>���7��x_cM��[I��+4`���
l÷������S�a��ᯢ32�d�p3.���ؕO!���p�	π�k���X�j �t��)sݯ��2!M�#�M���$y��*<kø��HN�e4r�h5�NS���_*H��|T����/BF��1:�ɰ�u�WJ�uO�,7M�y�=
����&c��Mp6X�;l�AY�	�B��r��|����m�D`��Kf�T��Ob��O�C��?�~����s,Y�/�F?>b�����h	�kb��*Q������j�+GV_M�O� O�C�j�f�����	t,���LE2'SKԌ�9o��-�}Ior|
�$H%� 0�u.6�S�1�����U�f�Z�!� ��Kؔ���hꤦ����DAo�U�$	�����㳽%� `¿S1���j�>�����m\�:X����:DM$ј�3�.�������A�p����!�G�L��9���|�D7���8�8��=�B<+���7NCn��L�0�i����\X�؈�oK�/d൪�R&'�o�g\E�1���3�q5���;��� �����ˑ�a)r�r��J��S�^a��S�1�*�YjJ���20O'�K�08}���njB��@��Pw�;/��c�C>�lY��Jy)��\+��J?�$Ze��f{��Z�(�{��Ң;K���2?�=*l�sS?L�8�����M�2��p���F~NeC0!�$��F�}�$�6��.=w-��y.�C�en�~��c����S�O��v�ݸM(�^]� ��Y��Ȳ@۶G<���+&����;��w�F&��BYE��w��x�_�h[�U���#S���%��&w9U��DV���G$ｑ��~Q�E��&'Y��T�@��@�7I�Uˈ(4���g=R1����k ԏN�u�=�ᩴx�Vc�qa`��K��hw&��U���z�L��Z!J�� �̋mHN�mC�Ǘsc�&洺�f��7a�P�#�)o��=�ۧk�$q	 (�*�6:�U|�l�2[A��8�T�B^:پ)!�蒝s|��L�ƹU�7�b%��6�b���@����y�,�R���WH5�jI�!-���RL$`S�B�@.̶���t�tH5I�,񨺯����2��C��pa:�M�Jݳ�A���x���,+}�oS�+iQ�PGxZh�r�.d�%��n ״$4�̌Q�
�F5�����u����<Hl?J讀2��'�틊-&�zd��[��,��ҘQ>Ԏ~���Ly��p�Y�����38��;�L,2�1���2��O=�O-KU�U,_���ь_�^����C��5@�W�>�n�!�Ud�=	C�}<W�1��H�&�0��.U!���RLh��qw�a�}�5�G���)�8ڔ��M��e-���&E�6a�o�j^��<�$ �r�DQOcZ������Űe��KQ�A�Z]��Sz?Fn�~�	�gs+Y(��Xs9���v���Q/�Q��6�Uк�	��n�<��������c��KGD�.�������F�J����E}�5al�
E J�%�>b�ylǜ4E�z3��֔+��b����}�Y�'9���E= ��٤�>`/�Y�a"$���^I|�[9��UZx6\������=�yD�d���sD(�!Џ
1�m'C��&1��4~\�gYi�!��K����/�いm������5Q�%x�'�-��^Y[Ok>�^�@.k�f���ؽ�8�z�&�I�շ���ڝ�NY�^�n�E�� ���DQ�]Y���)\��x}'ݷc�\��Ņ0���������6�2:����4M(2@��.�lL�!�}G�3�RQ���Fי��@����S��,�|�	�^�p��"uN�ˋ���Z�(`�$�����>Nނ�]���	��B��D:�@֧ĥ?>u�dֈ���H��`�XXQ>&��e���xW��\D��.�����z�au��
��}?x:�j���!�?�e?Sֵ���]w�R��[���xa��o#���|��&�;�	GD2*��������2�V�R��7�p���:�g�ޡyc�\��H8��I9{����ă����J�MK�^{��N
���\Y�i�@h��4��J��uM�(6t�y/}z��흁�Ŵ���S.4�A��8����`<�Q�-�qD�z�O�jM,yC�!����LA�/� ��������(�J^����#�^7�i�E1���=�`�B��2ZJ�d/J>e�KJ�`�lz�r�cwe�`߈�u��.���� ��(�>��!q@.^8�d��kɆ�Ȩ��븰���-�o�����{K�9�8�+����M?L��b.�r��l��� �=�7@��ߤь�S����
*f�H����[g����(���c��\�lf���Й���:�jx�.�.�b0���Z?_G`04��w4��oJm���W8jH�G�������jק#��F�ӔV V��Z�3�7�A��ߩ��M{��fbQ���z}���>�ߵ��l���t�J���t�B����&S*<u�d���sd��4M[�S$7�۝���	-��<9*�j f��?���KW���K�b�F[3E���%kPIl5zd���2�|tW�W���L�^J��g)�����Q%YO�dd�b����~FX����DB5���|c`ץ��v��yP1�7ΐԱ��H��j��f}>;��>�#�Yek�S��6������+A�/k�S�"�ј��@��P�A�������!0	/}`�J,����1L���_Y��@
s�w`��w�r7j�C����d�w�nI	��E��k��9���/A]!N���b�	�%��\xMk�����́X;p�*�bf��>����9����b���3��&�ã�Ÿ���������e�'G����F�'�@Yh��7<Z$�;9�Ͳ�M��L�����e�Մ���Dҩ2�K>�S�pT��5u[�Ƅ`-�Uk����eA���B&{o�>a)ꂫ�6m��>������ʜ�a�l��$؍[qj�O��W�V����JlP��!pR�)JS�{��p�E�e�Si����uCFy�H���)w�%��m�����yYw���,��.��Ȗ�X37����6����?�{ñ�G�=�67g�e`e`�ǐ�K�C���ᬇ���9��Q�^�t)q玀��R����a�$���ݦe�׿���me����5U$..uL*���O�d��t�
�~	�{�����W��䘌��L��'�_�l�3���,_8�y�EG�Zy��⃤�_W����E��4&8;�־�<T�%�GC:���+ׯ�Y^p�/�ފ�0�*�S�L�[�@ ��򠱨���+���̇�pBb�7JY��A"�	��rZ��d� ��cv
�XrE����K�3�~�-2�I�lC�XU;#偪�Z����F?}w}��	.����p���#�!h�5������ 4��!XI{��#���x���T�3hH7
&$E"c�銱�b�§��|.U�����
ؕ*��Q��S��8e��a^Y��5��s�|#�7:�Da�1�8�@|��uт�I��\
D��G7����Z�8ni@ywB�,���7��[,ATe"W�h�"����(,�Z��L�R8�'U��_�Z����z�8���x]�^�]%�
�|`��LW�9�faR-+�_�)�Gz��X��#�L�r�^}�-y�0���˨�˔�h��*UB��>�<ss��J�l�
�<7<����~��c�7��
�H��=E�7
�cq�V%Ę��ĖƋ?��8G.�-D��|�U�/oz��Wu{C-�:�����tJ�JQ��H�
�ˆ?{D	V�p�3��H5�!A|m���4��F;ژ�}�/���_ ��7:�'��cªjv��V
��\���=)�X"b'/�0��fr�X����9�q�y"�s�r�e��4�T���n�`�s'����%}���m���W,���!ɭ��0a��������o�زR�㳉�Hw����b���F)Z!�����Qk¿z�k�F�y=�_c���j��LƔg+O$�م9GF��0r��e%,�V���az��7����Y?���pi���MD����i5bm�[Mً�z+��gK��ΥU�O��s�$�)�!�)՗�Ag��C@�C:ui��얜_���؛2( ��+w�(Բ���׍�*RhX�ܱ���Ӿʤ�`�D��	����*���`�J��u�/���U��F��u�Ɋ��qQ#ps�%%f~`5�q��LO���=Xw!��ZJ;�V�+�h����{]�8�<*�&m��y)�;>�J���'Q|���3LL���j�֫����Pg�m�~�����jf}��G�B�@�>��#��Ϥ_����'��̨�8�%#+o�xTR��}�(��]��,�K-@1O�a�#��&V���Ow�ho���ڳQ�3@�v*�l�5[3p��B9��9++ߩ����}ӘVS*%��=�X�����ޓ/�5υ�o��	w̾�=����arg`���x��O�c��� |�bh�.Oi��c��plR"���2�	�zt��bN�}FϪ���,G����j��S���G능��\W��p�ﲼ���K���o�t��� /!̅�,��3�Vt��"KX+��Ʋ��pmb�K������˥y�5Rt�vк�^�tqB�L|=��qj��P�h��l-��'?ј.�k�,;ȹ��s_��]���㖟���g>��������]R��3��)mO����q:Y6
�e�����-�S#����SLΪ8,mSũU��}ЎK�O/����9���[�mG��m:��F
q$�tW�B/�:�)�{��(�qoh��!�����G�w���R� t|��%�(��ھ y���~ObG?Z��0���z�3dt�'��P&��s��0e�J�3�R���PQ��6����4%��@� �G,��%�7cR�5���3����F���q�!u��ul�Hz���F�fp,��{~L*CTt�[x��[%�����U3��upJ<������R#M���d��t5�"3`���*sN?����e!ݧ�n����`�	d+��)ǳ����\z�o��[�NTq. ���~�|0�<+Z@2�g��s��'����n`;	��<('�`�$�TU��a��ݨNUpk�j?β�G�.�3�)M{fz��М�qKȘ�/�w�Og�5�땼!����2���l~��&�-�ni��Q�����R�2���;�OQ8yz|����6�A��F&U
B/�~2qi 㳇���Ռ�Zo�Q2�}��^S6�'���":[m�gk�E�{_�Z�LG������� ���no��L����hK�E�4'�#�!+#3#D�̝x���<QC��ep)3�7��ʚ