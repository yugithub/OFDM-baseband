��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6>�M56�M�I�8T02IW���4�̈́ipճ'�����}�W��Ny-���^����� lT��h�#����gd�̗���ƪg���g�����J$��ݿ��gtr�v����r2�H�y
�5O�p7ʰ�xV��}���$n�"'����g�'\M4I"0f`�O�������x�rkN��`�4����%��&<���l����S?!�j�շ
���ܦ&j�M4�F��rF`�rȆ��E�'=��pˁkR�r�h����nX\�nQ�8<w#X�ѮZcb$�mЩt�,T0��⩂>�-A�l��+{�[�e�M#�&8&��ҽ�K &l�kM�����>�x��²#s+R�D8��F1��Es
U���&��-nhc3�C�[�*;�[\�ie�£$o�f�5��'��3Xd�MCx����l���2w1���р���6'j��p��#�p��	J&8;,0�Z�NOSO�1(��7&���_I' ��,�4t6M<ǁ��t�N���_%ԏ&.Y;��U�A��@9D�h����/G���z�"-��c�Z[�HB���!�5_�J$�%��&���B$Y�9�v�5��1@�fD��ڠ��H���x�H�X�N���.��&>Pxh�6���о8��>s���&S��5=Y'����j�v�6w���1����Uc
���d�ϟ�M�hm9���:�����6m�ٱX�X5G�� �x�oS`��d*��G��okV�	�3�o^�{ue�(�eI�W���0е����ø�ڝ|�/��8��m���)�[M�)�T�_��Q��U��rr���W��ú��[�کW;PKjz��m�OO����;�x��?ъK������C�`��H��ɛ�V�eڦ7��F۲����~	��ܪ����y��0���}��'�qh���7�q�0n�.\u�ۈ���zԀMKd^�pG����I�<�ù�D̴�_5��p-W��:��Xt�����glp�K;�` Nj� IXT�AZz�K��B�X�2���J�&#'Cn���Is�[*u��3��8r�z�����"��SUASg�K���ym֘�xSbo�!Ӷ¹Њ��܅b�,9�G ��9+\S�P*)��	���.~/��� �n]�@���P�SC倚�ۦ���a��"C��R�6���be�א>-�,+q��4�]|#��)��7v�ߧ� �W�Iqm�����T�M#��0yb��0�$�Ư�}Bk-��s��bwP:��A'�	.k�����Ϩ��%u=RHc�[f��sɟ`�:�Cd��Fb`�<����P3�;�%�bc������p��~����C�S.�a���8~���j�Eb����&�f�|��=���qƪ�&�<�J�����R���_�3t=x���`�t���:o�� �������rXW<�mɜ����#�H�l���u�1j�<Tf���¸�F�t~$��<TQ�F��.��C�Mx��!��F;/F�9ajP�J>n.�#�������HL�	m98�ǡ�Y�"���U���u8͠ni�K�#���y�q�5EX�T ����[���+��D�>�+}�ێ/'�M�9K�^8�$:PcU��?M���e]O�v���qI�9�|��͠B>� p�^oW�����y�\?ng[T�G�D�-9:8n��5���G�v��.��݇	��\�����{����B�>�'�q��$w#�ƆrePm�@�-�sl�$<��-�mւ��:�<���A�U=S��?�]r{̲TF���:z����Tt��=-D��/��G4J�NۯH�0����)�e'�������"
KJ=��t^'D���`	J�u���W�	#�f|#��D9?��*����M��`fA�Z�a�J��$]�$���S�à��t����8��X��Q�W�-�}���V�f�Xِ�>_�ͼ��v�����
hd3Z�D;�oQ�"t����L����ˌ)�U�CkK��x�����ΰ���^�zvQL;��y{>+L2 ��`RV���i�F�\b������4*G,�QS�������[���!3�o�����aR��X5c��@��6���]=Y����*B�a�}���8XK ���Y�0T�$T^�\�؄x�7��H�b̎3sR�Z�ɆwLV�'�_��^tج�b1�ca=z��g	���0#zȬ�dU��v̀�rI�P��Z�G@k��y$80��z�V;<~�
[[)�Y���g�ѯ�0�"�<Y�$��:���& �-G��$p&�L��k��=�Cи�/�L�i�|<4C���-v7�ڄ�?��\y�Wx��Ǖ6(XՋ0��kx,M��9֢\xI��~"��.^�ۉ�?tȔ{��ƌWQ�	֎27�\�������N�F�pvZ�+b��	a��bf� צz�v;2_��%E��֤�A���H#Sq��B�}$T�Xaw���O{� F': ������e@�[�	Ǖ�?��*�B�%�� Y_���0���9T$�w�k�㞷�LN�V7�p	�y�ih+��hp`HV�ڜ�J��7ֈJ3��1�L+;�zM"GzkI4_��[� Y��q }�r��U��
�����VC�hmi���b�P*��B�a
�m̾���5b��c��e��Vs�B����F��0�7{1p$�]�8d��~��ʝ�w �c�Sq�؎�em��M�����v-.u��� �a�q���FS<=z���OeW��?
f}@}|B1s�06�5���SF�b� ���T��m�3�z�j�X�����%���g%ҏ�J<6'!����r:���^UOQ�/Zp*w�C7 ��r�V6za�.�U��ma0�M�%�Z#�drƁ|wz�/�P-��8-��;*e��&�o���5�d2ڀ��Z�U7�̠���� ����qYU!9�G#&�.��\)�����G��M�#�Ɨ�����NR����h3���GI`i�-ꮯ� �����\��Č�	ّ'�@l��!3�icpŬ��W���k�F�n/�XjG
)��7�wH�#ǳ�^
�r�.��O�#�BeC<J��)�f�_�ɡ��5���z�4��|[W����G�����Yă$����V���O~"=����A��s�d����֦ݏt�=���U��F"�INrw�'4��0į+��b��� T)w�}EK��l�)�y �#~�.�G]k�݀A�N�7�\$�c��͌?�����t��~6w�o��U\v?et�,�ێ�a�iy��t��~W�ݽ��|y�~Ge<�J's�Fm�wN�Ϩ=�cr2�~������$��Չ���
4z���$@���o#o�`b���p�TB��(~͸�Ī:��j�:����xrmУ�ӑ�~2n�����<�z��^�[�����S�NX�)���DqY�s��f��#�l��Ⱦ��c���Y���)g\��W>��<8�8NP��
6Vr�@��2y5��.Q�Z��%���<}�\�,<�z�ͫ���p��q����m#������������zrj�b�еj3r��Єi|§��"/�Eb�CN���"�������H�Z��J��B�w0]~
Gu���ҟBə�<h@�1	^�1���.��xM�
u�n�>b��ol�o�Ӌ���kQQox��ٯ.�JD��:�A}�+�͌>S���t@h��xV�D�nrZu@�BUDv�L!����ie��TK�qi�l8��瘺i�� 0y,=㪠��@���6��e{���)�kL���yؔe#��~�N�A�{������O]e��O�x;���9���א��<K�W�.���c�ܦ�&Z��4��ͪ-�V���#���{��Wc���u,���vo ���p�<��Eˊ"��>t�`�X�4 �۵��{sV0��9�n��[�$��D����/�&�K\���*Q0���C���!N55S�E�>%�x�짰��n}�r�K�?�ۖ^>��9F}����*��iQ!��v�1��o�i�1�d?+TDӁ���R���{��&z���~Or�\�}�nf�"�8��R���� �r�o's�.��0��B���L�����L_��:ط�b�:��|+=��-���\,�Ձ;��u
�c�v51��^�诼��������PB�Ⱦ]F`��U��jC�]�^f���RsYϱ��DSe�1V
[{�j:-�t	�%x��=��&#�pH"�-�������f�9����(�-6邅S�Rd�n���r]�ǹ�Y�0�\dp���,S���"��0���5�8u�����/(˼�1�	�u	3D�eY���8:����DDP{k��1Άϖh��%����(��I�--(���1ޅw�#)���0$Oy����2�[M�7���D�P!X����Y�8��b�fK�������a��B �Ռ���.�ݰQ}�&/���0����a��¿DGc�.�b[�y���'H�Er�'_�=C������$��.H���Hhe`��-:�l�Frc����_u$σ/��i��ջ�:�Ğ�_}�Shڭ����:��[Ƣ+2���I^q�;q�W)ʄ<ʽ�q�Lþ �]���e�d��o��M�(��H]^����l7qw �׿9��z�H����k����|�(`�?���skj�g��١�:㨜�8�_Q
�y ՏՌ��5f���+�2R�%Bz��uXUm�{�O�[���]vԈ��`͇ƾb@�URvk�{��+#:-�~'�xb
b�rL�,j�mZ�Y��;	>oCD�wIT�__fgt����H;˗�md|N_��S��"tU�w�v�Qw
�R���I���H�S���j�.��MN�W�YKl_�:���q�AI�2���l�g����z�O�M#�v�v��&����H��m��{�4�Sv��;hx�U��<-����o���\�Q��#���%�	HR�]}� �m�A�"���} �"$�fA���q}ͨ��zb�4�K+7D#b� H<x��n��G�~��&�bb]@H��ľ�`�kܫy������S����E���V� ��Kj/ڞ�H�Ӭ�}r���	��rzkE�V7rqS,�J�dA�$��^;=��Xd�#bN�6��tI+AE�+lK3k�3�� �g\T��T�{̇@��t�֭�����^���1��4�~��)��Z$Wr�@pP,Ys��g6�7U��5�,4�լ�5�G��P:z?pkܽ������ၡ��'�l����V�n��� ��ѿ��E������tm�KJ���`Dl4V��z��Ǎ���YZ��Re2� ��[�K��%C�('|���Y����>>��5/�m�oF�Z忖��~i��NL��3�����m���RQ�DZK�?]j�\��:/$C���f*BX|�%�Ѝ�x�׼:���|�=%U�ʁ�3[����Ny� {�x��/��2��Dnw�`wn\�����o�9���ķC���ڤ�]��8S$Iԍ��F�s���2>�mW,�d̚j^n^��yc*AJ�ŭ�X�a{��mՈS����Uh�����)���Z>�4�f�Ҙ�����Ë�W�D�Y69��PƘ$��͔��J5P��mMe�z1)?J�C�:\0b�t|��#��k?l!�������Ssu.���Ԅ~��kH.1�@�u𱳇ut�]dvy����^��-_
;Z>c�"�Xa>`��f��Xė����J#}��L�rN��[�jO�FN�\��
�[P#�%���7��c.���3�=q'�H����qG�݁ ����b�$3���Rݚ~YW�	}����Ej���c����k�	OE��S�=�-�:�������z�?��/��WvE8�YK�=>�4X�Qo���b#��*1o��*���KO>6|�94HN�_/�}��p�N�a����H����nu�8A.q��??�������q�vS�6̱/�|��6He�I��H��Ԑ�-rnk�#���=�M٫��$�f�Ű,'?��DB�M0.��k�z�}���%�^��	m��$Q~Mz>j �+��j�.�����V{B͙��af�Af���@A\ehL�n���xb�I���ݷ)��|P���J�6h;FpD���5��L�Xd�3��!�?�� �{	c�7A�w�����Smc�CWk���`�N	�|�
�X�*��YŐ��n����)P�'��F�a���%��hm7���9��-n�����ݵ☌c��-O:��_ʦ����*) �H�u &�EևL�v������muȭ�V�0�!��D�����m�p�7��z��`�|�={Oဗ�1��4w��d?jڧ>�>@+���C�՗�rOH��K�e�;ȿ�
�z��0N_z�"�VM�دߘ���v8?x��xV ��L�����ۉ�Iw�j�1�Jd�Ͼ�SK���Ҹ)��!]81�WFZ�k_\��AR
���G�/ѓ288�EN�A@�ꓴ2�)V�
�_&ӷj�k��ƞR�	���E��]	�'L��*�"�P�w��@;���6ɾ���噏��%��3�9���m���M4n8HhN�l�����((��q^��OStP��=��7�p]% � /1a�F�K\�&Le�Z��S����$�J`�@K�3I��č%w6W�CS�|�3u2�A������ϣZ��^����*��}e�v�i.TX�j??���S��c��Y�%��r�2�9�XA��B��O���o!��N�;����E6����eϠ��!�')@
�>��,b�y"�9Y�5��ƀH�ނ[�:A	A=z�[dj��vA�>6ۺ �*�g��#~���gCN�l�Y6|jX��8>-=&���-=Z��-��j��x�I15�Wc8:����8or�i��}�UYkp�#O�o�t�<Ip�˦	�K��
f��׍�(^g�D�u�hK�w�{
E������x�+���h�K9�&�I����\]_3B�f��+�G#�'�B�I��O���'L����:�K��W�@i�Mry�7-8|~�5�I�5����{�����}c�$?m�T���Bo��B��&�SM�3���0-�kDd��ӳ<.,�i�	�N�`'�3��tʥ{?��~|Ɲ����P�W~)�`�^G�(跹j��([h|IwZ)BR����!e?e��D�^f�O�@(nd�x�֯�d:�1�/9����$��P��Y9��9��Haʢ�#Acn..6��D�����)
}�8�����c��4�=��b�?QWK�l�����)�Ҫ��!I��S�7ã_a�b��@`�X�GvA-΋Ъ"c4��9ㅙ볓I,�7���P�����9K����E�tW�8hZ�`B
�*`P�)���,s���=^���]b~��Q����&F�I�&&�W���{{�yn�%�K�
��?���?���5�,D��(iΏ�[+oᒤ����ϒ�ǃ�H��v7�R�o���}�k�ܧ�N4�q������.S+����@;�B��������CƂVWkC:��6+e[9���� b�������������a�g��n�$n�L?B�X�ທ|*23 2p�L����J�m.�[u���ldB�=�p[��ݭ��L�-�I��#�a�e�E�x*�EjZ}�4Y�ܦ%��� k��4`+e��L�@��Lag�a�l� ��P�>󫖯�:��IiKFg�/J�%Ҿ�o�Ô�v6�2��wuL91��p��7q��/:f��"�����aew��|��^>(�0F�I��i��%��;��4����Wut�$���E�]�S,$�\w/�PK�ɬ
��\�ui���yU�5����kGj��B�X���nU!?-���,�}�� 0L[�I���ȤDjp����
4J�j�c ���'�L��wV��ha/r��x��A�h������`.�CR�Uk��l�Έ�6�'K�X<��W}/��7��z�o��v$��-�`�Y���i�a��b���;�!5�MX�ﻍ�ba���5�ڔ0-��Ž�A��|�}�E�Q��`K�f��bU��N���15m�U�K�"�N�,`{o�M�j�6����UUFK���=�_~cO�p^a�@�%�z٪q�!^.�_�s��*��&Rq�QP%�Um��BZH���Yѝr�o��xJw�?�M=uU�=�mbS�m[d��S����Iy�Wޚ����!e���?�h�B����YCټ�ר��x��"��?]>9������ ���B���b<��d�$7�e\t*\��-���g� ъ��aK(Y�#ܡ7ZuV�5�i$��cWN���zck�M�k5ÁF?y@�y ��5�퐢c������7މ?�:E��5��Z)�`�kBg\����L�Z0�^"��g�b�z�AsX��6��Fh��L?i�~B�f�]�*�B�΄BjLD��T��i�����r���Kk���̍G �,���=��0�H��Ls��M0x���5b]�V�
�z}6��F4ӭ5���/כҳ�1�9P6`�ѷ�˿�L����3��tm~__k�g�)��u��O>u�2�C���aʭ�-�ޞ�}\��x�l�y�:�A{!_XQ���+����G͍y�Q�QDM8Q���2����@�Q�+���
c�I���^��)�=-�O�W������J�}���~�1W��d��Ɣ*��nT�W:��E����X���n�4A�>��R���֜<:٠q�S'AQ�w��G��(Ug��[k�ďp_���m/���DD�[��6y������!wXVeRF�rv.���Aь�iO�� ��g���A�];`9e'�����!��8n�%�*�}̏ y���e��>K'߂�*4;J�[�ƾ���/�e�t4I4T�H)s��5X^��|�A����iD�z��II��{,7X�V����/ 	 j����z+�J��[X�Ͼ?DQ8G���y	�s]'h�~�jZ�, .��
���k!�P>@��~ѩ��G��'��`�����BW��T:< W#�?"Բ�W�i�)��>���^������<ң4�Cp�{ޅ�/�������܀�g^�>%,|�&��:�2ud�!��y�ja�o~v����/�e�!�(�.{�-lH�,(*�s��'hM\Fn|����	h U���&�e��h�?oJ�W�:��t�̿����O��a:�iM
>h��#�+�o[��F�^��2�/����%~�
�ۙ��p�MGՇ��̿T���aQ�T��z�[-����S;k�(yS	d�%�����ȹ��ĸ}������Co�q�"�3�����2;��9��x����(�2]Sr�
�W�&�úB�h�X�;������^��Q/��T:+JW�\�/<�p���7�l�98�"PC��e���\W���c����Ͻ�ڝf�k��c�B8e��_;�R�O����T��1�V����Y�0���M��5(]-��=�t��5���X8�G���\Zf:u�J(��[-��)�`�����m\#�,5�^U&Z ��S�I\�<�^��v���@�����
�;���߼8�������u��ġC����vH�c�5! jYih�/��?U@�[�½'���\N�*y�m����|���2@�D�BW-y?û-���#X�nՂO/#�J�zT[�����r)�����Qv�n�V�d�un
����#N�8M�ѕR�l��+Һ��6ڍ��#�<+�.�ݝ�:b���	i�t�d�\ED���ԯp3��A�����#?
�����M��hI�޵M㭆�S��S����j)�.���-�VN+X-��O�lK�v�٣�����DA�=D��ϣ��[Rd#['�[i9;�x��x�w�w7�W���Ag�P"n�H����~D�U���Sm���⅕�����5��,@�9����.C�z��$e,
���>��B��m���\�J��k�:����!�{��/����8H=��F!�)�?� �C��pY����E�H�;6Qy�:���J��
K`��R���$x^���T!�� ����2*�L� ^Z"�'.O�{]�����E��������z뇈�#dQ]�c�p��4*��Sh�1�?8��\[��DkIP3�Ω��z�N��"3%��Y� �aTS� &�B�O��
��p�X�L�^Y
uS����) �讱:�㵝�C?ZA+�1:�?j�Pv���Z�Z
4���-�"�G�"�I��rlQ[������nQ�CL0�����bo=t�V��<ާ_c+�� �s�n�e7��5KO�J�tA �L��m�"�T72mJ���b��� ���V��&�P�%��9&2q�	,bAf �-�U�����W��/;�HuLLjr��O%u��9�mu�������� ���`ure�7���y�~�?)��v������� ta9+ÈD�7�M*��z<��Ĥ�9��K�	_
Ӕ�y�ם\G�>&��x0b�>���ʒ�^g�s�w��v����֖57:"W���0C�ݎP���eO�[����
488X��hi���G��)��
P:Ǉϑ䷁+�A	�B��⣃6G����C�#��:^��@�+�O�t��F�V'WQ�	A��
��>�@����.��b�Jn���S�I���p�����φxK�9Y��e�֟��~U�F7GS���1��U���H,�V*�\�����	�'z'�*B�!��7�nb�=���ȡ�Vac�\��E�_�"�dF�/�u)�7�����1�w�������/�=R��9z�#2��߲8%(f��B��Ei�����C��ۼǯ�@����_�c����)=�q���i/���ƛP�d$����u�9쪼e	�m�"�[4{�����v|?i���BѤkE�����ں�!wN�S��(����;���b�w�͟�Y���Э	��Z3�el [+��������?>E�� 73�ae�}���_��=�����KƼ��1���&S�-�ĵ�f�+�ЉG�p3*Ә�E<
$}���u����=��>@6�#��\+kQn�ha`�Vnzݎ>��Է�1��Ҧ�0_����޺�*Z#c5��m8��ME=K�Q�m:����NV4֓*��|M+�=i�pL=�	
���W�J-�d�;�x�y1��,���\�E���6�ya˧�P_#�Mt�R�(�A�B��n����k.���ˇ&e�F+n r� ��U��4#z�d�Vˊ�V=�H ��D�jqilzb萉�a�n��eX���:�g��;A�ky4���y�h�N�oѳ�_B���Em��"
`�[V-j��[�l�+�(z:׃�fJ�ҷ���D���a�"L�TX��𔫛����!�TT�G!:;oP�� %R!I���C�s;X.G����#Y�e�R���G���K;B$�yl�L�3��i��8�D�;�Z�jKc� ���L���u�?�^����h�쾣G��6�PǞ�Ae��4�q��
��<�u�>o�B�Z��r�ݣ���i�G8�{@m�M��:։�9k:*�f��0��bH^R�k)��	Fd�[Հ�R74&2.�w���1�/.�Yv�f1*5t[7٬V>�M��/�'�=�Oy�=�����b�+ϳY�ct�š��LZ�18#D��I�!�~	��0w���8�?�N��⒛ӁM�/A�<-�>���:�荏ۀ�p��Z �cs�@dYܭ�,}3\"(mr�	��P���W�q��i��#Yl��P$O���9H����Ӧ�T�.��c$�J��C�Q3�]���J&[��C�B�Mg�:�h�X*��4�NBV�-��z�RۑM�p-� �����ī�4�
Gޞ��XA� �ZȚf�����y>ⰻ��a�5��x�����o
�s�5��G>��I�"�?����0'�0���M"Ͻ�ÃW0g"��>*/����[���t���٫}<>$�b7��2G�Xx�h�'�p��H�>�v���M;�I����!=�}��k�! :7��]��sT���F�h��?�^���3-�� 3�O.U��Wh*F��o#�V둳�>�i$����u�w��&R���Bn*^�̞}�]�&�3�w��Q�8�=����hC�S����zI�.(M�����;���3)`J�$�n��7��a�i���"JQqEW�^g�Ma�V+��5�ۋςD�~a�3a����gC9%Нw�~&�%2j���������u��H}|q�*�o.� �z��1��ȁ2a�߾�	Ð����ZM�&��
�75(�Y�e���D����z���N8����0�)�qR�;Q���he��Dh�ܸLor�DV3�?p��o��*�L߱������zY��U��8�h�f��-�-�5�,�7sM��D�_˿P�dtb�h�`d��κ��q�6��&���ɶ���jsp�)ߢ3�K~_l�n-��-�)����%���ojv
�l�7|Ю��1S��by��g场���'����r3�� \qΦ�r�X�P��៷�*&b[��Lj$l\ml��*'��Z=��6d����y�8�z�,���.&��x6g�E��u1���j��E
�l2���$�1���:f-WX�2oE!��RW^p�(/�"s<V�[ܩ�Uow�]�������|�kX���q�tw�~��
���(F�d�*�,�Ǉ:l�F�VW��tF;q�'}��{��~;�j{W�k�$��D�����Y��ĺ��>k��K����̊��E�kJ�ͪU�T���a�'<bu�b0m�}���/��� ��˯6(1? �C�ۋ%f��) ���i�"��:�Ҁ	�fq���d��QP�����tT��3dJ�� M�����8A%�K�BE��
�_JG)���VZiW�?	�:������^m�d@+�� ���*C@T^#`������rMi�eH;����j������D^Ʌ#w"�^�iK+*,��Pk���Θ-*��Jͫ�Ϣ<,QaMo�3V�vy��NFb��n.�����j��d:-c��� Y�k�<��ry=���`���5B�Gqrp)���Č���S>��9>g�H�X�s����
� �-ݡ(bY����%@�o�G�t0	v�J��/�[4l}V��s���U `9��E�ܱ�! �_��	z�0���0��!��K��>����#*��d+X&(����;}�?�a���LpwT������T>QH,:���}b���0sAIe����ӃmZR�t�����'d6"�>��ׅrQ0s��X6M���X�8�}�AB��>�_���C�8@� ���b�<@��͗���,��g+~;x�8��z�n�ޖ��S�,ur9j� ���������]j���̏"��1�,����_�	��V<��6�K5�A�~�Mރ�d�ƣ0�S~�����vt"i2���c)�X&��27��x��a�|�P���9u��eE��q��)���8���0x�$t���!� ¤�lC���K���w�.	�9���ц�
�nSt׍�;�av� \%՝ �M�d���D��Nah���ܦOie��T9�0����=v�B^��wRN���t���2�"NM�M���L3��G}z����Yv@*छ>+��a��J�������xP��#6�y�G%m[#����7�,�������4
?��yv���K%I��E��MC�x��ʃ2��|���|*�Ƕ�+����4��IH���#譒Պ���)C'�l�d�6;?~w�"�&�0���|Ơ�?�H�Z
U	��~%tG�~���x^��'I0���Z���G��0�Dr�$cWU(W^�^�����o��=�6~��1��b����A�d��:�lL�%�|���u�Q�|�*�Q�5��G�E�.��tk�7�D|��IV�^��ڽf_f^�ƿ�F1���ϥj������eW�_!��z@�m�c��+�)�9���/>G�n���@J0:�������0\�;�cB��f+��E�㵁+��Ŕ]�Z��Ϟe5pE �q6`؄�w����`я��A��6Xe)���c��o+�5v��S�X��KA=�D�]p���q0/T���Tg��mph�&%��ȗjcB����$��*�LA���� ��l/U���l�����~��TPn�W�l<�|
Da*�F����K�������<{�H��cX艣���U���@28��,�ՙ?^�O	SnF��$�hH�k�9��Ϲmm���=��U��W<�#�����,�<U����:��+
���F����Z=YI���J* &Be��&�,p��@{1)�QwIj��o����e���=��;띠�S���{k�+:r�z:��{=$e��߃+O�z]`�5`� ��0��� �1k��D��?�sC@ܮ��¬�Űɀ	 ڇD��*���bQ�ֱ`m$�t��q�� n�{��Rkj�(�0x7&t���`<H�/��ލ$��1+H�ݷ�V���G4��K'��U����Gh@J�p����u�3/]a#Aw
M>M�uʴo�$�����q�m�뉺��aS	<��Ǉ�%P��?C�ŬJ�/��2���w>�����l�A9̊?�6 8�h�J�<�:Q����#��� �7�������S��#���~h�!N��=��Bʛ�?�-ə�d�!M?:�"��7����@DL�!�c�N<dV��фp��y�}{M�+�T��ڦ�3C��w	
�i�,���V~�&�5/7��-6EPR����j!���=������|�%����q}N^Ua����ՠ�
O;f��<W�	��R��cיu��d<�W����Ǩ���n��v,"�����$��@��	���I�ɯg]YA�?ŝ�*�ꍉ���!�P��߭,*,w���C�SPД�"疠!o��[χ�U���&���������T&���,���E.D��}� �0� �MIR�@aav�
�Ht��ߞ����;_C�I:�����m��v�=��5��A�ւ�a,�~�0/b9��9�����iſ 3�����}z�Α[��;�t<�,?�t$I���a���sٹ�+_����������	�-�W0���W�U���)���]U��'���wRS�&���Q�-n���~�L��侩zp.��n��"�iq/�k-HFjG*�9����& � @Q��y_1	LmJ�H,�Sg�Zw���B׽���/�?�"�>̩��]�*��#���Z�OH��V�~��{�![�P��rؓ0�F����`�[���;ʵ�O&�S(￴��Á����o%��?�wۍ�R(�=^�B#�'�s+*,��U��s�$*c�ѕU��<U�f�q��?�t,��B�"��.�u�t���%֬�19J4�F�ꃝc^�2d �s�(�h�J�r�-�����<<�6N��	��6H���E�_��!���^���w��>��:%.���t�FF,k��/ �f4������J �oU�'#��$Oa	$�P�¿3ڧ����ȶیc��3
��S/#Wť�jɍA���������@�F����j�kܹ^�o!FѮқX.�=X-kJ�ԁ�Ke#w�Hڧ�q��MT�LG�>��FC��r���� k���t�_���)7�N�� \�a�M�����Ja�#���%w��h֓���s��+��f<$�����U�q$�h(�tpi��!)~���?��5	�����*�+1s�	/�fAwO��ER�v������5s礬�(G���bn�*�Zl/���h�{�>]�td6�<���#3W�83�y�@2]k	JVba�T�q���Y��s<�,��TӁ��*��$����R'Sݬ�lV���lc�ٮ�d}g��O��Dٲ\�Ҋ����+?��R�RW,wv2�E'�pw�4�����x|����1��݈_\�c~�y��E��﹃fo�)����zp�=Q�|t������\�VZr���F�JjC�G|��J��nh[{�P/b�E���<�e��p���g8�^I����K\N6i��TW��\����D�N3IBPˠpQ�#�1<�^8}�{Vv(�M�@MD�DRi��H)�AZ#��aL�!KHg�����V�Ě9(��34-��v��4�j�M|���SW�}�M9����j��:AR<y��E�!lg>��5��2ȫ�8�q.zW���������J�4�];^xC�����=�7"�EOs��a�_��T�p����T����Z�A y���ݷu�W�{�R�O��¤%8��K\lR��"]�����=l�᪶aU�Z�^�Eȼ{�m�p%����:/�-���V\����7��zA���1��Ż�;Z� �h�w�E�^wk�B�f.�Y�^9�%�v����F�$����#�&���f_ts/�mՋ��"jl�!���?ᜇ
M�à���]5�\@����OA6�����poX��NmpMI�`����-B�/�a�ŵ����� 6�e?��$;NT�J�&8Sߤ7�Mq��4�c��įA�V��f��m)`�&xI����'�Vj��"ل��(EΧt�w���x�6�:g9�`yo�p �>@&��weٴe �����}��x�a�w[�Ҕ�W1W6y@>ܭ����-w�8���=��?>��?�"�Q[�$���=������µod����S�PԡU��Ȧ�ۨ*~�[�y��%1*��R�;��D��r�Ġ�gO���V��j�p��j���lf7��֐�>A��� ��|�i;�^X|9+��%�Ewd�}e�U�&X�B����rl�Ǌ�B��M>CU�p���>$�v���]�׋�u���kxsC�G%����H.RA ���;w8@�"�yd�޺E�����nw�	9�uK��&A��J�hs�WF��蘝��Q��^�
�O���=�M�xO6��/���8�V�&��)L!n(XƖ�_�D�N���޹���2&Z�{�F��T=�'`�'L���qB o�J�>=�r�,��$�>;�P�s���t�0z��s2�� �I�\c
�� �Υ2K����<�z1\]`��0�G�CBw�s���V?���Ͻ`����x���Z���ܩq�|�`�ה�B��4�򓬡F+��S��U��'��fl&�����h?C0;`�9w:^,�fp�<.�i���L8C��჌���?{�qǞ�`'4)�	F�4�/�W�����s8(�A�� B!.�d�P%��[S��,�����!���+E]Vnߟ~D���[^����E�����gRk�U3�pX�j*�ˠ�W(��p#fV��nN�fF��Z%�� #�F6C5 k2/EO��,������^�3����x�E8�Y.�OX�I$���A�/V֓��2[��IR����ϺX���93��vf:E����|�ݜ]	�AVf;s� �z,8̦��|�^�����G�}<QBz͡#���N{���c|oT�ZU�����9��h�ܨ�c'Y32�������	[�ڊ�g=�f��WA��E�=�LPgmj���՚��&���0�Q=}�7�S�;A��Ё�QY��� ��fi�>�H>"2�o5��L�q0����m�����"�Pҳ%H���<O�����V� ��w#
D��+N�ɫgA�u#v˰�J��IdAv�M��4��dXJ;ګ^�7��=�+���BQBi��="2��<�t+l��H�����9��
��C��B��D4��_�ҟְ����G��.����J<����m/��&/�d[vI{:!jOo��r��<��Ŝ���}] ����{���tH?�f+x���
H��'�#<"�i�g�u!�GՉU��gR�g��@v�O��!��	ݿJ�!�D롐��p���
�<*�˧ܲ����_��Hٴ��o��W��:��s�N���u��粨�a@�}�Q���O�3��'gL���猱j{�}>���Vo嵰\�W�J.D6�*�󺁩�S0$�>��V)�rl4k�B�?44��k>�����];-e�������&=p]��vn�4��K�M�tfR���U��]�0KB����Ɇ��É�'l���G�q�C#�O�p�V+ 瓷��N6�̤x&���B�E��w�2��9�L�
3�h|е7��>�ҹ��9/8:�!`��sk��Z�|j�Z���1� ����@�q�`G�ȃ���^����v�V���s�7��P�k�o�}�C�ӣ=���#`�P�6�ƻ�s�<�.��
��H�D�@ ChmS Z�h�����H�՞2i5�=�Vu��=�,R�ێ���Y���A �@B���[L72����4�e���XF�yԃ �a�?����i���ȱ��Z�����p.��5{>X��C�daL8(D9���1+����Ē�r�k�s_B��_A�o�4� ���mxy�K��V��1�?�Mwl�K$�ו.��[�t��Ý�X�����|}D2 C[�.n�7�9'��6�0?A�-	Y`O4w���5��,EC�˽8��nC����SBމ:��X�@�:{/�e�A{�-<X��r����ox4Tt�!)��E� �G���k�3��5L9��5�Qg�q�L4��"��s�=$�<Q~�P�θ�N�+�A_�^
��{�f��R`ׂP���3�x���L0*�"�������ҽ�C��0�?���F���.E�R�H��F���G����|���r�^��x�ծ����lU�'�`��hy-�\ pß��<E���x��`a���_D�V�9����9���R!<SC�G�*2S��:�B����:�@�N��b�>M�m͏$��<��j��D$�~��˵V�w�d��=��sh��T�b���������5B�3�z��m3���ꋜ�co?Iʯ�&̓Cml@�B�ջ$o���Gs��p�̡,}�W����N� ª�	�$�@�l=�����7��G0Em��@�F��}X/�.F�=��䣺ha�9����w��D�ō�����A�A