��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���}AW��l��&�zZ�#F��h��(!�b1�{pE{r�_k��08L'��Nx^`D�z������`��#�I��E\E�`Ȋט�;�����W	�		\jя�����{�h���q�'�ѵ��0�Dz-��a XQ��+����WT�n�Y~����^&�!���ߧ��Um���0鞱a���F��{j&��QCI��h|�E�:�=���:e�M���J`yi�~�p%,G�_?���:��I��>$[,�����scj���Qy��׏Q���:b�N��P��N���ދ�P�O��ã��k���c�k0I�ɰ-c0��9r�!�+(�<���[y�9s�8��]��Z�L'l�g�M�+f�|x��`�aI)�{)d�W�?`�����3�mbC�R�j�Ɩ�
C�>?��iZ	��=y *sj!)�nԻ���ǚW�@��X������h�l�~{�Eؙ��+_sz���
��y��[{Ƭ(Rؾ�<�����#���W��i�]�5E�N�u���̈ʌ4bǟ�X^@���ej�������-���oS|�-�Sk|c���;�z��b|�Gր�sV:��,Wa兀����d��EF��Em�$��kɽ;Kx&�h��̀1[P8/ߌ�ta��
��kT+JX�]E%iQ�@�V�4�^�����r� � d��G=�e�-�f�,��M6�wצ��x�<���Db[!
.�"<���81',�Z4�-�
Of�9YX�8�GYM\��>ﶉ���Ok���
������@"�֕z��������FEnb��/�K����0�)�B�K#��7�����X�tu�I��:9� �q2=�b��yR0S4R�\΂�	���p��4��"���*���K�y"e�O	oJ9����bދQ�Pe��%W/P��db(u<k~�HD�l�r�uDbi���[�9�wr�����uLt�L
���x�7D�q�B��,>y�[���Z�}��6m$��gtY/)��P�t���aH����۹�d&��]Ín��͎|uS�*4~{9�m�|ɿv.v7әpMm�z[�+��3���剾Ѽ�D��"Y;D(4��K�|	'4D*w��ܗ��o"����`���f���&�~���g,u�=�7��ub�`��TyT0��;��}gՠ�F�����|��I���u�	�j�e(�:;aq���7r>��V����r1�;\ �ق�\]筑�hLq��f`���k�'h}8E𚿝-ڗ��f-�g�]�����Xf�~o�Ap[[��Q�;�[�3�d� �!L���;2�)�ymɧ'�!� ���T[kع��.|,��Jt':r�L-���f�s28�Sqc��'�~+��2z�PE]Ȱ�p�������&s�v��dX(Q�ߞ�mx���OM���(�Ѹ���r��9���ӹ-j�b��q���I9�O��0�i�X��͑ϳ����ƌH�5'�NϮ�@�3�t��Q�2XvAC����5DX�E���p@"��� ��% (Ǻʼ�\Y�1���Pİ�M�R.Y@A]�������ٍ���7���{��߳Zg玩��]lY_5�Pȗ��$)ѩiX(�סe^!�.=�	���Z��4-�[P���?��э�	���u�!��1hAN��)����U��$�jc��
1Ĳ3����*O<ȶ?n�f�[���������j���r������h��L�e�9!�1�z[����vF�� ]���ͱ̀�\ŝ�KbY.&(y<�p�K�'BC���a70�/=^=A�3��:G�׹a�/�`$rU[T�����!�	�-��rD��{�,K����7&K|�y�H�nͣ�Z�*�]>5R������<Hо�YgdWC�.��U�e��1������4Օ��҄�G�?�z�����×����O�Y�Ga�*ihg�>�/����*Oڥ��T��fU��	E�8��9u]`��	�t1�V�^�aS6`�D/ � 9l_�+�E�t���(Q�j�x�������l���(�= ��%�;��Q5t~ݸa׻kL&�d����9=9���~�Y��AU$���ֵ���'U>��WڰP����
�;�j��v�u'��V�E�OC�f�E[D���K޵�x�ty��H�@��K����D�R.t�@�蓣��q���g��"Ђ�$��]��z)�D�,�&��x�8��� ΀��|6X�*7$@�O�۞V�rnߴ�,aoO��"+��i�q�`�R�e�s�����1y"C�\��c�
���[�Xy�����:SG]g����	���q�е"�C٪����A;�x��lD�ݱ.b�3/u��o��Z����C�Ynsr&c@w�!��o
*�Fv�(s[pq�$��U�d���|Y&b�o�9��x�DA�*��ޯ|2�u6k%o�m�I��Ï<\ ���ϟDEAQ���w'�q$���:$O���G��+��Z�P��3f�"�@��k0?��5%̰�:�����h�TRӪ�Ϣ++� �(��&��ҁ}k��q��7dZ���'S`��em*l�����$r~'v�7DLb
�eģ^[�4��������$R�`�Q�/�ɴ˯fF����̣����� ��=&���T�
��|�|�e�!