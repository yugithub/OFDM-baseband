��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J������`�>Wd�T@~���Q�|�w6�v���U��!��[4�jtw#5�S^�w�5;&~��j����lh��ҧ�te0��!A� ����.�3��E�O�[�߻>�N{z1GY~#(v+�d,����ğd)�þ�#�߲z�|�zḻ�?s�(rm����D������I��.����=rU�O9���=3�}">�ϫ��Ѫ�B\�{f҉]���P�vq��ﮰ��f�Դ5{^�Z27��R6���\8#b!����$�s�2V�n��-�o����]bj2-6Dr/
�),n�1�&2�
�d\	�sًM���d����\��K��U	�J�!W>d��Y�$F�l���Rݸ��Wh�Y!���"�E�%��jn�d��H>�,W�8�C8Z�2�r���	R�\G�&�[���t��Ԙ0�O�9ê�.(7��[E��L��~��v��;
V�X*��x�x�=w�|7Y-�QV��؟:�Z��}�<n2z��'�vz�������9M'Z�t�3�Ѧ��gM�v��#'���E=�:߱AG>��P�g�k�=Dq05��Bq���iq�i'������������{Q�>~&�!�>3eԫ�X9��g
f��~F�S�8" ��_�����Ҍ�����0�X��~��S�?���4A� t���t.��xM!�e:�_޻L�zS�E���9#ۡ�o/���������́�V���tNӦ�c�΁Rg��څ�#X}��^!Ί%�����ZQ��ÿH��0=��$Q������{�.��,6���k�M���0v7ᰓ2h���h�����3��b0��DS,�Tr(�-lӗ�^�cE��.!��(