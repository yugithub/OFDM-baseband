��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ��������LK��^v���5塞�1gM�Wp�f��	mi�b������=�BfK\��|	���69�]/N^1���>/��L;*b��䬑�יj�sN�f7"���9Z�&�hZc�¹7[Ȳ�;�CƲ^M��(�xϽ}�bk�n��e�.0/qڗk<�O&C�K�>�v{���Vt����&�5����U�R�t��e�6d!�7��y��&�u���K'�������˙r�  A�غy�'3���9"f�b
��N	���o��ѲqL ��H".;�=hx��T�$���>>_�ʡf4�%��4=C��+���qJ�)3x�1��e�e�����@�QlQ�Q��Ǳ�L������!@B0X:�����R��x��j�X_cv&H%���� ��V�ŀ)\H.	K�*H�*�--P�]�
�(�y�}�!EB�ǩ�gk0q�8�%Ak_Nם���/�s �F���a~���8�������n�ڢ�)<����æ�9�cgϫ�)q �žAK�톕qDڔ�r�<�\B`��B/y��'F�g�oу9���򬸫���h�̺�(�^��о���حN�g���s�=���U����OH�܋��ĒI��pt��C<�Xb-�i��G���wy�:fd��X4c�����2	�D�Z���Ռ��L��GrK�3	|����)�f����ߋ��.�6�9b�.f��H�^z��1f�����\��	�AX
�P�c���C�Q�l)\��f�~�p���{B��#�AC<G�g)A�Ѕ�M޵�WOx\���K%8���U�r���f�vⒺ~՝��ؘ=8�����s���SJhtV�ȡ�D�6�}��6h������k��w��_5�~�ێߏ�P�"���B��1SP�\��9b-'S�Z ��Ea��(8G�|�A�`A��"
��YP �E"k?u/5�Y���t+�����s�h{��~y���\��=WR���!M��'�O��K	ы>��14��Z�'*����.�a�M0Ǖ�v�#Sl������ �8v�a��.M.S-�9�gV0��t���#<������uk�g-k�r�1u3�p�8F7bO�9�ښ���$�V	�s�h��n��a���"k�5p99�?���@�r�ԇ�E6 ۟�uE.�՟��,�o��%�hl�
n
��o��[$Yi�խ,�!�~"��<��m*��������ޱ)h�,�J����7'~ֽr��e�r�я�yf`�^�8u���U]
'E�G�je{����Pz�t[=����Be�,�6f'�QL��+^���y���+�'w͊�eY�w*�&�#�% ZQ
͓�.	
c�=�@O��ZkP����j��<)����8&�Zș�3v���J����
�1�$��E�_�{b]�s�* .�����"����ۂ#�|d�O�έAT��y����ztD�4I��!W?��hk�^���U�*0�x�6`U6U!8���sZHjd
{�.&����J?٣�ҳ��{��H_�rKnPb;������ނ	��%�m�Z�� a1�WhV)GZ!eD
v�r"���%W����q�ݑ�/qI]0�U$�${Z�	r��l=W0�}Q��c�*w�Ϸ���|uXq&R� �76C��^�v��������J�r��\��r|��Jj7Ԙ���(��ɿiH�VX2�)�9�/��?WJ���iX,��iY�Q���"�I��� ?�6v2W[�J��L��k��2@�#�=<�r��	K?��7| � �fc�&~��4��Kw��y-�:�Ȉo������zgc٥%'Z"��~c�d���r���1}]vʰ�3�V a�I�����ّ�Kǵ�TIAj�7+�>��#=�ۭ�"
J��o"�ߵ���W���K�a��ƃ�Nt�T��$S��P�[^��'�����h��ϝ!z�����)��}��g���a$�5>56/|�G9P�϶���&+�$���K���U�RH��:��8�'ӹ�f��(��s�/>8��D�)���Yf}��Q �c��	W�A�t������194��sN[o�?�g�RE���������XD+�}�{�`�f<���+�bY����� �W�y���1×��j("��+�*�O0\��y�lZ���/9�`�t���4#� [B"��F�C/��2�<�53vu�Z�N[t�y�U*k`�hD��� x��JK!Z��t&S)^���!|V�ϲ���h��M�e���c4"Dʰ���b)�f'm��wbS
�i����N=�.9F����DfL%�5_!���'�%�x�FC!�=C"0�B(7l�\�M���(�΃�[?��	/�;�c��2�5FvU�N�����K�Q��('���X���Q�eԝl�?���1��!�w'�
n�YN`���锞5TW����0������S����)�٦9��IX;��p��c�xi��I2]�EP��B�7�/d�s�,叹��jtEK��Y��ٯg�S��Q�.ޥQ��"�����6;�6j�$}��/	������\�^A���`LK���/�4���?�e�s8���m��\
,� ǲatf�CR����D�^�`V�T/*Ӽ�-L�a�������3E/{���H(�b�(~m��;�����5��_rn9�,L<$x'u�^�W�����ۚ���RN���6��}4��KZ �"&v9��ץ,�(�W�W�N��c�$s������T#�\�ot��2>��R,���냬�P8�Yh��e�:qVj�c���׈�:��&�b�t��d
�JLC�˚0}��p"��6�D5����$�e:f�$���l�d��;�VO3�?�5��g��pn��/�z�+�0�Eq�/91�����3E�]�q�k)�6-�1w>�&G�� �i��g�t� �cp��M��;�Dp����$+6���	�����s��X2��h�ǰ�V�5�w4�q���sC�"�N�������5�ET� 2;"7�aՙtZ]��Jg	.\=u�Jt$�ۜ=>=�N����z��̞��[�=��Q����vI�*���ǫP��@ �Ψ�Lr����:y ��������TIX��3�R1?����f��?��q��TC?U#N��CڤS)H@�ڻ"����WӲr;}c�y��
ܹq���\��zQ|Lۃ��<�L�����]2�uUC�0�I�X
[c��IM��q˝��h���C<�R"Ñ��xD��Qo�����giH��&��Q��Ӎt��3�GY�V�`�X�����*j+��ACM9ZYG����&�`.|�M߉�>���K`0�*a����s���{/��)QB� q�`J��	�2���V�Q8|��Å�u��	ڤ�bD�䐮o�P���h���&~r�gdj���[o�(�Z�7�]������'�l���X�N�ug�80�����1!y��i�_��P��
"U����G��1\%�G/}Uz��"��2�A��3�FЈ�>޹\ n�ŘQ�6������{!�fy,��|��3��GD�:
Ћ��.��f�u�-LH���`���d��`���=}̞��I����H��U�%�0��9���?�(m�QuV}��o&ɿ�Z&?��b��v��i�L��,��L����@eν
�a������>�lK���P~H>u�io���M���:�d�P��c�ގÍ��[Z��2�����#.�ɘ�����w7���ћ5�Ԟ[�~�{s7z�{vtXd�4�*N�#]K�P�z��8����p�L�/_�4K���~�߸k>��*>b�'��q���:&
n*b���n�?��N
Q�5gp�.�2V����� :_��w�_�hPO�z�0^��*��޳�΋��_�"�9z[Bi���{���&-f�h� *挐CI��L�	��Ѕ�3��9z{es�3��OcP�w��0�H���t���}נH��4�f�K�D̺>�(�׼�ʛ��(�<hf�e�O��;4ꬕ�S`D⼃��znP�/P�5%���]�|Py��i�����λ��%)_U�]�2�|B���@����p�NY��������6t�/�@YO��E]��V֜�i(�P}Kzɓʒ�0]�I��霼�����) ���])��
�RW��v������B67˒�>�H�&ev�r�.>.i�����<Z�G�!�'�N�,RޜRbp̈9��S!��f��x�9��*�c��R�R	�q�.���Cn��\ȃ$#���HZsY�f��β��YS�+���7��Y�Z,��=�r�vώ|s弣�8����E%��s��ǏO���s�j�ĵ&��r�I2�EYV��aC1|��`�t����g��jlw�H�$��;�$vlZb=F�����S��l���1�E�]�J�f���t�̸&H�e����pA���,�4��rR!�D_f�K�ܱٻ���/7�.U�$]Tu�E�7U��^���B���4B�ehP_$�*��V$���O�3=}'��l�P9:���h k�� ����E���.�Q�<|pK[tu���P���"d���T/����y��Z=�e�����?��O���v�:�� cU�LE6#���; �pk���5a����q�<�\D��C�#H�8�d�li���aV*b���3�z���(V�e��f�p̑2���R������m���)�B
.�}�$od��+|G������4�+א-�<؛DTyA�AЉ�}�sT�F��gw�0я�y2_���ꧥߒ��Kl�y��Ł17}B�O�XY�U�e��)��e�H��w%R��F��7_���E��n��w�)�p���[(�p����O|�P���p�'��{�����Ms��99S�n��]%ؚ�X8_�C��z#��lx p��KPS�5x��9�jw��Q�(fi!�%����= ��L��}�t���"�cdQ����ig���`ţ#��#$O��'��2����h=�Ś[k���pG6��J�|��E	��a�3�4�2�&�O�5(�Q���a*����y�t���m���쁷[<?�ȃȅ��^2Ng7���,O�d�2�����x�:;�����L`6J�;�W�6E�x����msv�j���<����EX��:���4)���i��t�1i��9��N�<~�K��	��$��l�J���Hc��wÊ���`9���Hʱ�>x�C���yro Ge;)����>���n�Ujo�dq ��اe�!{�2vͥ�m��g�޹��|4����9���t*��sk����o�S�)�����#�&�,���n\}�i��R�Hy7��x�#1�/����2�C@�
�Q����Xp|�D�&`�!Ь�CV
{	Ԯ�5�ɓ�^����uE@�$ސe�3��f��{x�e�AQ�?������_
����\�+|n�'";@����f|��-ܫd�^��~�^	�,�!Pj�ec�"�����wT)w!j�g4�?^�f����L���L��C��R~~ld��-k�]�w5��آ��]�E����L����O�4Ӝvܤ��6� mޖ}k���4*U����N{�h���
1�}jL�1䫧A�v�d�z X��>
^4�Q��;<䶛����t��,��/q��D���YE��5%�8żf�ϵ���r2>v��Z�n���k��t՞Wך���n��l���@�Ը�����2��\, r��݀U ��v�f���3_�ܨ�	�\�?���Q��:�z���%�>c`p�gW�љ=n��B��|��������7�ܧ��ﱳ�J�i�f��� rL�O辧�1���i�1�9i��0^S;Nw<jmZ+����W,Y.x�5�g�
�Yx��\��م��3BֺU'�;y�J��~E��?��g�@�u�ܯ��ˣ�B~i���{�	~��?5
c��Z�����w�m\s�^��H/t��hA� @�/M�T���3g[`k�@;��ë�K��><Y��w��#��%93ȡֻ.=]�m�ҋ�/-����ZA�́�I%�PAk�\�)7?6��MD�B�f[��]+՞�V��!���a;��X[@��s
���؊	��i�u�hc.t�O'���gW��F��[ ��0;�S&lF�x8�Op�'� ��\�;^�Y�J]X��,1����;�i!�Q�x�}�p�D��7�uE�~�N���F܎�L��t��X@���d϶f։���"�Ew	7�sTD$�V��c���e)^wڱJ�U���;����y�5a����C����"�,�����Bg���&h�'�BJީ{d�+9�:T
��I�=��2L�_�}>9�&��
W7���^�r!dU^�9��=��p������@�1��yY��ӿ�YkH�<ME<�*��z&wP�i@�ʐ��
c��Xp 1�'��$J���s稪���53[�}Wbz��� ��d��[EJP���~	k�iB �����hF�P�2: ���p�/K�=t4�1���/��:��12\���@mT-HN���ĕ8[�la�w�v9�'�%f�ګ�B�P�　�TEK>Y5�t3჊�|��=�7����M#�X�;���E�nb�5����f\i����F#?u�v��nw��Vl.�j����ع�}\�p�ܻ�OFf�m>P�qԛ��;�l^*��d�c=�ZV�,3��8�
��xVF?��	�%�Cd��z�D�U=�L~���q^��i�v;|����Ͼ�x�L���H��c��d�9�r��Ì�}�x��)ef�
#�|h-���x��Z9�T�/�}���A��
P�ΰ�k9�pz��b��y��+�_�P��P�[]Ʋe��\D����n��u��>j�e\��l��	F�"�\�����Zʇ���ʬ���o΂F~Ʋ�ş�Ĝ�{�����3�}��|T˃�;�uA�`F�+Y��̓�b��o�ʂ'酆�Z�@a�v�6,=�x��
pd���s�k�ɗb�4��G͙���]����S��'!�<Nz�ű�����$�N���˩��s2��E)����t���:)��n�� 5�!"%p�Jp�����
F�P�G��O��@����W�3u�lU�s��
�����|O��ub��CDł�2�f/��ڲ�!a+cz�R��|��8/��@��~�_�E	)���w4m2��ct�Ȅ��ÜrIbg`ʉ���Q��^�BV��$�Ѯr�d�rV�,i�x^I.��fkf`.���a �.5{R_�����#9����G��[�|��2�O��dB�D�[1x�4�����,)]�U�M��/b�F���I%V�Ko�eo�~�,w��OP7a����y�xK+P��Lĝ�O�%��{S�:���lnf�_)k�4\��|��*�a-m�?(k��h�X�.����6�5�5,���Qo��<j��߾�����JP�J_���MZ��?�0�+E��� i���k'^�d&�\+�D"/�/]���W�+r�k,�����u<逤F�*�8�!����ϒ�u�q���0��;�Z�F�o�����W;�Cm�/n����MNg����`��1�/��_���])�`Ki>�L��*���BF΂�<���U��Uէ�=U��DJss�-{~��p!��}LA��*M��s`�����T6����s.�&��[�jիQ�r���0�`Ɔ3d�@�tǷW��M�ET�RI2S�ov�@ΞtZ	�=��ه�0mU#���y�|!;�v�U���Q��_?8�!�Q&����Nh[F�G�	N����
��M�-���j���LD.I�օ�\��!R}g/D�jI7P���c9Y�H�[�D�r�6�����SWO��飘�qC6xts�1���XNw�*����5%er�Kqal6O�*:A�Qu
��%:���!�;�q�xC�$�ڛ�V�LlN�����Aqr�:m�<C�̺$�?P�E�3�o�&Xcϊ�D~W/��`��D�r}3�i��4�;���whw��ji��Q"�w�P�y��c�w�[+lK�����)������U�8y`C�^��ǐ��%�21&�fT�`tv���ۦ�205����[�Y�/́
��r��^ݚ��͜l������ٗ�s�<�AK�"�����4"���;��>��?�T���6��3�2#ٌ��Zpě�S�P�բ�9L��X>IBC�(L�J�Hm�S�(-�9�ۦm��~�~Z:����Z�uhi�ũ'f�4J&~����kc��^�3��]����d���
{V~�8\C��d2v��D���S��e������"�y�|cDװ{�<�=��dg�ju�M.����P�D�gk*3`)[a�����A���ά(:al����yW�.��bґ�a�y�'�R�Os��sw��D�.X���־o�B�U��j�s�:��.��,��$)��z{�s��|q0���Ĥn�+�1�Y�d<oċ:���֡��'�DV48���Q���p�<v@�SdP�գ0Y9��{�]�[~������9O����`��/2�"�~6�ͮ����;�Ev�^ך�����47q�z]����@@���X4;1U?����&Y��8����rO���%y���Ĳ� ��>�7��ĭힶ(H��(��fi7O��� �|K�sH�0Wc�N�����Q�c��t;�H���b��D�����<����n���y�>R���v�N�� O3DZ�,�t����i>}+���X6����6�Y�t��5���­�R-�-��D�Wم��H�_�o��1��t�_����>w5�8��e�N�/�qQ������	���J��6�S�&�3��M�WLt��ޘ�H����{���+A��P��WV}���Y� �Y~�j}6',��s����Ʋ|;�T�^����|%>3�=I�,Bx�r���4�h�`DzR�u��Z�״;�c=�F�P�yֈeGۄ�a�qP��w?p���	+rO9���>H������bP^t�vK�l��p���v%:i�B��w����;�cw_��&�.���G��������T�4`��q2�i��OGN��������:"����@@��l� ��1`ݳ*
�q� �O�7��O�U�O���\�npa�$1�?�bH��H�9�K��� 2���c������R�-�i�t}�ì��g9<xpp��JQdAQ_5��?�U���������� �'���I��n���}�!��np��Q���?:@�HY��o�k��S�P��q'o8A�3Y��d�0m�u�h�kW���xh�@��5���J�2DTٲ�['Y$£���a@^L��6�����`p���/Q���b �q��
�" l���\���C��
�H�Ф���5�|�®b����3.Ϧ2���,�� ��2`�+z��(8�Ȓ��K� ��T��9y��������싩R9r㕧��F���s�Ֆ,��p�����ʵ���10����Y�\��ik�o
I��ɔ��k�q��[%�-H��z.wz'�0����l�b�@1ô�G$����M��9u�� 9Ja��WL��fppL&�|�����b�{��@h�õE�4;t�����#J��]�
�u�����B
8U%��jCM<�.���>�@�/��
��KK�1L�>ئPm�W�x<�:�	g�\��I4������k���t� ���k �����	��:�@��,#��mp��&{F}Gr�Ӎ렊K)r*%h��6f�����{/]'�B��$L�W����9�ǥp���4��;�~g����-��!���%Z��� �+|9~8�^·�)� ����&�!�y�:���5����z�,6ʙ�X�PZ�[���|++,�A�V������2�M���`EY��K8�I�ld��=Q��4+�"O�Ka�2�lf[L���/���f�����Q mϜi�����c$'��sM,��$ޭ\��C�+B�^�kf�d��H(��=�**�ܔ�S��%��,�B�b=���F� �k���+)a�&_�Vy�e��G)�;^��yy��pd���j�c��p�}*a�4a�yX�����4�Q�S9���G8(T�<�u 0k)�(��'9��%�F�QU�?#����j�M{�m���>��5^wzp/�����Vb���ޡ�O��o""��L��~��\|s�21B���h�*i	
��� $���@��W���	����}�B��uR�R#��Q!��H�Fю��Y1U�c���.�k�M���S��e��7;�S�P�F�|g�v�D�(�x�9�5U�����<�C�����~�<>R�`��?[����9
�Q���Rݢ�>~��T�C��t�s�ڃ�x�]�x�I�}2�6Fr�&|d��m�+�vCQ�-c��WD�b�]u��3?p0H^��3�[����O�C.�ȱ�w�'ߢ�e�j	����;����c�����~Y�1�aṮ�]�ւ�ޒM�ѣ�ʑzuW��)O��o��TOWCNԡ�>����/��,�F)���T�z����c7�b���5����@ ��<��t�_`,�aU� �r���Ajjh.��4j>�ِ�!��Ll��ef�9X�.����.� �ǴwV����6������^�H�o��{P�9��g���t��@�KvHaЎRt*�|�$��h��Uha��s/,�d�=�%�������G:���Tm-����S5Ys�oD_���*�3�)�,!e�:��&#�[:�.T�̓[J�O�A�zwri��<g����bQ p�z�cu�-�w�q(+|�X�J��Ҹ(���m����l�X;��ڐ�@�}㞔�UDd�:����ܙ>�J�����E�"x�=��J���GГh5lZ_�q�����^_A6m��P8���/�a�