��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ'���ugJ�߅j�4�4$���7��[��K~��S�#׼�8�8���!oD�KTQ(X����Y���lR���=��b�r1l4���i`�b��	���;E�;��������%X됥	��\�=�Q5'�I��Ի�,5�j}�DXo��\�r��DH�I��곧��:ҁAF�Uj����!#�/�����ѵ�DJ��h��!֭]��ی{�L{����5� Ԅ�A�9�$�&�9G{�xv��~�9����W���V��*�*G��nz�S�Rj�=���]�>���B]sg^@��䭠���#v��è�Θ�U���١O͞�0��`l�Z���c�����7��BP@�Tχ�C���+ϋ�.!l� ��"���ς���4�-�P���{�>�z�}�����g�n��Ò?b���k��P�lT{���qx�(�GWN����S�M�7bJ ���uc�ń�	��Z�����-���8|�P���.V ����G��+et�٩/X�`�c��-�~?I��A���Q;ޖ]v���'h��7��l���b(�-�y��+P	 �y�W��\�e}�0Fp;{f0(�:t�wA6`�����*[VR����2�=+{lr��>˰a��T�u���LV�"�u�������Oa����+wc߳�7�}I����ϲ6zH,�w-�_`J8����{2S
�kLK /��̗p���>�^�|���j^�~k.��7���b�M��k˗ҁ��+yo����E�6x���y��a[�s�.�=��_j��ϼ{s����ʀ�Bx�'ڽ���N!-0���%bV�\,ی�'Sĥ�t�b\N*Gl(Bd��-��v��B /Z�c�K~����u�5q�����ީ�Sz�{B�p�at�y �SQvL[�*TN��>���g�$�ݠOhj�45���^}jTׯ1+f��pLf�壆��z���=M�k�-㽁:Kͤ�d���U�g��߽�S��E��׈H��z��}�K3݀��͌�jpFv�ڿ�B��.�r����<*-�|�j�R���n�$EG�z�@�}�����������c�C�U�|4+�՞�V)RWe��Eƶ��rB����Jz?�>�:�5��x�+���gݨ^�2�#�r�������a#�$� ��}&�E�&�=ޕ��g�$�� �#!���NDe�7�k;��֓���9+���É��\��B/�Çɯ"o'�b9�@
t٣�R��9ʓX�r�I�
^~�tJ��PBDI   >�rs�W��n�d�vf�{۩�����FH�3U ��>�<��w�2p���ݺ��j�)����Y����7�G#Ydw&���a����(�۰�`���
��2e�F�ra�amPM)l���b���P�Y	֖G`�R|^���<2�t=�	k�J�dacsi�7��(W�{�#�L̝e&�|JZP��$W������U�l�;9a1�ꦏ��2��y;�"�