��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛD���L���`�')�0�V ����\����Yɣ���|�2�Y�!����3�Mo �@���V��}�&;���ar4�{~����7AvPDW�	�GG�"#�����	��L�&��*��*���xhM|1Z*�V�CF7&����<<��%����j�+��Ə`�!$��o�̦)�YPd��:���T�4�:Tsk��ܿ���y����駭Pb��c�A��m#���_�Z������֮���j+h\R��)W�s���BG!��Y�Ӡ�\�N0�J���	��b�|�����#�X1���t�&�.����Z���<#e�a��ZSF��*$R�SW��0S���􎡍������}X�	z�C��q׷U ~�w�-��E;�o����fL�A���ެ:�o�:�f�O0"�x�3/�m���ב/$u#Fro�f>���2]�G������ɦ�`��83�%�=6N�����`.'"��:�:@8�A��2�i&��J^�#m��2�3^=�p)̭Oj,��/9�MQ���v��- �h�:�T����$q!tf#���_���١�֡!�k
��J��`?X��E+d��w�t-!�4����m�G1����<W�452.�1f��\�dxW�i9�+�dv���/�]��K�Ɏ$�k�B�"f���o�d{�.�{P���s�t��p{�v]}�1�T��{��3���K]����͋���p�'���'6�r~��s�'"'��(0v!�:Z������ϵ3Ί�3va�N?��̴E���>�%�+�(���A__�]9i���or�Qbt^cvky[=��$u��Ü��,��:��IbF���ѳ��UC���l)ZZ����?S��\���_�Xs�
+I ��6h O���#B���*O��,� so�u�H
��N�->�"Y��0�Y�� -�2%g�O*?�3��gN� �g��Ю֦�JD��m���%�Q+p5n��M�lgN�[���m��G5�ؕ+���ë*֟���0�A��bVϿ��V�rw�s�*���B1U���-���z��K��,[��4D��]!>rc{S�f>auix�"�%N9�i}3�_�
�V6�"&nS,�1��"�|�hw�e�|mm�KN��މ=>�t!��0&e픉�A����ꊷ#S/2E�0zL���U*��a���9�u��Y�trK(�#��(�}E?O����鏜�](��ڝ�-,���
1�@y���Y�^0$���?yTD�� C9]�����2��#�O�:7{Updc�����d+<�R��SD���f8��D�s�ֳ�N㔁5,c���^�אb���*�z�9&d��ϰ�����В����d%�����J�5S(�'�=a�db�s�<��te�:b�9	������C�#Rz�_l�|���-V$}��C���Ow[�PeL��� ̆LB�u�#�M���F[��t�F��N�*e��+q�%�pI���k�RMb�]WXD��j�.v-J-�$��4�B��{���wnr��9d����;�x:��J~�=��JD6���p��6��$�h������1y��Cq�i���2$c��	�#l0'��_"�ͪ"f��r�ƚ�E+p����M_M���^W�e[����(dc�6��ݽ��y�zP|�i�`�X��PXR2ZvH{�O�#W��	�0��9ֿ�ė9qv?� +Q�j'/�����r��g�tR��Tw�,S�xr�Y�Gos?Y:�ά�:�*��cm�x��@ߍ�p	�����(�'�)�]�x�~��Eh�g#L��
Q^����w)�zGcR�����wbs�a��!�������c�!V񅘻fk���Җq;�Y�Үj�j�k�|�P������I��ȘH=±�$�.Q�
�.�����du�@H�Vm:�i�蚖���s�+��[�7`!W�a���.�pUf���b�vS���#R���(Io�ē��XZ�N�*�>���|��=�ʿ����`6��w@�,�pmw�*P0g��e�i�;�����|5���/������
A̐�w`<� j�0}��G��#�ʭ�H��D2IZ �K{MM[�U%t�tf5��ki�i��U{b�`h/��E�q�~ ���\kR#K��㙎&����J�>_�gm(O�<	�S]��
�����9�L�ɌVF��FyP�/��5;1���郣�b�E�6�;�kqv{����_{؜Ke�������mt���y��q,���5(P�]��/	��g�ᷕ1�w��Lz(�U�����8�s����w1˪z�!7��1�iw��j#��J(e�q�U�nKL%;O�`y�ӿO���@.�Z�rv��#�����c�7h3�Q�ӝ����u9'��I����n��!yZ�M�xQ*yм������2�X׮�ʶ�v�n%vY���:�+Ԛ�av�I��>m�z�o�^��
��K|&�����4��J�������<+���;a���l���:�5+��'��:H��>l�-�����$���}c�~2��0�~���@���<x��zΉ7���QH-���E�M�hn�����F<�|ar욖#/�q�w�͟)�!��wK�9S���e��:�\c�Gx�`� �z�Q۝�EC�	��c�S=�
��u=8�^����2���������PIKw��pJV16��˪�i���q��;l�ϴh�9R�x�$�E��O �L�4���@�(����#耨|{�����[c����yt 6�b��k��'x�ͧ��;��B�C�"���ϗ�:���LYq�F�i��t�l!�4kX�Y�Y4�R��[,Я/��L�$*?݃�=��`�((�S
ا&v*ҫ5��,�E5ݢx��^���"�ó �`�
�a���$J��O�R␠?�����5ю*���ȓ�㊫R�
��X�~����ۂ�|W��*	���H4~S��S1��`��� ���͒�ֳ{��	�����G �Ú��Bz���˨�y��˂�,�p���F�m�ċr�1n:A=	�L��QL�C�]z���	�s��IH��5�z5����������og��
c�������p�PG�uG�HM�5Ob���{����ifcw��~��Ǯ{�U,�A�dl�6a�d�fN��̾L%i��z����:��r��������n�o'Ko8�kEj􏔍��E�9�K�V� ��n��� -�K�Bp'!wɡ��j��6�����?�m�&li���6��[�џ� �+�$n��IƅC�O5�h�X6��z�t��	j�	y$0�܏�h�^&�9���||��N��#�D�&��v�����Ŭ����-l���S�V��c��"!��M�P���+-8�;N=��d�����NIP	��$����lm��;i,�e��t	��Cx��@S"��{s�Y;��׺m[�/��'�S��G��N��%r/�45 �|�[�xnx Hi.�r�hU�;~�籅5A������r��U��WLk���s�ˣV>R<�6*�?��s�����Ş�
̼�8�ì&t���X�U�	�zN� � ��R���Æ�ǻ"��&���cM�5Jx��V�[�Srۣ"|IlD�x�X����ų���!����=Ur-S$I��k�^��L�6�b?�`Y�ϖ4gE"�r��F`ϭ�%����������E2��x;[�ķI�`�	E�t�/.x��g��*��\Q`�P�� �q'1�J)H�4c{���\����r�+������v���Q���wx[��6}l�t�ض2��3x��<=Hi�P 8�� ���#F����l!A9��ii��(N�3����3C��y� w*q���vd�qcp��&�hNMJ Fns�Ũ�*�ѕ�)���W_�K0��|� ���\��#;Vm@�Ć�ފ�B��L�F����oNdXƎ��e��i�E�e
Vu���q��s����9g��,�()EL������ef	o��V�K�dEN�&�a$�f�NI�K��H�7�F�.�~>7�#��M�鼉L��5f��@�\x��럜� ��u"��zx�s!,� �&:�5L2FI}k���3,��y�1�	���}{��a���aG��%bb�FA��Z�\�\����L�&����D�[�x! g:st��]7W���ѧI����T��������1?q�KsW��(l"*E�F�A���}cPiwQ��GЯ�q �]l��v��n��vA�P���)�ym��3�hw?��) �ŋ�t�7��ݞ5�'���c1��󪧧qx)�)��xrAh�E�Ͷ�Ho_yRl��͝<2��-��G]�r�Aӌ��,�q���E�P�O��ʳ��NTH�z��/~��+�ᤞ7�9�B�z �Q�Ц(����q��j�ˬv��oi�pg�GP"�ܦ�nr�P{�J]���u��~񚃕�7�j�kS��<-1����_�d/&!6�[D�-��	z�FGp���=#��7-B�?�vx���(���dP+5�/�"�y�%)��3�����FfP1�k��Te�Z�	�[if��l|�>����K�!���\B6a�<$��5��tP��?%U���V=�QU��A뻰{2���/!'�P9W��ف��H0�O�4�2�{轅�J�ľ��Hv�y������(|��#�5a.;}/~B,��.���O'�>����;T�)��Bl��Ϙ��,�{��L�EKK���}�R�GL��v�VQ��wGyy�\9nD���6H�����U�%E��]��I����W�m�%�I�hGd���4���SI�u�N~�֚�?w-q%A�Q��r� ̧>K�N8��sѵ'�;l�I<��S�t���=�l`��b����Ӥ4�w@�x�\���Q�:�=��|k���%�
ǳ�8�h��8��e~߽> ��z�>�(��F*�c�4'cyp�������
�]�XJ2�?A@��/Kp���+|�T�Hl���̩Ŏ�q��9l��j�	+�"���pl���ko�5,�j��@w�׏[g����# ]�1X�
�B�Si�W��5旑��z�]A����P��U��7Dq��W@��<���B�k��0�G�a{.sJ+*<��i ���$��.?3��i�֌�z���f`��_Z�ͧl���D|n��	R�Us_w8�j��-:Ҫ��#�Ԙ�w�+(��;��3�����3�-z"��Ĺyk��8-��>�)т:��M>;��{��Û�J��e���}\�C��ٯ��Xi� ��ZqG>pl⑻�
���E@
���6&���crЃזpbr}?�/�W@�!k?��ܦ�ՠ�;~ӏ�'����=-�_��"9��NF\���o|O�b3T�sc�����y��%�XG�t�Mxܫ�`�'�8��}V�s��?B�U�y��VY&mڇ�A��G�����%�Ba",sP�y�gR�W!�y-R�t���� Y3�ǟ9G�9�D��Dp�
j�Gio�=�aR1�h���w����t���V.Ԥ<x(��?��e��;�}�7gҶ�2�۽�L�4r��@�E T��Ţ6��,���O���1`�&�U�a�i*�?�� �|���
�v�e�w��E�)Ls��~��fx�s�>W8+���5����%�tnJ�$�`����՘�;��'Nh�俀��!�aw�<(G),�kx@l�~v�����w�ף�'�l)��G���W{o�w��fR�{1熄�/��8�
�T��Q�/:��ΰ���1�6x�S5a����'��b�Gztn���h��Ɠ	|�ţ�d�&Ӣ�HЄ��#�(F�=��7B�f-%g�� -�����7N{�WCJ؎3�����JW�ʒ�1m� _U���)�������m%��c����"���P��@+P��=6�Փ�~������[�w�	�f_��{�񗺮z�F��M��+�vm���I�ݏ�����:@��H�ry��PxPL#���|}]ƛ��e�n[�ұP���-3�Z�b k5���� ��:�eY<��n�P��X�#�P��WY5K�V���đ{�{�L�liY�@S;{�A��3N�zg9!Žϫ��3cbf��Ja�5%�� �"�|Q�5td�g�ʙ~z��(�i0au��[y��^� �:���h�$���!�_�Rݫ�blB|�R�p��MS���#{�����y)��5�I���yi����������&��M	��s�i�%s>@�x��t���F�o���S�4Vi8�g	���S�p7�����)�ԧYHb�C
Eϱ����'�"!��r������B9����յ;MG�\įG��Ԕ�j��ǒd&0������uڠaK�����v\O�U/�V#�OR�E�T�!O�;��㌬|p�Ժ��0�>QE��r��A	�K���о�NO�n��7�3�� A$<�b��!��;���1֡|%���k��^N��|�<�}��:U
IV�7giL5>��度&]�x�z���%UI^��+@�!oT���"�}{�m�������FA�_�����ɖ�h]�Ğc���19&b������kֺ��fG��W�o<+;m�(�oh�D�Ê���}hY�{q����,I֙�Fl�>y)��|Fyk�"F8�YCR��GN�6!�'*̑e�-Nt߹��6W�/��h�2M�=.�������h���/���Ѱ��Ne�M?¾��+ݎ�~,0YK]���E׌GW���|�K�U/a����\���VF�A���FY���{8	ݠۀ4����"uX#�ߺ��T�\���k�}��Vmdo1��� �e�͙,�����8U���1|�o����O|$;� ,�0^�/�q�i��V�cj@c�pMS�HN�R�>�'�ܖns�s~�+��j��k�Wt�
>Z����&���!�^� ��S߆e�)y���P3��:��:��5�H�ᤤ#��6����~bF8K����Ѕ�*�*+��a��q�����2��Y����%�L��=�;��&�rq�ĝ��*���J�0��|Y�&�.Mmx�i��=��)�b��I�)v��m�y���&{W�y�yq�	��޷Nt����,�FXvyfk�V�a�|Qk�sy�2c�~M*ݬ&��_uڙ����@�\r�T�c�1a��(�>�!cA�4��ɾCD��@b�s��;d�U�fQ�
ۿ��r���eo�<�6�ʝ�5B���ڪ��Y���\Y��K��kv�aDo����ˌ�� �+����n �)�I��ŕt�f��𛉈d9N�Y5Z�٘n��L�KqOx~�;ũr��h�̓���;�nM�\gusC�wԈf�m��I�"s0�6d��7�֒ #�謞�ΧBl"�9��<���`��w}����7��:3�y��Ѱ�w��-'��u6�dr� ��&-��m}_�3+�.�'���TJ_�����7��gS�c��u�@	����l{�����u{W�[����P��o�zZZ�ĥi�۔�A:d�雮r�O���#R��*�6n��l����=���Lr�aժ��w�6?��Q��!��wL�+�i+f�{M���E�9F�ua�ݔ��|���)�ՎuP.֞��g�5,Q*�.��B�vO#0'����ϝ���)�4�G�sn��J����:S�w�OF:�Q0�v�;���FU}��V|���c�L�5����k+X���&;���7q��:& :��k��P�@�ܻ����|�c�~�t������R�8y�Y�Q��+҃C�����*b��)R���y����k歟�nA�& *D��K\���z�<��ҜN�Ow�����#t�ݹѧ��j���������H�[���[��l#�jr瞵j ���F���3=�^��T)Ň�~}�X��O:1]*`n��+��D���R51��-rP|}{C&� �x���3���N�J/��^��t�	J���7���K$<�9xG�R&0�5��i���������x��qT��Gj�ݤ�+j?��l�<f�@���7���7K�pbb|<�x_�/��?��%�KdR�Ⱦ�~�5t��vJdC� .�:KG�;g��̹1�I���e[��q��e�$w����TXk:BD(�|H�%�n��d1�`,�٠����}�bXʝ�	��\��w�<���(��w�z_��n�b�-��B|�Ծg�3��C��-�s�Kj��7XNH�����D�SY� g��qyT�Fn�H�|�.jY���Sʿ��Yxn�<B/�S_�>��@u<�g��2d��H�����,�ֹ�,����3P�n�K'����Q�!��'��N2�g�������]S���u��\��"�cV�FO� �5������|�]�5�m�ବԟd0�ğ
 ��#��n�8pL)�d?H�G���?f�q�e5eb�*i�+���F-5��(}���V��S���b�"��I(�9��lF^��"�!F�U��ܦ���iF3������t�\�a?�ނDCV��㱓c� ��1	�m��~�b�/�}�����['��K@G#=�J���Q�R���ѥx&k�1]��>&t�n�lZz�;����H�Aэ�ˮ_��7\m�P����'"���{k��� ����w��#�����*�j���X+�Յ�)���!��fu�CX��<�l�F
g��utZ������Al�,��֊tnA`p�3��b�Xθ�H)4.�$�����L2!�n��Y�L;�����e�$�������)�])a^гى��!�h�Y��/M/チ��l�=f6�hY�����F-�vjؔ��i�^��F�����j�	$]����U��@w��f=��^T˷$��{����	��
M.�bqxL�&
��9��®���M�
S^�$ɜ�"X���\��,��X�:�W~���d�c�tv�-�I̍��SeǹQH�@!��IPϗ�����"gaL���R*��J#�l��/��Ɖ�u��LT�� (��FB�ޅ�I3y��"��ar�[�|�K�cj<�������hkl;j�@15��	��/o���'=�6Ҹ��u軚P=+8j� ��Xtx�3,����ԏ��eO���Ld��>M+��	��R^��)����Jp��*�77ޅ%#Ehf��c��6�JM[��T8���R�}�hk�:���g>̺�F��I�@�#���RVV�6P�8��p��]�YN���^��6�{�5u�Qv��䍔�����C���I�k<��� �� �
�C]VKK/V҄���/g3�XŪ"%"g��X��ݛ˰$o咞�:������2��.�T┇WE�=g���S$l��+�uH\�P���[��(��F�t��U���kr�eH�x�ۭR��Y0�/���T��z������<�,sEƦ����8����2v�E�C˳�F���"���Z^�k����F�56�"p.�N�9�;�r���PsAM�9�Ӊ��§��E�0�� I�t�:`���	4������i����i:=n�P;	����*�e����`"獪�	�B)a�q#]R���)�*KA��O��rV:�_Ѥ�nƵ�E4.~7Sns|-7=M��k���R7�+Mst������X�YC�*�}�]���TOae������\�l*��i��V'uk��<�X���z�({�DS���/y��.J���>�	��_�z3�+�U�8[��m��pWgy�-Ehfh��J�U�&�EſE�G�u5��1���S��4���	��������&�Ly][���-��S&7zB>�g\0���c��K���XCy2|�w��j�A����ŀ��+rm�*��,(���&?��3�ڼ�-r`�׃�Y������m���fFn��!���D!a�U=�!nT�~A��\V`k��}�L��������&�@�/���EZO��O����f	�ВT�h@�x�L�-O$� ����z�5ٙ���'#�c��mm��$IU��5��7R���k�\*��*?�g����Bq������P���f�\Γ�q�K:>�&�\����|�
���j�Y5�e�4ifT���TXc�Z����������h� n!ȥ/��Si��ρ���º�ђ�ǅ���~�6
V����g���L�à�f�֧c<�z=A��W���_�>i),��䦇U������NB�辟}N��Dy�H������<lU�=���=/`����0Ph�Akp��|;
d�������7�I3��-n�Sך������W�w�y���r�0��m�?�S9x��ߟ������H��F^��-a+����^��1�d]�y(|R̯a7�w�����ܥ%�.ؐ���X4�^C#Z�����V�G�	����8���=5Sԥ�x�͐w	��`�i�?Fw9L^�ڛ�p���j�tD�%��y���/l���U�n	�T,Y:}�����7�~��B�\\Ѯ9Q.��)���o�_�E}�_38��W�8�Y�-IIz��|Q��[���C�D���������H؉R�
�|���?�{6.2�՗��y��&�gnm3e=)��_� �C�wy�kZ�nڧ�2�}Sr��@ջ��'P2��DFY��k���ˬ��\J� �LM�5W�<���6����)����W� s�k'{���m%�TH��T�|A���kH���gl����.�Ɵ��ba���I��
�:L���<�9�w�I݇w����g���,� T�
?���i��D��ٞbB1�4�D��4?���>��9u��H�Zi.�W���[ܷ!A��Կ�p�պp%ډ3#;�y{��8�k{:�>GIƞD81�A�����h=���]��	��~<��m�B�.н�ӥ �bp��g�`ĺ�%��Ah���������#X�6�eE��K�$�)JZ�'R����4����H�'W�(�m�~:��-w���ׄ��5��&�Q>p�I�bB~�]V���䢳���8 ~WG
T��M�1�Y��.Q�~�·]��L��,��F�R�]+i��=��rA0�s��յ神!e V��񆏴���z`��D:۹'�E�kK��\\�O�q�jM U_��֤(w���O�r-�t-�2
�4+�ߕ���%�7�쳷��!� "N��Vh�!3���Dװ4���C�2�������W�m1>�M��y�6��Ă�AG���q�	m8�1c��G2B�=�_���"�)᩼6b~7����������LX��~�����'Қ"gq����G��̕c���{�ݱ��֎j�ہy��J��ǣyݾ↟���8�v7�4^W��SI�F�Z;���:@��֯~�3Қ�6L*��!�=Lt�mD?��zޡ*8�����5!�����t'�P�#�Hb�[�d����2�>W�[����K�)5����Q�dl^RJb	��[!��@�Iz?�O��0��_y��$f5^C�C��6.��(���s�5j{�Y�o���[��@Qc��2D�Ӊ�����{�_F�T�����d�W�d���s�\'[�6O�[ U�U���t�Ci�����o�?U�����Ǣ�|�)�<uiu3�����H\�|�EkS8��UyRˍ�����|Q�t/e=���j�"��o��n+��FD�B:�ܠ�m�y�ْ���f<Ǵ��S��fM���aE[�YE���NDx��E����~�Z��3�wݗ��,x�[C5n29y�&/7�n�.����Xr�1�����ml��
��P��Z��Ei��*3����n�+���3hDW��7`x�h�c��H�i�>��T���#�yUS*UI��<F0�m�oB8j�H�̟��XW9����R�����!�XUr*V<�p|Vj�KB���7TwQ�fΑ)�v 9���iD�Gu=�/e7~3(�7���]�,����P�?-=l�#C��(��$�ϖ��H%�[ՍB�(��y�$�j�����Jd�H;#�"�܏}��ٗ�ci.L�	�3/����_$���l�܉m�
��Qh%F�6pz6"�@cPkJڗ���Ul��m�Ţ�Jo��3��K
�Ĉ��q%EݬS�A�#��^���p�o#�����s)�8��:z��0�ڟ�Of�'E/�T�c9���i�RYڇ,Z0d�_,�f��뚚t�3�����#�>��f�*���{h�`�4���;�%[P������_��Ne��T����[�"���2�
�C����� ��t��뚠4c;�r�W(�T��;�ߐ�T�W ���G����D���Z<;6��7�L�����OОL� �&gj$Q~�*�R*6�i�^�_׺oʽo���SMq	�� #���#d7ޒ�\d�ta!e�W�j�<�j�(�x�o1,Z��yL�R;�M�Ă�а���C�mlGb�:�'�`7}ϩ�i>����U�5�̨rp >��B+���� ���`q�������5�����dO����6���^+GAϚ�w]ӳ�L�-���M�I���I!�R�[��|6 ��G�o�)��,�/t����v��w淞-$��YW�u��p?��6��[%��y�`ד@LZo���K(�O~hp�-�A9wZ�_����F�?����ۭ������٧�mǂ��{L�܂�u�Z�憧������{WK��A[����*��R��E�f�<�{2�۞c�*�l��Ţ�i	��'��z;?���U��!�˟>En'�	��7e��������BlRât#l	H�ۡ��@���k�R8��{Z��.N�{�F�Z��W5��4�|�"��Z��b]m�Zr՗�Uʡ28��³�?n�a���R������ǲ���:��/��n���y/?�j��� ��9�p��sd�[��liv�1ũa6�Z��0����9���A0Tc����l��>T�Dy���٥4r ^�p&��^�\G�j
�l��\]h�m'��ltF���0+�y^��O��DH J��Ar8�~�Qjur�u,
�b���Id/�G��h���Q����o�mZJc�0��[%TwmqH��O,�1��5�0���2(�X��c(R,��b�*�ur�#��s����N��v�J��`3jѫ�_��F��ǬR���y|:���ϰ�e��I�J��\��x�!����X`�d/���]��O��rL���7YX�e�V��@���"��;��Yzv��7L^ђy�u����!}+`� �x�\��?�X:g٩�Z�w� �:���TV�C��J��0����G��������?B���J+���A� tK�BR�V�NF�k��h
� s
�&Va��qnk���L!D-�����`�y:���+>��Y��o߿�L#"=N�-������?;s��zL�'\���x.w�6��b�I�2` ^�C,�Ѫ�jrq�U~TiW"��@����S�r}@���@��,���л�p-j��k)���3=S�ߞ���G�����q�����̠UY��̉d��-�s��K[�$뭭�׃	z0��s:f�-'��v��N�69B�a�z�ee��F3��!�_�Ҿj���Oπ/n-k����ۣ�6�~��㄄�;!7|�_ �b�U�����#t*�k�;�'�A��B��F���I���5D|;�M�wjѣ?�Fa�u�Pwk[{�9��1ޓ�y�(KwӅ����������)����������f�]�,���#0�bZ�-+�%)�t��R5�&>%�`�AW��'���0ɐ�׼�C�DO�n=S��w��N��L��5��=� 6�y���$����Zhk�e*��E��;8g"��i��gy������:�o^�)�(�7gύp�{���Eҏэ}�>��r��q�}Xa��rh}B�k�ޝJ�_YW$�w�,�b�;�~�b���gY�/�����M(7�^1G�k�@�5��o���w:GO����o��p3BI���f�1�ʍ;�yda(����!H�8��̇��e>���W��!`����b%��ޞ�kl�S�|�?����U��a XN��h 䓮�o+Nn�=�Ԁ��:Ye]n|�5()&D��ʭ���38;`����t��
ͨjt3�	�	��N?�^_�؝�?��o�"n��G�f��;�t���3��1K�c~�~���޷�q����q�N������ղ��(a�t�c3����A��߼,:�8��x3ӊ��(dȑ�pu�e΅��O*#�l����^sG�~����$�t ��b�I�?���q���Y������Ts�z�Ïc�Y���� 8��ȪnHB��G������<.��%6P¸h�Gz��%(c鿎�<�� �N�P��^3̵$�eؚ~!��&T�옝�Ï��6�:�9ļ9�UI�Z�Kʱ2Jo�Ȋ48�71�����r��uyC+$�����}�RW@�q��l�Q�Y�Y߲ ��)�Bb�	c�E��ʝ�W���ګ��	��gZ�kR�G��J>�"���n�ť� �C���Q�(y-m��S�:-9��n�	I�&���s����ŒA@�����.��FI��ͅn�
���߃#��ٻtc� ��k�8����g�W�U;�tN�O��8�;�ɧڤt}c�
~%k��!£ׄ����� ��J鑸�O.N�Mg��v�Yx�'�K���r���~�,�Eb�]�e�_3;�l�oL3���,4�w�-l������{\���r|�}��Fԅ��U��M}T[JW���z2�b�7���8�Y}:�9Bv9��tv&��ݹܬ�k]�+cA#nGU����9��
���o��in~�b��k<
�"i*q�A9����X>q��B:��Л�GH��a$)m��|Qw.^��RxΙ�#ժ��"��*2-!����]ӌ�d����I'�vK5�r�m;6J�A���w�:n�P��P�+���X��2�i�y�&�I1u4'u>������t�?�MS����T�Tž��uK�ȬJ�=K"�>>G�J��[�x$.9�[:�(��^�;�e#i�8��*1H�R�����6l�Cp��]�z�8_���i��R�Xvv��vˀ����&���E��9�J�1�ļ����d��?cÃ�6"����˦؛��1�ub����W��+���;��<�aБ�[hS:+�|�P�F�Q>��Ͼ$X��"�<^��on��:��Zgd���Dǡ�Y�%D��@��Ƌ�"��:��^��˷��eR����>͙\�h	%�>��c=Ծ�������a
r�֏e֑(y����F���"��"I��t8��;���T�����(H��Չ_��y Ȫ�\Y^�6%p�&�(@���(�f)|���Ŏf�f#[]�@[$,i��Q*,z���U2�pm
�U��l����3z-H��jTc6�A�;�VZ�|�ʣ^��v+J��=�	�粗Y�d1\�{� k ͜z���Iqo�9n�0,v��썎wȬ���B�nM�������kKs�q�u&'��F�%U��{	���7v����~�\�<��Sɭ���p���9^
qŭ%ﮫ�푦n����SF��K�eđӋ�3V�i�<)!��
��k����K�r|�Z��p;g��g�V�Ѯ����ϕI�(���d�a�&ZD���	%	��Q�3��ta�Eu�+�M���6�r���y��Jt[�^~~L�>�iE�x~QM�B@�L�2�&L�C�8OwL�&��Ӯ�W��zc7�Y�{�A��o���v>ic��3ȵi��(���Qh?b�v���yPCmm��!��^�������w��q�@:'P�]��$��x� ���a��� �Mc&��f�z�cܲS�ur���Sb,x�38%�q�On.����b���M���,��b�����|`���5�:�V��ͮ���XU��z�q�"O(��v����8�z�r��^^T�����SO�S��T�ox����!i�+�i�<�c�?�]��\���I'7�B��WJdQe?� .�'e.�,&	'�4��Wul��bV�C�l�Nϥ<|����ZS�D�W9�a`�����v��DxG��W��p����pF����P�����a��VC�PBi^.G�S����J��O�d.޸���E�Be��S�Ul�	�ao|;_�}V���$�b46b���f	��y�e����|�Ҍ6 )V>_�(��X}���Fp���*��/	O�{��4�əw�'>E��ѵ��1d`�^0�a�����/�1a~8�)��`�oBa%Ow�t)�` �7�hRV�e��G�g$�{�4�yם�����*��Ϗ8W���5��_�GD�Ǣ��=O�j!�����j9�@u��weצb��Y<w���۱(N�1�T�bG��G�7ј���G�����4o��U�~��+*ҿ)0��T�<-bN���;�kx����)Xi����x�]F��:�W������/��%��(������q0'�A�A��⠙��f�O���/\`9�� &� �=aC��GjE~�SVW4�$ĤJ><����%�%ϛ�{Ρ�asD̚�`m������d���)���/���?��@\(\��.0ز(}��U�MH��Pr?�`�ܝ�dw�y����YC��q���Kf�����9�~u
��ŗ�w�1�{�q��SY���\�Q7ȋb*kFi]��欢�J)�H�ws�'�}?�&���`,������[�$�<q�����V$(ȩ���i�Op�j�h��A^Mk����̡��S��O�{�؈�[S�:��4��2 ˥^����G�tí|f����:�pC��}��W|]L m�q@-�D�M��~"�f%sէփ挝0 �:��8��"�u�Q�6%A��7S���`maS��S���0�A;�ip������яĴ�](��3��~m��vx����nMT9�rG���:Y��澔F0��%[b�ݛrq%-����s0e�:�@��Bl�'#,�&.^�&���\͕�[0ȝ����c����m�u`k�P�@+��s�V�adυb�^;Zr��2xqe7I��V�U�$@hi�H$��?�����2��hO�3�q�օ��;sf�Tq$�~M�Ʋ��n]��"Κ� ��hZJQ��S`�ҏOA&���gG[�u�_�v�9�E;K¢$�U�Ec�Z��UB3~�4�h��	Ɂ_x��xX�̚H�%�:1d��)��[
,��Z$O��I]]��Zi���WQ3l�կ�^��أxY��63���A����R3���l+\��E��av�z%�f�[�:AeVD��SpqaJ�䭟Y�=�(�b9�/��^hn;M��7vVb�� �d棙�.�ؐgf3,�X�R�������=��,��H�k �Q�h�QQa�\<-�"i=�Z�f�~=@H4��M���m�e}IJ@��ˣl��B���0��<A;\�DR�2�u0�~��H�W��y����S3�e���(�ʙ�����Ʌ3���?>�7�&1�橣�*�RH���+H2�&!]:�lZh��
%-�v��Y)��"�<��G�4� C� 4pb�v5�~�g)�+k�w�24_�A��׀�{.>�¼_67-��U8-�6^�C��Z���W��$>5L>O~�?Ѷ�Q�����aF	�Hz�xK�E
���dN?P~f��yg��b���3u�>J��AL�b`�;�k�k���pDѾ�7#�<��c���{��ja7y�BѬ�?̋�\�=�M�ԙ�Uv�"gf���;[���e��{�������ҏ3�J��{~]{�~0��i�� .�Ϯ���{Hp�o�k%�����[���݊!EA�FJ=~6��-�����0�/AL���@�l����1]�K�GDTVsXR�����q����*K'�Xd��SO��H]���>��hmԧ���R	��F�+�_Fd2��dL��B]M��*�Z�i�<��I��8�-����t�������h�Ȳ�\Y);jt�����B,�����R{�6e!*�p��sY!>NV�0�b7�*n�yDB=�T�����מ���/C}����%�#�u��4α�:�+W�-�U8q��-�ʁ�G_��?�ä���Ƶ�X_�0����b�Ѓ������a{п�^�l	�C��}K<����'�F�?�l`w����՚����-f����u�A�Bqv�ҧ֦zHkn
��;𿤃���m8SQ5)ic��e�&FI����i6�20x��t���޲��r��B��r�t=����
��^�x2��Kl	�r}����[}W��pd\�L��)Z� n����Ha�z��c���:�ТͯA,$J�:�R_7>�(^b|ɖ;L� !|1q�B���Cl*!�Z�#���%�)�v{��:����$�;��b�)��f.��Wb!���p��*�4D�iY����i���T�X��kW����;�T�@<'��4IU��N��*mh�j�������cq�μd��D��+s�V�d�P�J*8���W?%$�y���Lo��{kX�������0 39,�8cm��B��rN�V�%L(	$����J� qgUJ��!�X�(L�R�'|���ht�圧��v��#�}�N���#��~�`�\ڦ^�G�gG��%h8��o�_J�r��x��%`A���T�*�2�6e�IL�@m��4X�sh���D<�:��LW����\�S�� w#�?W�X��h^����,xx�A����G͋I��`Ţ~��}��*>;�I�n�� �%�f����w��T`��l�%�0�!-�7�l����2��03wz�x��W2�]�g�<| ���*���|�wˆ!;���{A~\��0���U.���ð�B�����S��KZ Z�������������� �Jh�e2r�Eߜ�r8;'G�e/1N��]\��1��S�ʕ���V����b7�y�p��\0�RЁ3��Ms`��@���ꃫ��U��U��x��� ����%�����\忼w��ѫcN �9 �',%�[l��hl`����	֏��l����_ͤ�d����mj�Pe\^�t7�5v���Z�v��}�2�u�*��dq��r�H�&�n�Ơ�Hm!����W]�p%��˩LW�E� {&��Z�݇�%�J�mH��waa&�θ~^EY۪�À�mM�U�sºfL�٢�Q.����MpSΦ�&☃�����J� q���P>)��TM�NW8r��K�黎M���` �*'k�H�W�!	t�l}��ž�{i��SB���=E���̝���A|IG�qу��h���T��nx�����a@��'���W�D0�S)V��n"��%~c%����9%��"��q��;5!B�6&��/��t~2N�ϣT�^*�Ys�{��O��E�-�`��(�G��sxq� bBQ����x�!�6[� ;�mD���#��P��A�LM)\���B�)sV9�"�fm�����Ii�4�Y Nb�b��$��
ԩ�F�1���c�vw���u@z�&�?����4����zZC�d=5?'E�ޛC#{�4)���� @u�ƍ��޻��wy�û/���-�&F��;ſ���Z=�4�`�s�>."���?�6�`��,9���lD^�+���[� �Zv6�S�\
�b��i��_Y\�Yy�Y�"S'
���
2Z���5_�c�8���J2`����/���_a	=.� G#�������1(�� ��c��$�-�~e;��ޓ�e�J��q(��r�ѐ6���
2��� K��q��T[r�7����5?��KK1;� ��Y�k�����e ��,�Љ~�/�Q[�&�S�U%-}k��+���Ƒ�C���ԙ`eg0u�t0���Ó�Kr�)V�)�X�i�S�E\l	�#Ա�j�()���GĶ�te�t���2?��Y�J�!��{�y�KR�ڽ9�ڔt��by��\1{�2��jJ����'� 7,���p ~����+?Ke�'�4��9"��D7��=+�`!�EQ�u?"�,����֠�UH�3�.s�\���ZlT6���\�ld��,�����^z��{՗����ę�2$�E�^!�s�N����"�[�6�i�����z����%K����$=(,+(��rHX ����w+�ϻ_=\�|���&n7$o�c")��D/5��0�ƏK�[(�t)�~�DX[$�@���*�)c�W(�O7��Ө\�p�JqUL��]y��E�
N�u;���F٬�	+"{`DG���Q��|oS_z }�&g��5����D��$5Ud�9DN�)�f���:L#O"�s���g�-{e��j�x��>����9rj�k�-؉�͐uqG�X���ZC��y��0B�z���b��}����T�N����*C��u1-�o]�����N��іֻ���y��M��
���K����?�u�?%���}���+�9��z��ƞ?�l������� ���ƃ�3�Z��Nnhd�"�t����_%������c}3$�s+���W�3� �c%�����ϑ�o�:���;����;�?�C�aG^u���& ���,UH�r��*��������L�k�u�ev�:�sV�-�����K�'P���ܖx&��qa������o|�<��N�`w�ӡ��$��֕Tja�D��@�����ѻA���n�����Y�*7%�u���ʔ[/�ш�\[����^	���"&��ɟ����q��5O:��D73��!p�1o.U��`z�)&v#t'樵X�1���b�|����Џ0��n�c�F�<�D��22J@�KG��g{��U�X��q�O*���ho@Zvx`rH�By��m6�͖���Y��OP�����Ĩ`����/��B��Ij]n'!@w�R�Ԣ�$4Bj֕j�}��[���gǩ�����ԫ'��q���@�����}��+^D~f�K� ���N����]�
hP"��P�9:�_���B�����L��IR��d�MY�U�+�oEQ���K��MjYo�"�u���n�������ɚ���,H��>#kGȯ:�(����u��X:E��G�۹��bP�5�s�Ӌ̥H+�7,K��Д�R����G���ܪW�Qvu��9���C��T�4!�ç��q{��C�O�)���O4!F���;��~�S%��/���-�lYw��ƭ��v�S!J�� �h��A�_hV��l��vLO�]��"K��7�1�i䘚e_)����f��*���l� J�ov� ���g�ۿ�|��{��Z�=�TY��8Q1s6�t��P�d�(�U;�A�
3���)�w���7W�`�R�T܂Oy���>�oaM���
S���U-�s�%�7Gr��DPR�B��_��H��X��8�M����E����&�JAZ��X��aWg"#n>�߮%0�%��
?*ΟU1-NO��s^��Y�(�r��{��b:��^:!�>[8����;�Kա�L�n�b}�����C��
�^�b6�[�����ֈ�ΐ/�$ØH�[�Ks!�D����-�zD6�6��9L�3VϞ���^���Ѧ4�y��!���\�-:l߇iHSZ��k��Rָ�ꌠ-�%C*V-Y�Ьy>�y�&h��`I��sK�|1��]X"����ŝ� -�U��u��i��l��u���?S��9t��Ũf���=Hs�\bc��[��r����b�?�rJ2Y�:U ���c��̛{�Qɮ�A@B?T�>q-:<b>6�9�(���e|b&�41T�<�}ԱQ���Z9W!Ĭd���� ����g���;��ZF��HB����ei��&T�P5T&d�G��P	�ț���=.EH*A�{>|���.�\�+�g��?n��eYVЫN���3Sj�o�m�T4��c�}������!9�-�G�8�
�����P*�*1�'#]Y�w��\T�Yev������B�3�o���J�(o�~��(��D�Iq�
���g"pA�r^ 㢉��"�F��9����ᤠ˒xoGΊ�r�l0�X|�2bbC���
Z�=��[r-bW$�
d�J�K��6.O�P\�NeЋ���*��&�����f�k�\���; z�T*.��ȉ+�&��Lg�H��~���f&l玐C��Fh�VK1Tx���o�> �5�x20**�,�e/@�%`Ѷ��T��f5�*�ȍ�NE H )c�_�#����y�╫�4s�~=��_W����2;E]J��D�e���k1,Mq��FZ�NCs=}Mx�@}��`Ԯ��@.4Uk<�?ͧ���X�t���7���ج�&���e�pU^��Q�#�<��<__�e�=�Ѭ�����9=R��]��*M|h���O����66�������b��������&q>6���Xu�:"�Xc� �V�T��C�a{�{��̸Ά�5T܈���;��16ٝ��q�.�FD	7V�r�� 8ѿ�2�-�w2��.�����.}ٲ}5�l7.)�H��q�D����c1�ŧ�k��_v/o�O�h��.��-m��[�׉x�_��6X1�iYsAJ�O�iy�`�d7�x��Y�)
���y�;v��7A]����'�z�Q�&i��>B
��!Hn|3Q�o)��)kУ	��Ռ��@�-��i��T�.���������~��ܡ����J���&��OK�����6�O��,rHv�nN���-��O}�xz�l���Va��X8YV�3U��f#�N%	��Y�V7�pk��(�����ƥub�N+�����Y�V�w�n�SF���<��߯m���,�f�S�k	�����Y�����S�,N
6���o7Z����v�*ka��N,Sڶ��-�C�v1)��ǴN7����]�pd�1����c,�3D�9���[L�8CO����h_7����)P�و����d�pVM ��ok|x}T�Z���A�(�V� �nV�^�+�ʷ=�&�Ze�"\��q�����F>��_������#hRx��b���"����0$]����*���1\�Klƥ�("KHO�c�BA�o�x����m�z���q�>��*R���t���1(�iA�L�;�*�|�d����:�Y��3�Gg:k��)�=�Q�Zx�&#�J#r�a�O_�����?�0N����O�=hLI2��%u��L8�~�A�L��=����uU����L�sW���CJy3�f�e��},5�d����V�l��q�����WI+�L��7�O*�ŏ�q@��b=0�%y��OM�~px�����l�8��v8}<I���Y�/�ga�h������� �?�����S�xZ�l��X�c�e$��&^��g�����,F7��;W�|1�f��ng�5��P� z}�#XO�YR���`bn �RŸ/5�u��]�Hwz��cNG�wF,%o�8�%�`�(G+��VR�Cuk��>a5ۺ���D¤�Q-PfP8�NsN� =N���=��9�_�O]�?�ї}�0,����N0�,��M;�lD~�jK���T�A���E���'���r��I�J�9@�vMz�F"�4p��U�n���x�gS�Aǣ@c�@ p�Ea�� ���&��r�aBT��|�(7s`�wC
[��TF�w��-a��V"J��k{�/<o��E��'U?Op��o�'�fg|���e�K�����^�]9JĿ̒�I�ZX9��e��)ǯk^٘�&�B�!��?�"�y��X;��_y�,��K釣��|���d?��
�4� �X��j�2�"���t
B���y{_]��y�O�jLl�&��	��3�$��De�}���M����v?0M���q(��_�5];����m���a��ޘ3����V�����H��bK=��5	g��(��Y��q���R���!z�>�mf�a���V��+W�|�{ҳ��	t�ϿkU�˃� 3PT��LV)˯�-+nn	p���XS���_���t#�eY)��1[6�Ŝ&����P����X���4��|y��)�ʄ	w�K����Q��QA����p˷�O�g{��x:%�����d�@2Y��k�c��|y���W�%�̄��J�nGLx��UQ�	�0�K{���[�`VL�q���t�,�~�B0E��1���%b��ʖ�ސ�%���~@�5j�l^��lj@���c��P���xچ���[��������� ��7AW]���IU7?�0}�.�L$`��H��O&C�ROob6�,��D-W��M(��+�$h���Y5�3'
�]� �t�g8��0�\>�[AR,:F[�B�0O����\�#^!�v(��n��԰�ޫ��ɮY�~����7�}Y=Y?��(%��Xc�[[��E� ߦF꟬z>�������m�l��O����45���s��7�	�F8c�-)��Tg�����]�R"��A���N>���;x����*�����:8�[gjQ.�� 2*�]V󣬤�9��k�l�?�Bw�iZ������>\@DB����FWn�78�5� ��E�HŒ�����!�s"�sq�Y�K[���7Xt�চ+8���t���$ɎŰ���/g��	�)"A�{�h�Ѯ/x|�o��~��LpƝӊ�J��E�T�����A�8f>V7/��d������4��x�臑���w�����+(9����<)�p����0β��K#�XX��l�|+O�F�^�U�Ñ�X�S}*�Vm�����tϺ~S�6_�_*�{��K��򂰢W�l��i\������6��^�i��:cねݡr؆Ԕ1� #� �]ξ��d�Fg���⍫�:k�q��(��:�V���S]��R��Ů�3?�9@;�bN���,n?D���嵑@�~ Jݴ��c6-&��=�򻘷C�R�f��W�&7��l����b�1�j���lv纣r���'Q
�A�\��  �^Ы�Gy�Q�)K�et�����0Q�`耻�����-��B��ftg˃6���%C�.Ě0�4n���#�(_~��Dp�����d��5�Am��V{�A׮��g�m�! ��hTA:����T&5���ھ�}�WQgEC����36$XN��E&���ط��?Υ�.z�Tp�ulېD�FX�mgJ���9g�h��n��z��^�ZT�e����NԹJ�[�gI��s�aq<I�L�|�/n(�7�8��9B��]�`׵-d����_�'��3��y�_���N<$����5�]k��n���,��A5�&A����!KN�]�Z��^�|���A�H����NthF�(�(3�V��:�8n���tya�k�LCc7�@��;��O�� :R=l��.���%�A�Z���[)�(O�q����4�އ�����Vv��D���Y���WQ���w"P�kw�
�����n�� U��J~��9,��R���+ޱ��c���-&"���{�A~���)j�d�So.�ݐG�����Mar��ɑ�y�ˬa�E�Jwտ4VV�W¬,�)��85���-p>����r��(��2���h}�p�pnL�G�8�R즱�D$wǾ�Jܪ08˸�J�V�wsA���
�/w�-�Kk�,��j}1�z�ӄ�+���)D�ȍ��P���K�	n��>5/�PPL�K����+)zg�� y�ԕ�]�a|�~���hz�+z�W��`C�,�Fq,�I\/h�v��pqU�9t�L=/�����v}��Gû썾yk�6ȇ��/�l��F�����D@=�6ص�9���v��e� :�L{����a)�4���_�g��]�X4��0P[<4���.LZT�6��<����'���02���+0�x�lb��>.?b=���A���{o 4�~U�6������X���Y�}�4=�	xٙU��r(��參ް��XW;��L����|OS>����O�� ��5���ǵ��0"��g�8O�N����gU�Wf�-Y]�z�a?+*C!?��o�|cкC�NI�b'#uk����PhczLƱ�E�Z�3u�#��V��(C�h\��1�2�B��&����r/:�Q<n.�t֋�>�.�p_��l_�{7�7j:�c5��-"��$�>�b"�v�||�O~��z�K3݉�����1H�g�Ɂڤ��Nzm���`�/��M�������0�)��+�g��g��h�9',����V1�A����,�#�2�&�S��%:3J�.�� ��hL���$�z��fM�%���rb�󔀂[Q$�,=�W^p�(�X�/�9եT������OKW��m0�E�l��9B�D2HM�I_PƮm:YsaU���	 �q��mZ?dn9"�DEs�U.��77�UJ�>��b�o�y��s���� ��\��p�~�>�p2�N���<vU�O�Eza��v�����NL��E>T*/$��ח����vW��zmH�0.w5��B��7����F�������ؔɃ�'���Ԃ`(�)��O�P��jdIi}��q)i��?9��e�`���V�d�.*L��D����u�HH��gC���sʠ���khY!R��p��`1Xd[��e]H�4ԇ��~Go!��L(��խ�$8�G�uA8#��X��d��TS~�X`1P%4X��챎Y8��ũ"vH7
��Y3�:uc0�h�����z�Q�7x2��e��4�LN��ْu��
"�����PǄ�/+U�\��i�(
�&��eТ��7��=�7֫�Gl ���V}��F���T
D���NV �/X@��d�$�p���F3���f�L T��&	��\�UTb��gK}ې�X��a� a�4��=n�����*�2S0rdQ`�����j�m���8��AN���a�<�gƺ����, ��'��t�yʀg�Aj��+-�d�˶ŧq�����?B�jO�D_��C���<�A>2î��F6�`Y��ݢ��Ó�yp:d���@�L�������'��˼�y�^[��~����}�FB[ �=����E��\
��]J�G!E{�o@�Y��y�Ι(��1C��f��K^K�n^m��-��+��i���6C�5���2�Vs��)D��<mlN�~ca=���G�7[&�N�����,��T`t��:���|�R8㋼��MD���:��nS�F�(��fw3[ӱe��/��pl�P ��b�q���i*���q�����k���!!�U��D1w�<�-�>VZ��'��w��,n�f�NB��Ù�''�2�ic��dC"��}�+�v�>^W��X's�b�'����  �J�ƙ
��As�8��S�MK�Mt�2-���$k�R�����/%ಶ�ޤCCf�J�t|��q?DA;����gܖ�^��K /y��[hϸ���m������
�S&EK��ҿ��̲j��.	���EM��q�y-պȓ6J���w�3�������S�k@h� �3D���b�7���W��$��:�*��ϫ�J��D(mH�K��D�W�}���kӲ�x�\!IYA6�C{}�=��S+��]�̡�KH}����%V�1dz��ݳT!A����4�ZaӍ��u5�������h�{�ˮSO,�,�F����e^�2ⴹ�_��F��zжCmF�Ҋ�T��Ž���L�>`��-�g$V_���b����}�˅@�������sȁ�~^A�W��]q6�.��AL7�N}i���+���sX�eۧ8�eE٠c-K�p�l�=\�~6��C
�(v�l|���4h[��#���U��O�~��x۲M�r졿�)��}�d�P�G���e���x�<`�1V�dH��uD$�O��:u�y�Dw(�Œ��H1K��=o<��� �䚠����OC��N����s�á�qg)��u0�h��i<Q��޶�=)/'z���n�p���^�/N ���&+����	5�����<��ֽ�f�ft�V�e���nu� e�^��Ԭ�T_D3��P6K�Z�-;^�[�(�&�M����W�7k��?�R�&�	�HW<���A�����%�h#�Bh@�5'7 _�b {�ksLȣ�Y0�,M;���nE4*���P2�C����ps,���q��!����'�%7����x▻��j��) �Gv��>:En��@5Ml�ǥ�<@���9Wa�<��};@��_��d����b|3e��]2m͂ߎ\�%t#%����`,)����qj�3)���M�iJ��ɉ�`���v_�,;�?{�s�Na�.J>���/
���ryG�~l�jP@����r��(3#M|�Y��bV<�0!�L����՜B�27T�X�۵��"��6;�RG�m�S�$�� ��<�81���)xk�l���U2��9��BM�Mj��m'��@����w1�4G�j��NM���?��mP�m렽��R].�?���\2���e8Y�_�.�b����l�^1�֋1UTD���\�R�p}ʇ�n�z�"Z��7Nb؁�l�C�=$ou�Qv���A���e���@�>(l��Y�ar ��� d�ZY^ö����#
Uj�����$��� [n��f���Զd+ B-zDB���#�]Gw�	�FnS��]��E�d��^vq����%������B�v��4IdT���,gB��T"X��U�ۯ �-�LE�Ӣ��r�a�_=����J���ϧ����'���q�Å�pg���#pA��rl���6[36�*�
#�����.��%%�~ߡ�d�Zkv�xĘXe�T�O�}��5��l�t��N��c?�� �}�o���u9<��L#�T����QU#��V��";�.M4C�ׂ�%���]4�s?��ܑ��yN ��J�Ì�^���-���9Wy{��m�l�e���m������@�,���A :I��t!�U$,TQU��I�zr=f����o�1��������������Ӥ�#r A@ �sW��/��y_�]�<�������F��1�(��e��M�3Up����Ko�Ka�;㋋���W��h0�{pZ��7��e�C��,��z���^`��������d#��Ѱ���8��H���pVC�ƾȔ�gtv���Of�%��xsy�2��Ӎ��H9��`P,U(ֆ��u��G�J��6��N.���2��+�/v�[D��0�n`R�W��'�e�:�[*����o�t�>^|�w5�jr��O�kD���$?Ed�Ż.*�t}��x?�o�U����JL3��)��k�$7t�Wc��p���q��^��/�Z�9��k��2 W���)�D�"}��֩�e>(����f�R��e���ʴmwU#'�>x�Җ���@�{~J�D�S�������ʗ��]��	^X}�OK����ߏ��;���g� �%��ǡ[3/g,�p��Gq�̯�_���.�O9�����<�?�;�K��F��K�S�c�������ƕ���!j䦿��$�5��M�7(
 f#W���*4��in�>B��V@��;J��'���n���K�Z_�z�y1usM��?���Ix��I5h��"al��jB�#�`T��Ì��(��C���A����u��`�l����?��uU� �։�c�`n��,=9<�Oр���oUܲsE��GCw��S�yD��Vb��ƌ�L�����#.�]��T���fc~Aӌ��ÅO�6�"yeĝ֫�/4���đ����VB�[���b���5�g����Σ�U~�6�Is�g����B�M��E�'���9�ݹ�Ȩ=�9�Y&ok"U�z�1.�#�0���A��������ky=���㠪nٿ%�~8�j�: 6]��:�₤L��ga䏩�Uɀ���$��Uߛ�Sj�b� ل��;艁�X����2�����%wȝ|M��9�0� �<�>)q��c���5�u�vZ��1sVH�L��L���U�/���Qt�fH�*k��Z�>M����ocMf=;e�:��tJ�&WF�`Jx4���@�V�r�$6���3���;�J7?|=����ŌW۽��=��E�S��Z���.˧�	��q��R��J�uh[I�й=J#ܠ�	�`|d� �ҿ�Sx��+N1�������[e*��9b�õ"��G���PߵrA��V"W��f����$�����C�n����b4��3�Q�<����7`�gJ�\�6�"�����,��Y�p�u�a�;I����A)w	����Ǌ4~��=�I�r{�J�G�廅o���H�K_�d�i8;e���xq��������`r[w{���i�:!��P��{UӀݍ��z���Ӌ΢HG>�ɬ�1tb=�B� "��L%��Õ�b���*+{9��zȍ0����ψ�f���Mu`��(jǇF	Ql`���	}Å-Y�hP����\F����Q����dz�����瓇��'�!Y���Cg|��N�Cg��<�k���{ZP@������uT�l����ѡtJ�'UlF���,�&]�.b��89�m��0�܀1alW�'Uþ��Ate^=h?|�b����l���}����K-�^&sGf������Ϣ�H��{4� W��t7����H�ҥ%ȬN����W��}�B�$%�]��mr����s�K3g%��<���R��Z�/h�cV�4�q|c&*�b*ev9<S�.� �W�� �E��uG��Q�`��]��Zl��3�H'OR0�����
���Ǖ���J��ǺZ�����8��GZ�7���A������]p������e2��R��+�9r��#d����3��:o��8�/�;�M�wg#Y���9l�b����	�8RFK��XVb�C�D�0��܈P[���a`���́�FSL1L#bY�r^�`
� ��]�ܩ�x^��^te�	�������&�UV��p�<��=�c�Q��c�wJ�x`r)	L)|ı���-n{��%�\������)������0j��˸���tp7�Zv03��*V�O#6��;��ҷ�\M�54Ǹrl�@� Ɩ����Zd���4C�'	����yҲ�	��w6.�]U'M�_��Gm#�a���b��:03$�"}�˛jJ1��>j����{����=T^��qs�0x Z�w�$�9�֔���>��KU{)ܬ�������X��m� ��rF��HS��U�����]�X�`�#�3	�s�3.3�ن���s�kD?7���¾�ӧ��I���N��5�vH;�{�.]'���B ��IS�	���㴥Bn?�琥��j�X��ψzv��(�`E
�p��!pZ�Z��?R�0�l�l�5cKF��
q�L��#Q��o���\�^$E�	p_���ڮ>=V�fI�3�Q����,d	GI������X��ǟ��Ļ��� ��?޺�ӞmBz���-�x�a>��̖9����0$U3� ����dTL� �����baS!e<�T�JO�!�H��m�FC�Ŝ���:��/�<1	�������� ŕQ'~��N��6�*^ʜ�ic �C7i�5��Ȝt�I�$p�>+���9�~i2��Oj�K�)N�ad�/�f%Us����=f��"��بN�}����NսU/����1���Z$f�e�zo$O #�~j&��Q�E�y�JS�L_��hB��'͆-!Q�~ƺvhg.�a��j��ī���f*���$��y�؍>���}���?���R�
�$PK"�S��[~>�X)�ƍ�7c��z���i�C�|�1�7YZ���d��M7����T�ȼe�wְ�5�?e�5�c ƕૺ��da/�w�JB@�S�����$/�i��O{��jL��P�� �.��G�w"O|>x)f[�>���}Z#]���|�+x��QT�CY����C�����J#D�3q��� ᓘ�����!k/��H1*� �.���hkK�'a<�f�b����ت,�k=a�l�F�]w�P�s��b���o��{A VA�����s,$����p����G^��;A���v����lB#�]��owW?��*}s?�W��s�\Z��J�Z��(EMu����R���5cT��J�2��⁠Y��^P�/�LF �T"�2E�@F�p�tٴ\6�/ *=:����u�7Mׁ!�BS�ok���pU�(����L�Y�*IڻG��*���l�h�w�,倌p�X���%PB��(?�s��vם�)���d�2}�25ڝ��HK��E��%�s��g�L�w"���3U�<���"�5�[V0�0��)��հ�{��J�Jw�#�o���cǙ;.�},8�7�+Z���MSF;@���m�ׇ ��;�UK�zAq�T�8w�u:^�����LF�E�B�	�3B����ǋ$w�u�x���_��F�9x�����Y�>]�?�Y�Ɩ"�b��lX�|��ݑ��u\i_ʨF�� ��&�WE�P~g�bː��1tgKr�
cC*��Qb��KLdI��vp���_�h�q�vU�ԡ���O�ȃ��3����֧W:��էU�\�bI�gSF�"H�UH��ch0��ߋM��{�Q�0�DEL��F�#��%/�����Ң��Qw��+����D`���G7�^IW"��v�m2�C���L�i�,��2��1A
���V虦��n����5���k�`�~%�oo ��Mo�X�W٢�����:VfC�'!�*�����1���(�����r�.��3�q
���R����e�(y!`�ப���#$N�Y �AH�c�!wӈ&�4�{D�n����3�� �Ԝ^ ��#�%�@��n�y�=����)��9��u��ɳGQ)�:5V��L�1�Z�,���G�:.n�/8w[\�͢�͢6q M�1�CI������HhK� �i�Fd@�#�*5?R'޲�w&�zf�~��3$U���ĵ⋃J����.�t��U��s�u��1ޫ�K�F���ix�ɢ��q�]��l����c�LK+��J�K��|���o_�`�lP���K���ͤ];��2Xy�NÝ^��#l��_/<��|�/tH(��_�9�Se����T��������^�'r��ɜu��M7׌+0��5��s�2�5L<e^��x�̥5�����|PEʹ:Y�Δ,��(FlQ3��N��mVw(���ޗ�Y�*
�9"��}p~o-E���\��3jH���4��j+����h�L�P� �Z�U�S�|��������Ť��j��d���^�5>����.<L�nlY�	1�k�D��2[��~��ׯK8��Wc�O`9����x�$��U����3�t�]��+.���!����i�r7�34�`��`���
�mU���M���'[ `!`�w�uh��a$��`
OnLꉤ���\j{��0�_}G9��nlZY��ګ���L�
AjpͬSop�L����bB��?���t�T��*ޔ.�3�p� �
ё6܈��~� (n���ڃ�&~ ���x��)�h�ࣥ3X|�a�d�e��2�D�v
$_�+ ��3�#�դؑr��p�
]� ����F���k��R��?�ߡ��ߛg����<V�'�Xq���S$Z���q�����t��@;�	�W��U�־�2�����b�{��� s�� ��n��=�a��x�D�xU@�X�����D��t�+6���Ei�� ��A�QkX����U���f��;�þdR��t��E;�IyMF��&Pb������ċ���\~|4[H'_hA�`��Z�}h�n����8Wˤ���q�t%��@QI����X�v�.ܱ��*j����7�H�T��3�2�C02ʹ��j��X�IL!p~W:h�qg��J�"���j[ACC�wvk�q���P�l�,.(n����.�D�����SJ�	ihX�Q	r�&�t��$-8�� ���@.�M�����#[��V8����0_�z�����;	Bh-;�"~Q��Ӹ���:v� 53��Q�E�e�FSd���:��})�/f��g�S#dQy��vg]�$��$�zZ��E�º	��Y� D*-�݋<����b�jmz����t�d�|fĉF<˝�*�#�~\2�CA�δ���B(&S�]��o8K|x�.W��/��H���I�Z-G�3j9e����R�̒��Tk&���&׉VQz�©���;���������F���GE���o/���s�E5O��0��v�`��C���z�-��>��^ҞK^`�i��Cv���+cb��X$dv�Nv�����i��.Q[@9w����چn��}Y�Z�6E
�:��} ��-�"�WS>rX��4}t8d�h�١{F|o�ʗ���6��Ok��1�^d#a=d�eJ�Uq�@w�$�On헙�)�3xB�ʫ�R#�sB��S#�԰�t�E�[�S �h�s�Y�Z�����+�	�T7u����>�G�RL3�4頖tu�<.�̣�s/"�@>�8�0!�8y�wC��+�.� �>�O���`��$F�x6�0�k�0�u-*a���
�k5��1(SP�HZ�_���}���g5��r)�t���t8�a���]u��謆N�4Z�1h���:�t"���ŗ��� ������u�߁>��'+S�&�o� ����I���sfc�(՗���w��t�jWX-���k��h���܆� �e/"�9�`DQ"�fG�zh�d�@�|V#bBˬ�:C���2���W�"�!q�$+]e�wb��E���X�D^puc�]_3Ka.^�T�U���ny�ַ��v�ޟ�	��I��Ք�g�����l?,���W'��`�^e�W���$$�K�w������$5ɜ�ъ�rN���򅾳��-'�,i궞5��m��%�v���~�8��|Y~���)�6 uC>j���Qߎ1�y
ȼ�{�8�}�l��.#Fم�P�	{�Ex}�Rx��rD3�
�����]��؅��#�vہH�N�9t{a�o����X��N}ya�2�\��q��iK���V�o��E@��6�[Vy3X�O��ޭ��ټw�/�V�}�| &�T���X �}V3��1�Ӏ.��Qu�C�2�Qbàu��W�j�w��#���Rؑ�����Uk�^N�uy�=�Rg�P(��M��( S�(��y��uA�5.`��ZbN�e�]0r飂c�(˒ЩBL��R���s�mrԛ�+���[N�ri_u��٨+�mq�B5ܦf�V�!�/w�z-�~"F�>���K��ߓԒu��,u�јB���|����2�;��k�11s$���$�߷�,��DC�{�s�y����0tJ��}�5G����`K��HmD��׼� j��x�T戄d��h.���u��!��o>���� ���ln�9��"1^G%��!�)�)Lǧu]w=�Z�����eG�?:�&����oj�{����t�W�V+����X �S�Zz����{{v�sѐ��	�h�4K�Q���)L�c������d�I�f��;Bv���%���`7
�z�!�]�?R�t\�.��&_rHģ�{6c�bo)�ܽԉ�
�����I�I+r�C��߯��{�Sm/X�u��������S�Uk{�8�N�r�Krf p�!:O�<O:`�\/��\�����TdY��-N�4��C��ZO(%ɟۋ�W7��oA�\��ُ!D��0�e��.�׃nF�8cP�U���UX�9�^�I���B'hH�h�'�Z-q���S�|��85&S�en���饘^fp�ٴp���"WqV�AX qr'�@e�n�>�v����E��8
�<K�pgyP�����c~�/l��֖���|�e���9����t��GS�A�P��AXZ�=�k���Cΐ뵓o����)0�Q�@�Вj�S�N��ĭ��M�^�9ճ�Q�*����g�^�\�޸���첥��8?ď�Z
� ��_��̫�$&�3��|�&�D���s��sW0�rk9��k�O`��.#"7m*����+Y3�x�ƩW�<l�(�'����5A&j6���Ы��ji�����'�ˢ�74vm���3��e��X�O�<+�k^.)�M/~����A�:��<�yzy�!�!w��MtE0C���ꞅ�H#P4�pB�l9�D9�a9B���x�j�㩰��UɮQ��RQp*t<l�y8�@: 5 ���a����bt.���f��W�QO���d<܀���z�ʤXH`�>o���l'>��Hi�J�7s>{\�(�C�r5}�oF��	��H���>5�2l6�"���=Q�dS�g��2h��` 	��u�.�GO��˅��}�4���c�C�BF�q��A��Bѐ�н�ޘD9[u�͎	22K��@����!�|y�Q5�~��.�Co,i��8[�RuL�����U=7�3 �h�,#^cd@�w!��3���{�g����~�M�H����b����,M����7 ���I����j�Y�s��I�a��-H,�g��H�X��W�Y0�:@�*My��w��v�yq�+��#EK�E�ǼR��o7��
�xF��ؕZ�/�;��-f� 1�d*Έ�-�:�6�ז�����q1�aňd���ſƷV�z�X�c�ҁ�'��7���n�H~H�Z�u-�ze��}t�K�)=�7 ��)����S�D����e�d��S�X��OFXA�+�	�ƃ_���,�e3���а�/![Dv_��;�y��zn�GA�N�6vv�ei��蒣]�"��+�TK����j�!�S�D�.���ͱ�*H�0��&)����=x��WF򦡞��f���㍭��X�:2w��N�����B�
G����E]7��i"��<d6.Fr����S��Q窹�)�{��1�\F����d)ļ@��� �@v �V����B�>g[W��ʭEns(�{�>�N���%K��&P����/�|+�AP��v�rHy׶��ɦ��	б&[���Nv�[͏7�l�5F�{=�p��@?C�r�sTU-�JA<sΕ�Q�F�(;�)s��%��0��ph%`���E��˿�^y�^��c���3]b����P���k��1=�mH��(w����O��6��$���Ċ�0fjE�m*p�-��]��1)`S�Wh'�2�A��.����4�S��j�-cp���5��G��c&��k�������q����bV^�vqn�w|�%�.�z��Jy2����*{�$z2�7�����~R�ͨx�k .5��bcV�F�o�ߘ=�l��5�hq���'S'�xҮ��ۚ(_�s{�A,�&����sq���RDT.uol�ߍLX'O[	�3�Np�wUMWC4��/����H�#�	�©�{Xm(��㙺3�++�7�r���$��r|���T;K�D=E}�(�"��!!d\n��Msq�یMc�����Ӗ!��֤��N�����n�_@jH�9��_S6� ɬ�CB�T{���Z��gvx΄Dݨ~Da-,��}�ĥ��9��܉��
4�A���=n[=��n���s$c��C�E�pqy�T�ɓ�B���d��9/?�lm`��5�eC!��@�$���Y�WCɾ�@�nݽ�����=r�'�A�v��y�\��B&�B�
���a��MKrr�c�����ro/�����Y1�j�+R,"������IN=�<�nAc�e���UPiJd����Zo�4����1H��^�'8Ӭ��O �Fo��hR"�*<������c3�VJ*-��z*�[._���RL YJ�a/��N�<[� ��*�T�>p�&����I�e�,*K��������Xκ��b �F-�Z����%�;&��n�c�>��-�o��3k�}0��a��8���!�\y$�����!����|<u�w[�*��D�8�����E|e'�,���E�{��"]�$!ۏ��ܧ_��E��T�ѳ�,�n��T$"�Q�`� �돫��g�g�jzZ�1WqEV2����-2�1���Lj�3ͯ8��,[�gV�U���~�K�@�(�hē q�ڞ9��'�]�ҘYO��<������~�J$Ԧ�Β���A����ύ2[��&g
g��QvP�N�>"����;�O��t�����4�	�%���U�������y�l��ڮC�m��A9ZE�6Ť�\2��q�a�����~ZP�F�ݦ��;߷�	�,�Fm�;^3�d?>cS%��*T��&���3L�õ��y�f61�m�=�ιd���L�w�BK�]��&�h��	�w �|�l�R8]HC��h�Pi����W�2iO�r�2Z/�V#)6��//4�E�s�w����}��S������ j�:����e5���D���S��{pm��<�~wv���/�]��i�Ԏ|ƨp�d�^���qa�W��U*6=q�]@���~�S�����-�� ��f�NYM��43E�%H݈=#���s6�O�Q�w�e/�V�Q���c&	�خ��Ld�����]bǲ�ڦ����=�.�-�L �kI$��"*ڢE��ua�c�0��v,��Y�����:ڠif}�?g���c�O
�ؕ�0�Zow�6�a$��f�M�k��.�B���W�Ѱ2�!��A�(�!�"i��7� ��Ȑ�?1���5d�I[��.\�L����W����	��[s�����dg��N��.�*L�ƫY;`Ō�n=�Qؐr� /}d��1�_=e��zO* s����$�L幞�s5�T����l�(���L/h���K�$J�/� �j
c}��Y0q����J�ݨ�� ��B�o��M2K���ab�����<D�Jc����a��\ ��e���ӗV��Xy��y�G��;�Gݱ��b	p����kE�ʮ�a��|�1��js�e%O0r�^�����d�qEd�>`�$�����謾r�au�U?�1���(�W�� ^� ����8CGқ��;��{����Ͽ�5�~}�a�������&��8�TiX,v�/���ʔq���#�V��� gS %k��x�~/�j�R��m�ͲJ�_���f�(A�e�/Q�a�3i��q�Mf{|���<&���uᲈ���E��~��lyXuf���9��aY�ƕ0��*�Y�}z3Ez��b���1?l.�ӷ�����z>�29�^���L��� �����r���ML������4�~�C�ef�	r��
�:;y@P?&����@�!FG�y���x,U?/�?f�'��;���Ŵ� G�ΐ�� ���~�v��\i&>s	=����2=U`Tm����Q܆�=%�I���ʇ���h���4@8�C3<� ag��T�v����T3T���FqW~�	c,��,�;\VTzmꑸ.�şn��v�X���"Vϫ�i���O��`����K�w�:��V�-�s�UV��+=P��zB�]�앮�؟�"���N�NQ��HAJO\�A��ʓ�Ԩ�M)�>	���>rE�8#�t9K$�M��@�>�F��*��mrJ���N��'�݀˺^��qV��T��0�OM=8è��հ�IƮ��TU��~�T���BAGV�p��\�!Lb�������r��cj[�hD�˫,��82�jJ!Ow?��T�mh��mC�L�� /Gj�u�ID��3D�2���pkt�7l�;�VX��4@�����4(쒤f]鈠� `=`e��F����7�'�D��х��*���C�")~	A��%:0�2S��i4�eQ�G�4'��$���PΔR6�s�.��J&D����'�����z�r��7�E���:��>^p�&�Tr�u��G0���嫖�=B�<�&���V��(LF
+i1���@"g(x�W wu�Ot��ڟ[J��/�X��R&"r�tp���lv+�Mִx��%�?Ng�R�_�^��{��O/]ӳ�i��t�
o�2�*��3eOp�2�rC/�G����%<�/M�	f��Dd��w����{ᰐ���~	Ϲ-`)�����x�Q�5������w��Y�r�ƺ>Z��^�� :���ڈ�c9w��_{mX���A)A_h���aΘ丷�o�B�-��{/��Z�9b��p�>c��"���KF4[K���7���TW�<���{���,����<��g���[@.5�C�u�+Iʌ�o�3�V���+���]5Be�q���P��Y��}�<���R�&�>1	�!�蔼���R�wV[-5�D>h^bB����	� �`�N��)a���~���4�����V�֋T���_���˾]_�Ċ!�Ժf���N�/(Q�@����r�NP�h���-���*vƵL�J$ a������U��� -/�� ���tE�D�e0��^�.��bG�4$:��ڊ���^'���jri�;�!S��C��?�g��8h�M�����=�w��}�W��c+�ugڬJ��^�i��XY�'��gk�m��F�Ǥ��aK���y��'g|_��V�˜rP�K�x>,�o���A��o��	p�;�H�!���nF������sR<�ou���/�f.&�-Z|�4����H�v������q���U��GQ��<���k>Q��`G�y����5>�Qg�b��][L�Ԋ|�s�f]K2�ݽ��3���W��#�e���0Z��zD�C��J�}�S��I.F�� �����	��9��##? `�=荋�q��� ��'bM�/��'�1�&N�~�\JQixl/ә���L��Q�#������c{I.�������O�[���(�n3a{��-�����W3[��뷵r���O�+l�]�jkmO�SD�A��vS�E��p�C�l��Zx=o⚰���sn��WD�u^4��;�y����5���&H��ޜd��H�R$����x6z6���/rW-��D�l!����Z�KA	Lve�Tc���a_��k�Q�����O%�����q�8�4#����.c��@t}�yQX�sIF�+�����0�6o`���f*��R���o��h��P��o��\��̉�^x��dӀ-�[d ���/&�IO;�����l�Z9�diB�y{Jb���{�h�������d�H�� 5��0އ'15�;vJ�jD#�	�J%�5%29"ur�J�;g�:L�_��L��x:�JT_�<i��r��C�,��z�4q�5��ϒ�A;�j>׹���$�N{߾��L+�F�<�P���;���,��������#VӶ�^�^�.�֘=�������!��u?�~�E1�	dW$��9%T\ߐ���z�j������6F	}���`��k ����e9/��N�1���·�Yg�^/o���5�fS_@yҗ�95a��L6���S�f����1o)�l�A��Sz�? �ҁ~�����՚���dGML]�r��\�}��c$c�,��Kn�q�������� yvg� ,l@��!S�G�� c0'�X�C�d*�ԘS��TdTu��L��e��z���'V�C��$���x�|Yt�bE
���;I�8�ߋʉ��;@�=��7���� Q���r�n�P�z�Ur��i5���6������9�k�c��B^��x(E�@�+4���%W[��Y��;@P��׼����+'H!��
�|�X��r��F����}A��/F�"\YB �#,�N��Ÿx�k�(\�it�L�$�]F@u��a�K��""|�~�T�e<
Z#�6�ta�0U0��'
=F̻,P�R�T���6�J�o��l�*t��mۡǩ�������u�uR�F�(�:���l6��~&9�Zh���\s��
�'�Y�]��Y>z8�z��G'j��� D�RDE8T��o��?{�5Hn�0��+ Ə/�!��4��w��c�|=�P W�6���5=3�Lk�Dc���v&3�r���hъ� ���.O/�3Y*3͂s7��_�⍟󠮒}p_��K�#~f�4��.$��t�����Sl��n4ҋ�֋EO"6^�]���^�#F�"Ю*ñ�I1~Dήh{�����Cxm� 3�=�m���|	�%�[��ƣ�#�;�ɐ�;Z���������II���er��Ei���p�$O-B��C�M��csEc���­�����3����{_�����+�B�%_/C�ќ�O�\�h�����,��p ߭8�
���@�0�$O���l>oG3�h�h6�h`��^a��)�Q�O�|�Ė��R�Bа�\9IP/]���1ښ�Z�8��ԩ����jRm��\�gCcaԬv��b_*���T�6w�w<���Rf�8��aE���I�̳ڏK(7���L�-d���SLf�g��ݧ'F^�N?]w>�u'�1���|s�)T�O&��O�IK�a|\L�L�)���HH��k;a^��t�����5%�q�=Z����P�B�$�T
���Ki���8��tCd%Z_{#*s��߭Q���~j~�Ԑ�T�������Lo���F�Ԭ\	D&��J;Y���=#����8��7��}��ܘ9���t73pE�~�bNV,�<+L<��(��|���&�N��ȅ���۠�}D��:	��FY�՜�޴�΃]�2������R6��oؼ܎�^)�SBMr����p�����zJN"�S�m���B�Z_���m6:�=�&�O�<^Tdr�����$�.��2���ΰ���rt�I��cd�QSA��^,n�pب���y=M�0�wy�ٯ�@ �o�@��{����}�v��ű*�K�Cu���W��)�^N�LfȖ��oeu8�ry�4�
Nº��� ��M�.�0�.��R*����7IdP�L7
ʝ�D	twDŒ8b�g.�1+�Vw��Gxjh���oOJ!���#H��m4x���R�rO��J��Z,b R暝���ȿ��g]�쨡\�������3�۰�U�$�Z��l�ÌA�%Z�*��SUW��)s>[8�P�O|!J������1�	ت��	#����s=u.s3��Pt,�)���(R���o�S�ϛ���b��j]�	���n��16���,���mp��1"�T&��i�c�-�����Y�1&�Ė�m���0���$.!-	j�,'T�b�	�d�������>kM����եϞZfɖ:��2ç�wV����[�H&ﵿo/�6p����Pǵ�e ����_gN� ���8~�E�z@�"����׌�Uϕ>�m������q�� %�����������A�"�jX�(P�]��RS��=��&'�`�����[�
~�H�����a�Lw}�Z6� <HA�h���Y��{�"M���	�H��x��
�c�CF�Y	k������-)Z)���(����Y�\o�\"��R&������!��Y��*~��_��vxn��h*��M�N��T�q&�Y\P��Op�t���H�k�
�Y���+�w,z�E��z�ʐq�]?���<q�0����u�&7�s����p�E��;\Bz�_�'�X#�T�R��=F�*�W��IC*I�%[�U�y<U�J�΄�T�<�G�0��ӎ�M���r�ﴛVW����.�R�<D6����q�bf���
�3�W�$�y'�&���Tζ4!���fQ�m��-А�������ݞ�] �
��l���!ҁ�oU;Q�;�?BM�c�!L�F�� z���5�u�����>�R��'�{�g `+�Z3o,	:����f�9����v	S��k����8�w��@�f��5�}�；��x����w����Ow]�Tj���e��W`��q.��2x6�|��"�B��L�!�����C܊��u�	��J����(G\g���5��'ޔ?�
���m`@���=��tm�;�ƺz����&����[��n5G[����e�n���wFT
"lc�q"��	E��I#��PxD�y��D=�Vz!0WL�tmرPG5��O�k�K�g89FR �E�^{B�I����72�6�}�bUr�y !���eW�JbB�����cJZ_�z�}���~�����Tnh�X��N�X0'Og��e���)�m{�5{8�u �;N2�p�T��ʕf�t��˶t1͵�Ю7�0���M�%�6�p�b����!F�8R"8YV���4��ZI���ލ1��;�
�j�	�2�߇�`�y����^�Ұt��U�(T��R��Pq-o�v�S�(�Y5`A(�b�c�r����^��+a3���  سPM�)4�N牃*^M�4#e�a(W��̨��-u�g��S�s���ld�4\=<Z�3�T�a� Խ��6eA����$��
�ׁX�+�?􈾐S�D�����!�/����s^vm�*q���H�6��%E�IQ��+�a`|���k�M��!x9�+��f�G�P���.��ue�jiֶu3�VvP�5���������a]Z�>�W��wb����\���R�U	b���MwD�|:X�G؟�wĄ��B�?�8(�p6����+�LgB�c�\�N�O���q�v�����$1V�y�P"����"t�*�YkL̪ކ��|^$R��-4X,,�d|��o\kLcaM�`���@84�n��R2g��}�n{�M��p�e{�V�uX��',��\@��$ :����21�'5&�Z��j5��14�q�5-�2���4��miꅪϱ�t1G�m��*b�[5MZ��>۵ۋ�
�#���S;���̉({�nI��S�,���?�$��Sy:���x���Jw���Da�����ҵz�ո�i�2�k���K���Nn�K%�|-���<���jٚޞ�:=\��и?
H\?�:ϝ��ݮ���{UmG8�W�%���6��8b�ME�d��\L'�1Up������#�>�6�xv�=��l1�����)�|ı;	�p׬s���
U���Y������Gs�	
ТT��Ԩ�O��<�.�qDH�q������
�8�h��g��v�,��%G�.���OЇh�`���*˪�"�?�0ۖ�}�6�5(�����J�bؤF;����kuX�%��?9�w�����="���$�wҾH;��l'A����,#�\}CC�����z !�gwqe���U��Vw5bt�Ɖ�wc,��DY�����9�zV���i��x�����O-�΃����j�,@{'����3T"|�X�o,��<ŁPe��G!!�q:q�D�_F��CZ���ɚ��2O��M��8�������V��n#}�|\�]ؤ$�7s�A����T��с�~#�yY	��G��?���$$���A�oO�0���	T@����04Zch�D��tP����g�;у�dr�<����tC�������8���^�ѩ]g�ެ�b>� �P߶�i��Ff�o�S�W�v���-��Gѫ�O�o��պ5e����˖���=!ƃo��
����_�~q��
ڧ������#���Z��N��A����e�E.�?�u�N�ª̮}���]O���x�fW%Q�z�7�g8�e��Q�ԯk2hըz�`��.x��6[����3>=H�)����e7֟r!�ɶd�g ����A��(�8�O���^�|�h�ya��b���qCO���� ^��mfv�Q�"���E��=���Kq�k��Ji�$�>��=�"�61�)�]}�X{�(>�~)�X���]a�Q�?�z�}��U���g(Ή���/�'�^��͗͝Z�h�O�� �`@��&�%���6'14�����O���� kr?Rm)"ot��v����~U���R�������tRPcђ
�n���1Ė؆�֩"�Y�NJ0I�^��ͧ�W���B��(��v��(p�*�.a����NąS~'0�������y7��32zk����}~Ǽ�i36^��*0P�yg��(GuOJ���t!�|d��$=��W�Z+
��QI܌C?��΂�j3�u�}��g�n��b�Q])��65�q�W��a�6̑��7�|L><V�&���z�x�h|�$�< �����T�K�������g��1��|�и�I{�b�+Q����ϱN��(���asVX��������%8��;dw� �O��R��RZ;��D���Q��,�;t3���8����2�Q�D��T"�Zj��X[�~�f�Q8���f���bw�_x�v���9���$k�C-chޓY��Ə�X�VZ�M��b����c��4�]���r8�^b�	��֣��uf�<�e�o�N[,��=$�e6��8���,Ħ��V�6@�BK�V��j<!?�/������%X�fy�̹0孙X{�;"A�N���x�����[���\9���e�
,�L`��9LB �Te��gco7��!��n��ǭT8����8]T%,�k�Y��5Z����V[�>��Q<w�&A�mc!(���u�[�dŞc4��E6�/���)�#`� ]C�"���;U�I�(��N)�{��E�*y\�~��M�@u�`��.'2EKE�U.+����,�Iw99�L�������C�kS(�;ģT4�P@�	�X	ND���@q�7������@"Gç+û��:���>�5�C��~�{s-���8�B��85�{z,"柀&��`�fN�����L�	��
z�58x%*`f��WP�&�ꔂ�[����B�,���m!�?'ˋz_&.���{qP�1������7��&���-�6/�ML�VgԄt�Qot���z�M2�k���	c0�\ǥ`Ǥ[Օ&�a�8b�`~�1����ڸg����q��&.�.z�\Ԧ������O�&��h�5M�^�c����/���ic����*V��Vy�����܄F�W�^%>����g�e����7�3t8���0�`Ȧ��Q��j�s4�[�D��<� ��U��=/L�k������������]'��#�MmA��.&���<ۮNo�?�<j�.�F/��t��Ds��O�b��Z+�<
t��Rk�Qu���	3">aґJ��Ӊ�!����+�I.�Rv˼k���,�J昄���;m��<br�҉=��y��tl�KC.�r�H%��1�eN�����d7-Őo_�S��?7��ru�p�W�Ht�%�����Oaܲ�5E&�rr�h��_�.��t9&~���3�I�W*��
Xŷd����5����{�H��U�6��>a�	8�U���X�ft]byc�2�.�YHR>:rJi��&"8]_���@�!��/��f��F7�9��6����}�g5.s8=)a��������I��ī0��m�	c�㢨C��B�#`������#3�,m/�9���l'����O�u�8�5 ��g��.�}I�ŀ���N.��F�1:4���V?��v1��z���].S*7�F�SO�ړуQ������v!Bv��Y�@�������;�����j��:��G<�z|RM��blR��:�4Kk�#�yI��$��B5�3� η�;���T��%�(���N3���6i��	�0��bb�C���+�ʵ�N��?��kt�+N��#�Zt�LI�?���K�̰�\$؁i���|Ǻ�5�0t{�H�W�h��M[Hr���@1�v�!��%�;?�q�C(�b�e�}-���� ��2Z�s?2�99f0�C��`uJ-,�"6ED�T������#?Hx��[X�nh��.��Wo��u�wЋ��Κ���FeRa\I\n����A��8������xu�3��2�_�ν�ó���ʨ�Wc~d�����H|$���1}z׬':�w�!m����˞.��L>s7��	��zLt����S�zZ�7w��31���Œ�9�7��R�uj�鸽���>�ӏ)ۯ��P,^3��Ϸ"��%�Ng&я��`~c1�{��2CO��h�^��������c6������~���!�G�S�n��������f,0c9�ĚWb ~*7���x`&��n��X�U��L(� ������C^$S��A��;�>��5���7P�|z�O;O��5���Y�^ z�� q����v t���64i �̷�$7)n��y�WU��k*��n���l��|C�~�w~��X'sc	��%��X _ĭ^.�h�1�I�R�(�#&tS�z;@����-:�LIG|Ğw[8�ZLN(7�oU�]v�1NRD�=���"�Io�����oq� �Z�C90�/��1���i#��ʴ����Ux+�Nݯ�>�l;�yc��T�,.�73w0 )6(��F��KS̰-�9Pm
�$�E�%�Dp��;K����}PAD��[��)Λ�l�~����z{�T�6D{R�jB��fGE5ȍ�{4�*Y�����L�v�Ե�q� [}w�ҿbu�e_�=���A��@��j[�@�V�ٟ��h4W�1k"��Ж�jڜ����d�+?-�7�O���'� ���z�~h���ױ��{�����E%�B�uV�3X�5����Pd>��)W�ڀ`�I�<���5i����p�����O3﷖��<mL�ɕZ�_'���w ��|��lS��ܪ��_�M�Bc"�f�@��*Z�x��8�WWA�yI?�V�6Hg=t��~Te,q��J�{�բ�\q�#��&��x�l��b�_ u����\
U�ܬy�YM��+ �Z�b\�#�~�1'XW�˒�I���0ʎ]]5�=�w�+c��X2G�a(ڣ���\�(#/ju��dh>���8f3F�b��+���x�d�?���e�߬�Oz#�}=b�ͯ�SVL;a)�@��~Ss�2Ί.�֧�!J�gP�W��u�\�5�}f�'�]��T5$�����]��%i�(��{u_�� $��$��1w�s�
�n�fAD����u|�YA{B���^q�s/���ې�/��!B@c�a<tR�d�9�����'���a��9*�m�A̰�&ol��j
�D��7R��Ҋ��gcP�r�t��O�|�m��z���HϤ��ZR@:����9���z�Z$����b��2�3�@7�_ǵ�h8B�HF�苩�:��%�WMZ�G�<PS?�M�v�\���� ��	��1WL���c�=��*��Rn��y�=Il\�l�T:�g��	�i�:���aN��Ib��8��k�"i�&s9��²W;3����p{� )����0�\f`���8=^�����w��$ F�(�\���`A��,�FwG�U�Y��~*;6�p>o�H�>�k�0$��T�U�w�E4  ���,�){PU�-Vzvl�߮p,��%�;DJ8��x�nxo���(��(�-cq�$�U�nRs#�Ġ�;�n��+E�v~i�b�`i1�:WA�?�kxF;���+&�埉>/���Պ�wY|�G1�N��(¤Ņ�'!7zu�QF �EmJ�$�����;o��)Wр$?;��j��ŋ�vm�,��Sz������:Z����WM��2Pi�Q�	:2|�RcUs�+1�;P�J�Di�ID?w8�iޞ	nf�������[�OwEXx����!�P���f��l�fA�����Df,���YQ�s0��	�<��'�@a�D������_��4��5�w�5غe��Hd��̱qQׇi0�/.�/�Us67���_�y����%$t�g~�o�P�YO@7�����&����)�����zd���,|�s4޹���Jy�����d�<�X���F�3�Y�Ŭa�9r�хZ�72cҸ!��%Di����)7�w.���h��CBWG$U �"A)�Q��}�O�s4L;�ȍ��!���n���ۗm��k}"O��J�(;���ڹ�HuOG�U��co�@�H��Z�>F������\ ~�e��8����M#K������P�G^D�%ƙ�m`�t�Jx<|��[�����~��F'�7>Kw��P�T�n�c��U�\y��S
��T^�K?P�ŋ�������)n`!���c�x�sa�hȖ�&��~n  ^��`��rp%����w	:7j��c�.�z�^z �\T����H�ǖ:Tk�����Ұg��\���l��QV���O���U6R���@--+�����͟�%�o�+zr�S�2�@�N� 5��X�?��P1�{�`�:��Bb��<�,��љ���΃W��_�3\���ՔXM3SH�+:�Ӓl#@ITwӄ���$�}�'h7T!%�5���A�}=[������d���l,���ݱ�Ȗ�  �|*�,�~�)`�"(
.���g0l6'ڰe����d�i��(�4(c���潍A���l.C$�k��w���($*�V�������gn�b�^�C��G&��U�H���'F��5`�-\D�$V��tI���?x���ԁ��A6�*�<H��1�@��Un���*��&�R�C�#|)�,�E�w����[10��#R��3��_%MJ�T�{;y뮑ܺ�_䕂��n��:�<rJ5�Y��4�����=���.�刖%=z��;�}/��	�fi��.=۴�J�Oޖ�z�l7���m;͊���?eq�*��"��ENE#%@��U���ڑ�^�,�]�$���+\�-A��BB�%���;г�<�!f������(;�_^T��P�ԇ<�z~h�XF��c��k˙?Q2��2a��>f���)t@>a�Z�p�i$�����bn�=�w���Գ�uG�����*Q���q�h�P�]�=�>l{�!�X������q�>��O�K ��'��"><�,e.Ņ�CQ{]���BY�bM�u����?N?�DB�<B��z�L���6*����G��=a*�g��3�S�ҋw�(�.2y�L?��V:	<h�Q��4�sMX��9���pй�yvT�E˴�L#s�������կ3Z�+�t�ڡ �~ف�@?��c:e�qnq�_�/�ݦ�����y����s"��8����i�e��ђ��H���ϻ��s��{89V�*�ne�SZ�dP��"��� I��@�� ����#��;�/*�c��"���A+�}PkNr2�,�����+���A��@
��fIK`���khW��j1�)��m��[��Ր �p]ϫTz7� UU(׋1�Ó���O�	���e΅b���Ѐ��N,_��u{�Gls=3�tZ����c��	��B{Q�Rm� v���n��wu����[+%�]��d�&��&���+Ȓ�$uŬ��dA�y��V��<Akߡ����By*q�8�"��V	�J�������"���L!��q�����4l�j��qm
�����b1�Cj��t��KG�[t�k`�o��g�b����P��u�Kvᒧ�+K�2�[{7�� ��U3Jk�g�����hB���.~ ���Mz�5�1��%��fG��t��7�6��F��U���?���1H��{M�m��@�s�@����A}X��Mt��Չ0=�>��+�t����R�&�a��s~�wt��N���M��"���.��4B�$M�,$B���v2��h��LVgx�g�L�v,.K�u���ZN�����[�X��y dڟ�eX�e�V63 �ll��W��-�ON�=(����BL�J��j:e��r���	� /-\A$�	0a��z�R���&�-Tɰ$KǳR!�Î�ʿA�|�z�\$�`g����汴(��� �O�'6�n)�(]B���yS
�T��P� 1�eG��4E"�O�K��ZX��
��n�̰rӓX��|{aZL����Y�)m�Ղd�&����B���:��TD'J&����b�bϢG�@�WP���ך�E��q�,7�«V\퓈8I
��/YXDEw���W �8�
�="������M��BЖ+��P�^����mso*�r�u��ȖQ��*�����W� �d
�"K��3�2��q�L ԰
/Ѓ��,ȩ��*�.���u\�����4z�չu��:��^�j]�f�3zp�2B�j9�!�ғw�a�}"_)���f�<G�`�62�o�T���Jh�f��۹�(w�t���
���N<��n��E"T ���e��l^�S�HO���V&��ڝ��3ua���l�tJ�'`� �}1��n��yS�㠁����j����M G��O\j^Gj+�p�n����P&�l�
����u�̌�us��6Ṇ���Z�0�TJ�I�?m�W�b��C����I�&�H���'�?V��{����V���z1��`3��c^�Vyʊw]���W4�H��<��1ɨ�_��j9���3�>��D���R�X ;�6eN�yT��
D�b�dM(�)M~�TN�q����:W�i�tc�'jw�Y��P�U�o��s�[Y���ob�S�K��̒(:��Hz�"Q#D�8j�2Yl�[b�e5�aM����l�.`8�ŉ �>��{o+��.��5Y����"�=��[ �H��ʭ}��""7���Ŏ4����6
��*�J,U2jYk+)#��TX�df��m�vV� 2d;�m����4.�܇r�;���X�c�s����R��4"f�<�c��V:�y�o��Kv��y��p�ѯ�?ߠ@O�
�;�OjU�2-`c�A�MuV*Y���DZ
8&*>�����/���R��*տH|���p`&;�2wh�2;�ؾ���w3x4B�т���_7�쥁,H���2��$�0���T;�����o�xD��]�y�`yp5%����o�Ʃ�P����	���a(�*۳�i΁��wjo�õz��!��3՘-��
������������b���={�.C<��j3�9�����#UOF���^rb�ie���% ���Wћ5:�n()��%��`�1B�:����,xїG!T�h��-�2U�6���y�P�\���>�4�F�yP�Lmd�z��c[�m�����������ͩ޶�����Yb
��E1���,�(�T�W���+���r���!r�dSv�R�:��.mEM�]j:֘-B�̀����_o���f2���@�x9��) V�;��q3�@Rr`�j�|�.Xw[����wR�+�3�I���s �6�5�M��H�S�G�X:���A�c2�Z��A���tK�V�@%aR���laL�~�
O�����{ !
$5������J��H_���>�1�������;���&�t���b]���~[\}~ͬ�GQ��-�"%>�ǣY&���j3OnZ��u8�]LJ�b�����lO0��	_�4q��x&ShYGlZ2���*Bb�V���w��8L�)ο}��_Qj�B[!�6?���j+t	a6ho�y]ٜ����WҞ����Nz�0�S��gc�~�:�X���ag��a��8&}��c�4�M����H}c�ѿ��n�M�V�H֕]d���p��f��� �4h+�V��J{@y�L�Q�=��l<�z@�������Zo�CZF�a�_�R7���i�{��hAC51�+�D(bq�k =a!�#J\��m}�K��h���r��C�^ Q��s�-��B�bo~�?Po��|�+&���h�\O��5=�"�kO��d�~�SIggQ3+ѱy\9�iU�-�@����� c�_3-�}f�s\s�8��5TZ2R�Ӽ֒뱢�6ʆ��~"V=r5�HT�\L� '�B]d���a&��O�ěd�)h���z�7�L؈����r�NƦ�@ h��w�_ݐ;q���zn)0�s9���'�n�15�&��y�I�;B��]�5���m�%f�t_�*���)�RY(���G/A�x�=�|s�^�L����6
�h쒪�`ƐX�V����}�U��MXE[ͱ�ƍ�#����L�$F`���KFR����X.��_��C�O��{M6�������ǘ��j��^����Oia�_bX�/��%D�t'7�n��]_yp���U�D-I���]�J
$�o��]���[ָ� ��@��<�N�ߎ5D*i$��}A�5��Y���zf�H4���t��L/2���d��Ht�t_[�~(�z)����k�d��+�9���.��)?+Њ����i�9�ER[X41�����4�荑�+]!�jv��j����!����Q�	>A~b�\�)�jܘ�W�Y���ڑ]�����m��D���Do:�}۟�r�P�НV�G�G��,�r����ψu�.�rEɮ�L?E�ݦ����\�i��z� ��I�A)ƚh�dz�e�!�N�ힿ�$���u��cd�$d�$��;xE�nڞ&��lXp�`��?>W`����D&����1/��(\h1^����ia�}$����j6=�أ��(l���b�\�k�'{���[�
�a�J����;��ƻ6�.�VI"��K����>N�j����9��6Vj)�GS<֦S&�����w�� &H҇�k���	a����WR�R�S�*6���`���U��EXyV�"X�hV`n4�rR7�Y��Td���i���=SS3pȾg~��Xߣ���*mMrsJ�¸�վ�'���&���E��@�߿�W
��9CI�pVf�t�Z
a���I�L�c�\�$8&�rn٠��������躧�_�kk0��K��9#L�c��sh^�W��Q^ �
0�2T��lf����O=���(��=�ԾҸ_��5�b��NLqc/r�|���`+���\�cd�W��f���0"��ϺO�ǺW�L����{d
ъ0 !!}�ZK�[
�J�,���a�Oi�чǟ5����;�B��W��K�dz��}jۛL���'ml��n꣼y��@��t{'��ȟ-�Bg��D�]^:Չ��Y3vX|1���;<�"lj+pn*H�N��$����؁��jN`��S��=m�Q�Z�A�(_��68���@`��5��9+�o^C&�ʧ�vd���6s�)3<��$�`��
�g�4F��|{���>"�wf1�&�ԋ��+�ak�Й��u�7����=?�|m�P�1t|�ߴ�K<��t�9�(��/��������K!��͚�~"���Z��� �P�D��E���jZY��7Ļf��y��x�V�8�S]>%��̪���D@�w@EX�M�^����2!�m������f�R�c�R�W����Dh$�9�E/���u���'��p����I��/�|ةJ$����Rڞ�� ��>�ZY�iD_ߖ_'�M�B,�F���?��`:�2G��7�ݫ��W���S;����,ݓ�%}��M�{�|��@��Z�8��A	$�ZdQ��r����%*ۂ�a�>����=����-J2Xl�jB�l}�+l����W���5ͯ�}�q��t�[),4q}'j���Q�7qյ��UM��`xm�mh5�GA����B��G����a�<U��������:�&�1b���&���W[�'3Ye_�Y ��l�����M�o|�����������l4�Y8I�肙�*C�n\鉹G�"+ӗT	�����j�n�:�]ҟy��Ae쫮�c�k�ϙ��>f�f����~C���ÂM5@�C!S�́_�Fy�4^�d�R���OȾ��\S��%p��6����33Z�wf18��X.:��5G[x�a�����zA/��-58�_T�K��&�?��2��P�- OG��h���������@����	�w���$�v�L�$|C.t�x�B/�����KO����M�*,`D��Ф[N��.n����~5z}TG��NU9A��熘���x�� Y[����� ��Jj��� �	m�՟1An�t�r�e^�ys���6S\��qj]��˔m�QcB)s�§���>*��������oL��suk'2Zt��B���������t��qX{�k���m}t��Y��ٰ�Is�Y�P�~pH.ۋQ�xj�2�w:K���g�
���0�(�U�ֶ�!~
��$B� ^4��kb�u��e'|��Xb궊�$�c�;�!,<x�P��b�O�M�R����-�c�V��2��j���@^^�.A�b �W���/,z���m��!�����̨���#`�z�d2Ŵa&&VA���<�P5�!?�m,���"&�����v%����ÄՈP���y��3��y�"������H�y� �����(4��I-�t��K������~/��1� vY���AnWgRb��|�`��_=h_0\�#r_^��t�g�G�W�J��c&7�+x5�Erڭ���!ASg''=�^��
`��!����_�DnG�]5�b�ECt��ם���~R��~��
�2�Y 8�&s�0�H���-(B�Ӱ���oӌ�C?�$�h�}Wn
[& .w���q�@�x� �̟,��ρ�>��q�ihy�9�c�W�ت�F���	�]N�]B��c&l[�dO��\�b�fd,?�ry^�s�G�z��:�WRHJ��>-�ߪ!�(��*6��V�@�(���Y#*>���>�x���#�����U��`�� y�XZ�ס\I+(hd�>��ʟ�(�e"��a�ԙ�=�ѳ$E���q����$n}��a��]�X[i ��x��&Z�Lb�՟|�2f�:�t<��S(��c�8�*�^����Y��#e~��j9�?UӴ�&B��J{E?��{4��\����C?�:���(	#`i�s�@p	��vv5��aQ�,3�1���������\�n��]+�O�Tt�Uq��P�)��1���g[Z�r���K�GLBz�CA=��(�����y��iw���ܣ��Ș�	�<G�;Ȱ	��?��^�&�֐M���5�ӆ�B02R�};�̕
���V��^N73n�{��J�T{���Н��0��0�hx�'�=��4���N(����i�P��aS�_��9h��&cr@�LW6��_wV����۫�!��H@��wx��]� ��Gq6�6��z�e����SK,��j1@]Fi�2�W[�%~�+��C}7��X�亥����Y�����HSi�X�� ���LM���Ք�ο�^���b�5������G{����v����Ya@ĺ��9�'B�����0�'>��̕.,���'����*�3׳�t�Eo'`�؂�/��R�r����\%�Z�`D�C;kt��9�v�#����G{uz�y�kI~����в���)�`/5��eDߏ�U#ES."�J.(����׻�S\�B$.d���Mژ$D�$
g-z�l��&�'����S��n��̪�5�	��exN.
�Z���Ԏ�rȁ���KqJI#�b�B�a�r����������h�=W�m�UsTb����e��'����%�M��q ��n8I>�1#��<��b2�~u����߮_��F������x&�QVg,���{�iy�&��=�.��q�[B��(��N8s�\��p) �^�� ~�C����痝��,�\�{x������⏩he�)8��N�՞�X���*�J/x�P���=#��t��d� &�B����wa�#�TI�$�CތJ������Ud�7��^l�-"Ǜ���4�嘏Ϫ��jW�^6�ޅ���kW�+�o<y��LU�bԾ'Ze�}ec{��8���Z��!-׹'C< ؾf�I�����[��9;v�2���ze�:Z-L�@��8�����- d��u�����<�g��z���uσ�6��.���цW��
}��k_*vQ�^xlM��ӽn��ekr��!��=+,��Da�6�h����d�/ e��X�(/�
`C��a2X�ELu�����s��뽗�Hx��t��&C�j.ϖ�K�Z�L�-1��4}��j����T�6L, �r��|�i?�aM<��M{|�YO[V�Eڃ�T���
�DO�P�q ����#ӂ��-2/v�n<��_fS����g>m�C#m�2Mp�Km[y ����CG=��䋴�H���$�m���ro7&�َ�J�A��1F����x�'gp���$������ ��� ������U�W��F��8��z��T'����!.�F_��J���lWy8#&��Ş�E�Y��gcWe�Z��s����~���ÃT`�Y����іocw׺GU�;�:�*�NQ� XP��K%��>:�E��7�8:���$��܏5C��x�$�L����}#/�P&j������ܒ/p����8�GE��K%�: ��P�S��}T�	�/B�8���\	�Qy8�Y�X��.�]�|�*t�@�p�<��?׽%����	�'��t~y�`��T��>��(�.4U��]��BJ�M+�\��]���ϝE�/�,�Buҽ�J������/J�+(��M�B��N ���{��	8���Ơ�z"x÷��s2�v��JX0���mb�f;U3�@|(B�oυr���DG���]L���D~�s�F~S�pΜl�0����J|#4�7���J��ߊJ]� ��B7�b��]*eo/L��9��g1��n���Ae�M_��m�Hfj�8_5�5e�=���4A+mg��x�d�x��d��j,09��(O�_|�Tc��6V�lƩ]iv��xx���W"R�7�6�7�.�~y��;g�N8DQy�
�s�mg~y$��fɄ�WL�e@� �L�$G;�95�VA�l�	�=r៰�8�/��0��?�-w�36�A$'Z�ɨw�J)��x���9,>t+o������	h)GBj:��ъ�{p��B�P:�%>jn�^֎M c�<��x�Nϵlg̊w5	B��͍�˩��A�~������g�nA�FG�	��=�}i��f�m���W�(��9�K��������r��ޥ{�Y,������q��+	�z�aQ'���[��0�`�2��p^mH�A�m+���� N�,L�
�����4~����~��V�e�b>��,P��u��6�����c��uw��d/`v�6'��+f<+�pd���>��kf���u�*۞ѽ�G[ܘ���
U�X/Y{ruGeNņ���q�	��jV����h6]#�cR�*S��;7���˶D�cH�K�=��T�g�����/��é���`-P᰽�_C���}�gF$k@o?}M�9YJ���Z�����Eu 4�K��i~[n��}�]m�����*%�b�� ���A��Fв^�ʱw8�f�V8��]�F��ODõf69��fk�xݟA����h��xi*G8o�ѩ/�������*�^�$�:�&f@���d.Z|L��PGйݏq�����W��;j)q��8����hI�uId��; 9��,Py1��t;�!����>fZ��(���P��H����j��}�a��A������sD=�j�^��e�K�U~>S	V��r}<��7��<�[�<��ث��BH^
�h;���� �'�jD-��-	"k_�F��t��BI ���M�������=}Ii�ʀՂ�
�|��L7���Ae.v�y	��Ya渃�ȏD?ʷ	GR�p��X��;&3�(��W�G��9����o���
ӌJ���K�ִ�`��-tS�F#C.��!���t�s�FTv�{bpO����O(�!]�b!���Wb�n ܌���+�W�N0�u���q��z������\Kx(�'�A��<��*�n�/�_�(�;��xK��O<�)���'{�����W)�v�e�Px�E�EN���6�F`ư�C�h�u�s�iM��Z�Ž�{7/�x�Yy�scU����ٽ�t.��rR�Y�h8��'+I}��ֈ��­�D�A�͢Tl,�A���t��<�"�l��Ō��~i{y���i��s�-��{^t[��^��ۅ�hz���U�,�@_�ٸ��-)v�-��oXz��^x�Ɯ|��$���TE��9�;Gh�S1NRp�5;�j�ю��#c���K�9�|�S�^��\IL䚩Mdsuu�=��ej�C��[����)�c�r1۷�aZz�h���]�#�(��;��o�m<�Yy��4��R�1
��9j?��'�#�Wg�+���	���ԡ ��۪w�jI����_���-جXR�rZ� ��XMb����|���xO�7H�8�y��J�V�24J)|tw����n�j��I�����)�K�<$4\j xmB$Um�� g��R��D�!C���;B���K�/�"�տD���Tؤm}�]�:& =��B�="T��,Ͽٜ�����0���Z�J����B�^yZ���ͫ�Qoݷ2��`\u&�S��3a�K�w�>6�|�5$+g�a�=��R�`���J�ސܸ;�����a����뙝�� ���I]j��e���ߕDq/ɚՃI(����|v�w�I���L�C�cx�IA����9x�8i5�w� �u��ȡ)�n,��arַ��J�t�:�}��M�oyP6
ꮕ0ĹB	U/f>YY�n� 
o�P�ig�5�x�N�n4��yo�
Kߊ���i�,�����"J� ��Z��2a���2p�l��eU��-��Ś�Q8�ϫ�;�__5E��A��#X���a����!��{�۸BeI�)*�mX��!Uh��2�EҖG�K�����j��&��eY��{,}�f�f3���.&
��9C`/��t�8+��W8C0>��f�+�{��A�j��F��%�0\������SUH�Ф�a�	������U���0G�P��(����BZ�S0��zW&��a� ;">��x�L�uS/�޲�H�Տ���Oc-p�аU3�2�g:��gI�,���^��a0}Ԥ�~ o\} 5�P)upa0r�A����t���v�4}RZ "�VBJC�.���^yxD&`���@���8�,���q:�M{7�������}U�n#��1��Z��K��t�dW�E��|�3�}�SʐY�1�� V�i
�4�̓@$��kha��7F3�����tY(GRI�.����`b��=
s������I�o�+��g[/���?�P ͦ�������Yk�j�Sc���D���g>�o83(�y89H�p�9'�d�b����b��`�3x�l@��>���g(3��r�CDE�������5�C�3le�`�M#��8�O
&���z�V��N�f��D�`���[b:�)O+���e^ppJ����.��n��G�!hğr��̚	G����N%ȣN_�h��f��?�	e�<�{2(�q����]�0�՚j�X퀽�O�&���
�0�6+n�&���Ӑ�Fd9����]�h7ˎ�<����&��+v�cdwJ~,��������������M�N��ɭa��A#@�t���`2��'2�$�)xi)��)�S)��ohUh�:<c���IQ��o[�t*y�m�5*��K��E�a0;H�"��d,(x=B?ϯ�/��'h��ʴ��cg۴�馻�LD�b#�Vt��v�F1�,��.�H}8'b���劏�����4�~�#�
��|�,��fW����2���s�Eu=�v`��>C�q�*�{�qHt�B�M�KL��M:	%M����]�� ��<��k�r�4Mu����K�R$�t�R.%y�J0U���D)��'_��W��v��`�0����~���F���Mމh�_���\7(#��<��{����&����Ŭ:����Y�@�� P� +^�yi�{���l�q=�-fZ�q���l~r�!Fz�|��C��* �?�ں�#�` g�hv崎���cקu(�߭-��; H~x1�`!��C�-6�\�%Y�:V���*�g��),���k��Dc!�Q�b�j���~�8��ACi-�$/�6�Gܭ�Jc*�s��,����,;���gK����
B;ZE������ �c����a\P+�������e5c^���0�P�+�È���dwx;��C�6N0��=�B�l���ʳ{����dUuKr�W��Q;u�3�\��f@��#D��(������U�ή���́F�Ϟ���bN�
�V.��h�����R�5Lj��J���NYA�`�Z��ջ]��l��f&�IJ?�b��+�č�!�kҩ�)��%w�>P�},T�G���w"��8O:ͼ��Z'Ğ��T����EY$�F��v��G��:s�tbG�?I�ʓ�jqg��75�:د��*[���1�5��8v�m�l����.	?����7��iv/h�)�Y�)����Ɨ*�|�YY��nK��Dz�`npQ_��5&v��@�\���ܶQ��2ڢl�}�;R�V�#E<RR���;�H�{Dh	�Z�ftm�?Y6���[��Z6�M�2����\�T�6e���	�$���1	G-C�'�%�t��UƩ�J�m��>�H��tp`4}��s'q�� u�D��R��b�+p����L�JB
���j0�L��ʟ�V�����N��P7R��M�F3��>���{����R ��Ă��5~�#�<rh)hMe��v�X�YW�8e��ű?�-�v�q��b����+�K��[�9�m\��l���MS�*9���
y�o�M#�	oǍv=����&2i�Yb/�X_X�s�Sz��{?M�C�e�'j;��y��KZ�)�Fգ���Dl5���,�����0T}��t*��N[����FAY�ߗ$C�����o�4��q&�h�	^��ُK cJ#=�,o�F�0&6��h��c_��g�|�����:�(͑�B�B�� �x,+�*�|��w}�޲����"e61�e0��I��]ޫp�P�5�����牐�)`��"z���l��-0@^)���F�f'�R�m���}����{I�� 8E��>)S�A~N�S��2�"Q��sc`
?`ŤG�I|��wʥ�e7ʂ��H�F��Ѿy�2�32�)uI �U��o�y�K��,0��z���D�n���ِ4�^_::�����)&��%���l��������w�Q4�l��ӳK��?Ɗ�J_����Z9�B�Y��1������
�r�F��u�s�"���(ˤ��aT��[g6������ZW~9��^S/{�8PI���B���צ�x�P)>�J��3����M��M���1�����2N��u?�.���\x��ɦ̀cR�3K/�ީ�C)M�js�[Q�	G�5w�ݠP�q�ѥ]1����ĺ4u���a0�>K�$?a�L�C'p�K��+Uԡ;8��5�
$6�a4hz�ib"cx2���A���#İZǤ��J>Q��B���L`��c%J!u4�&Z^�b��=���]q�-w[,V���4eļ���)s���`�����^J�Gn�e�_�@������G��e��g�d.��[@Q{ʬ*NLn���6%C���1�f	&����O [8�,��>��攃.g��|ɣ�4o�x>T�Z��!�*�J����Ӭp��R6�xW���^�x~�~����A�My�tk���1j��;��$PB�v5��� ��T�Oma���=��hx��gBP92�_)��C�`�e۹CU)K<��[�?�^��Yk���?�-��Ի�bL��ob��ؓ$����B��E������g��u�U���-3g�YD��.D��yc�����N��V���(�	��|A�ॢ�p�m
��'_)�L��q���g�M�ܹ&��T� +��
�0�7;L\oE#��Ht4�>���[�i��.���K�<ǈ&k���N7��.>}�)�_��,��*"/6{"��u
�'F^#|�e�8����Є�Q����C�2���,n'|�f���J�V�&ge�1��6X0�q:�qx΀��T�.���/^ґc��觱B\�U�ن�����C����CsS�"�qe\_
'U_[�s�n�)�W�҅OŏݱE�d����.m��b�␷��IJ��O6�'�H ��X��N�C�WA�z^'��͑��G.����7�};��"�OR�>oN�~��VN�ς��VC�Qxņ�O(��R�L�<���ھq��Ϡr:q�H��?(�� <e�A$�ۚ��TA���	�ߺ�R�%�A�2���b��Jʵ�vY�"�4^��:rk���:��	�³;B̒uQ�[�\=шL��W[����v��H�;��#��!#t��J��E}+!�	�LqtP��<���%g�7��5M�T�y�|�	踥i��aJ��F�{�7��\�b�xe���<�����N!�YS%�M�׵b�-��z�B#��DŊs�BJQ�>��
���W�"�ԗ!L������<�.�a����Ѹo>���������V�9�ռP�VY��#���]x;.���S��PT�%�k�<N��VI_�e�i[��x6ͷg�O��uݡ�O
�9)���*[�}p�����NB܃�&�hs|��~�/�H����	1+��Ŕ�������Q�:�x{X�ʟ�ł/��}��9�hd��U׳��pu~:��_t�b��}�k�F�Y�kN�FIЮ���#��q�3���YVU���D�cT�Z���se݀w�еHbA<�k` �X����^�T'�.�����h�P�C'�1=P) "��y�1��>��o��QU��@j��+l���+܀W�&v�"VJ*��%��F�,T\�=s�}�֯52g��� �r��B���p<(�.xzm�Yk,a�cP�����q��;�d�9���m�n�Ө�;J�G|^k�w/p�k��{��t���c_���;��M�����R[*���L��xz5B4JY�&ƴ���;y�.2�	^,:]��j���/΄?H���@Ģ�,�l�N����f�6����)�A�-ý�5������A�ܞ�!B�A�ط	4�֨��U�xG@�vm�|��B�~6�%��@�^w"ͬX!�������( c�hZ���u�L\fI~"}ކ��v``�%������p=�*�X�:��!
q�t@
���ޝ�u&�f%n�΍-�A+�����v8��OV��|1���Y7+ߞ�c�;y�_'l�P�����0 �,:x^���гҷ ���_�d6=��'Ϥ�Wk.k�6�8>��b���y��F���Sm��d�+1r`Bm�T]��ʡ�3����$�pgU�?wÇCy(Xz̦�\t���G��&��9)V�d�y%=:�Q��y�x�E���/ł`t+el�O�S_^�	uw���vx"�b�vI>�{B�7����!y��A>��Z�[F�R� ��c�]f�j�A�$u�����Y'���I-Ǻ��!����J�~D��Jo�6[����[��v�����G4�<�w3�X��o%�|T���dfX��@«��X��+�ѧP�~̟�1��MI않��.�T��	9�ݙ�/������7��
h�R4O�VZBm�>3��g,eI���q���S3s���q ��W��=��V�K��P-�?��Y8l�@T��!y�0\��Ud�Y��6k�������	��
�(g�0���ŜҼ]S�:N�m\ �=��G4�	 �t�S�"0Sh�x����8v�e	�w�0p�1�\��� Ü������eS���r��īS���Gn�����[���
�ܯU�R"e8�ר�]�3W�?�0z��.C B����Z�%CS���)���F�$_�rc��Z���Zb:KGφs���o��C_��4�L�.�B�2g�����v|M��j� ���2�]d&�<�T��2�=��9h���2k�g��g@80t���#��s�K�Y�ϓ�a� :Ĝ-���^~D7�!��GGfۄ]֚	�$����M����)X/|���et>�Ā��j3�f����Q]�}�#�E����g���䇰���	���SEr'����,�+F�j�JS��zj6c�@ӄ�Iq��B���L���4N��y���<?��O����ވ^\r����V ��\t�퀜����$�D�y�Ֆ/KU8�A�=Aܷl�S����y����C�3�J鱮y�P�g�(�oX��Yd<.��>�����T��A��P��>b��MB�Ę|���S>�!��af��~��!��j,�?+6n͵}f'�h����g.�#C�rbL�L=�GՃh�]:�F髆{��?l~�%\�yx��z��;��KY�;G�q��v��כO�lo.f��J-����jκA�"6EoZ����3���X>6��l�P��FD��%�֜lUO̚x��p̙!�27��*.>,�U�P��:���+��U��W�#ͽ�Ek����j�l<�[���^D���h�Aa�g<��($۰@�N>�{-�®���qQ��H�9A64&��Ov�iۚ��?޳�M�gWu֕���m�f��Jt�l;�,p/D��Z�SF�F�,�N)@@XI�?|����{d�8�~r%�����e���;](�xP\��I[��͚u@ln�M��,�h{ǘ)��`�"Ɏ]^J l{�\���*,m.�Ωr��َ�&x��;3	�QW 2ҌA���Z/�Ӕ\eK�:�&����@��QP�;�*�_�e6��8�������x�@�V.�Ȁ�Ԍ%�սV���l`̀kצǿ�G3��8�szz�W�j�|��k7���B4���B"?l���G��;���Tu�N��
��O����� 1nkv�n�*pY�
��K�[*k9Qۥ�{!�k�w�T M��k&Cң1P��ge9^�Szߓ�Phz�]PPN�M9���.$�Ѷ`��;wǄ��M��mwވ:�>��'�<ҿfL���_�$Q�G
 �5LU�[� �$��ዉ0k	�5YM]�N��ut��8��V��f�r�02� g�b�t���C�� ���K�=�8:���=G�?6��v+���q�%#(%�V0�q�ʵ�>1i;�e��#8�IFm�1��ED�K:��G�Fx�*;!�3��#@�:�.�/n:���$U�D�iw%��K8�2`�-;)+�k�8!�N�Ą�vf≶�a�I���	)�X>�ʻC<�{�<߂��[QL�E����S:��JQ�Q$�6%'3�Ô��9�h�~;�~�4���%�5Q� $��["�^KDKKV�G�5X��$�ܰ*g!2�V�*�O�	�+��,P�k�p�I�V0��|�_ϥJP|h]9
������^��A�`wɊ�hҊ+�R�^&*+`�9�j&A�7�y+�����ǃ��<�V��/9�@Z�ԓ��H:��C�9uce*<au%\�7�nɁ�ϯ[5�!k"o�k�K���v���	���TD����Y�Jw��R}㼒�Z�T�	��B���`uVi[*%����Z���� �@5������t�a5�\�mK�K<i�k�>2�tХb��]G�A|lV���T$�ށ9�a(g�@rZ��!"q㜋Ҕ��a���R1�K��O�n�,��^�*2k���o�,���g[~���.eUc�h�m���8�t�~�iUn��%�+9ӣ����x1��=�����g �<g�~��ք�^gq�� ����5 �0^��]R�s�{{<u-_�m��>��L�ӝ��^m�Sڏ���fE(0Þr=��l�_Ý2�{e 
[:�ܶ�+��6]�b���S�CB���%�^*�Q��)B�_�I₧c��}1����y��W��[Ą�nn����K��T��Ǜ���d�L.��ٓ]:o����� ����t��IY5�-k���/�.a���~"
.���$���44�����?F�Ȩ�<�����a�濕/݄RN[֎�z�&n�v<��$�A����t�%X�pO��xP�%��a'�D�\j���B9��[��ġt{�|2��ç-<���i��6��s��]{��ƃT����O��]N6�"��p�q�J+��eK��iND��m��no�#��a���<rԩ.9(����z����,���G���{�/n�U`c��+�/� ݻ\���r�^�u*/�p���x�U=!��WG�g���3l`e�hf|�Hx�&�t��^Oo����x���rZvw�����[ʂޅN��L��S�����ż"�d�M���M���7b��J����/w�K�^؅�w��������5"����+���S6��J����
hm�!���|���k��z���v�C(�36��̽���ၲe���v��t�=�!���?�12
_�X�ΰ'��}���<BR�z���H�Txl��7���Kd�eV�������i�Nd���0�[����@��������@q5N����!�hpQ��RMU��Ŗ=2��UHc�b�p�eαƂ-5��W �H�e-r�S�>u�S��G9M?`��>���h_j�����	a�$m.+��H-��p��X��eh��"�����o͏ɉ�Yx�_��xÎdw�'�ƈ������f��'��[�E�Ft�+�d��V��N5���▆���摀}4ۅt��$L:\�ć��2�bl����Z���z6���~��H��E�!��9^��}:�4��1^:��p���.V��9YH��t�H��9$�0�em9,����[�#���l�g�6��./��M�m�/}Ȟ#!�i�(�N��	f$+�ډ�|SO	\��6`}����m�Zſ�od{w}�q_n�Ƈz�~:�K�bg��n��?\�G-�q}��z6�R�k����F1�fry\����˸�g����O�]��y{Q��+������&M����&�Ж�L*F߷�ߣcN�T�J Ī��k5(1fs�l��'cbw�����c���|0v� `!�7�t�n�c���u�ž�,�Eʙ톍0��SqU{y���v졊�D��mqu;0G"n��s�\rNMŉ)��^xM`��w�*����Pm��@B�*H��O!���;��s�Ej9�` ,�"�=Ŧǭ�Х7��}�֜��n���v����@bS^x�Z��_2h�3O�t��B$�1�c�W�hA>�ո� ����N#�yZ��{��R�~�|6�C�n��|���g�&���PƠ��3E�.�F?1��)L�*�?�I�ߑ�+p�''+�]��$�"�c�V��(�ԯ�e�Ԁpk����LbF{b堅�z�f���ahYFĮYC�zH�N72�O{�,S�Yb�JP[0qš�n�3��-͠˚o��[�oV[ \��3%�v�v��^������լ��`�t��BA7I0�>r�f��M{T&� q �!,'װ�WjF�C�/"�^��JumI���3'iw$�e^��6`�[`����d?v*��A����q�
�GgS�W:�`��:Dk,�3J!����V�f,2�ۂ+H5p���O�Y�
����҉��:柳��d/��xy��]���@��yNJ�N��.ϟ���5�-��;�iZ�#2�.�^V�����0�n�ŗ␀2��9���ᑡ��=���]:p��IQ��̲��[g����i���r�ܣ'(LG8��б�
e>*�J��C�	j����K��HB08bגM*��t��ݵ��bi�����p�=�J�a��d�,��w��+,>n��&��눧}~��YZ��J3=�w� Wy���k���H�zռv�L6Yu���)����[��b�s�1 {�ԲS���IN<ƻZn�����i7z+S"+�b�F�]t.qȳ�TfU�tc	�"H�(��e
8��;�Dڴ/�=�t���J|��-;b���U������9.P����#8�L�hgR�/%�۩�0�O|G<��Px�Hu��� �UM�YG��@Ó|�����a~���B ��UΚ��� 
=�DL�῅�ɝ��D��!��$��7 l��_�y����r��^x���%_�8�������9G�6��(#:��>��pz��.BV�O�c�B�|M|�^��,��8�נ(p˭c&���	L�f	N�F�!��2�2�I�M�)[[<���K?�뎽3��Gԓa<	��r�X`�&�h|�� �θ�tX���N���o%_ײP�n��8?�b�h&�2.������ha�����4mB���m��N���z��@�RB@�83u����	��?�������(6��4�^%_�ABt���������@��v��/��w3<_��ㄓ1�"�{�9����B��-�B�M����*������h�l�@�����w~�tr����~�"0'#pE����]�3�;_�{��-A�R���r�u��%�R���B��^��P*C� Sg?���ތ{���ݴԢi(+��YoT�}�%.x�D}�H�B���:kSl�N9���ԍFFR��f�I�DoK��T�m��j�<ؿw� S��[�ćH9��8@�SiHoyBx[�=��l�%��\Ƅ��K���j���L�ͫ\�_8���p'��c;nÉ����i�=L�yl@�#��P^�6uo��� N׮�n����q�[����$�z ��Ocuam@+��bQއ
�ˣ!���u�!��QÑ	~�Cܦ�|��� ���/w���rS8�j,���ǚ"3�H��r*��z|3|dB�v	���˼�q�~�تє���y�]97�Z�oy*6~>�-�[�^�5�,�z}�Z��B�*7�#l	�=�!��Y��H
�n��D���Qe~����9����JH���/���ƛ�=bGP�zJ��ܷg^�5�ٷ~v�m��vAݙ�����f�4� ����NOޟ�M�-�_'a�ְP�8g=�1'�Ф]�R��IRdJoI����@JEkJ1�X�-"�%<���@��g�qO}_)�tm�ӱs:�*,�N�<�J�O�\Hh�����J�2�!� /�V�iRh�	����M�
Ǚ��ߩYմ`�-�Ԝ���f[~?�u �x��?��\j]��c7�ὅ�����*+��.���K:�2.���7ZHȱ����kȰ3�8O����u>֖ԍ[w `�W���B��/�P��l�Q�N��=/��.�6���?Y�Fq���Ї���5JFs�	��dM�tY�]����ɒ6	��C�t��U� �R���3CmTL�*�p�2�����&��݀}������g>u��b���L~��=\�Q�x��+�
�!����Gsh�:�#&�Ɔf��~�9��,���9���Ї�A�uh�g�ԝ����墭��Q73�g�K?�ÿ���!���� �D���հ�9�/@<��8��~J�^�XR9�_t��L�}��[���2P̤��WS:1,߁P�@�܄9؀�0�g�	�ܠR��;؋;��`:���z�?���^Ҧ�p��5��+ "�V7��K�6KTL���P_���Է�6m�����P�US��q�ocZzd��P&��gL'G�Me������NpX	 9��O_��	h�_ǌ7����Æ�U�}�B���:y��'�R�f�������?��6�s6�-�b��W>O���䀀�(�ZYܷ2�y>VE<�BnYEA�Q$^���`갱#� 6���P�lϝ�ٰ�_F��6����&J�z��I�;^�d���� �zȭ�Y~i�M��ѴP9Xw73��%@!~$9���XWi��� �,��j��D�A�q,�g���1�K�Ve���&�D;���r{��Ubq���
�.`�_����Ӄ�9�Hs9��bLSo���UA��1��ܔ�2	O؟����@��q� `{��OШ,K�̏g�D&*������h<���\8[�N��w�$�^��7dS|iU�"1+�R�9Zk�Q����0vl jȏ���l3�J9����o�tx|��D���#�~�����̤����}�'��ֈ@���2�Nr�S)'��L^o&�\1,]'l�Ό�4�lΤ���z����)�R����N7ʼ�y�Pg�J���PΊ��vٰ@YX=*U���m|QjF���~^��O^��ue�tݽY���3���T5�x���h�Lk��$���*��a�/\�3�O0�ܚE=����,g�-�~k�ն��}դ��5�hZ͝��v��Ԓ��.�T>xG���W'��DD'���9u���Ij���):R���A23�te�7�z�q��%�pw�:�3��2��v�C[�w��Y/v�\��oR@^��
R�2Ou*!wĵ����Q��t�urm�\�MR�n�>���W	�"�D�ܞ/���]��}�Ϧy�%�AcN��f���5oɺ��ߧV8_��T�f�<�L%갌!�<]�q���=V��L��˹��[�4��;d��<�-���,�,SB�BF���6�1

��#O	t���b�`ID*`�u��0P|EFI*���mB�/���,�������35NX�ómZP)h��X�Q�1�3e�`�4{�0��zG�
�6��g�?yͣ�o��>,jRa����v�F����"��f@"�C��2}[xo[�H4:����E�5��`F/,̬|y�΅:�G�$9���ģ@3؅���'caA���-���F6��_���؃�#�����d��]��~Ю���8~�G<�F�=g�����{���a��!���'�3r�!�R�:�c�N7�N�9�D
�����2�.o�ov�܍.��צ��<:������AB��g����d���:@#�Jp��{n6�Q���[\���i�G#�U�U2����IvTH��L�'�H9��}��T�D��zuq
�i�\(b`?��+q_7'�@Jǧk*��p��Z��K5e0�.���ӻ"%��d���
j������p��2Z⡯�ވ��Q��]���@V��*��_\����"e~C�`���k�&y����N��-�N%=C�#?��i.�L��^���#�>eV��D�uU+������|,żI�����k��Y%�@�O�}��!̀������ϰ�J� �� p	Vy@=p��l�*��"� ��<Gg3��^���Hpsoʈ#�(�(�̯�����ݑ[M�,�(�ds3��|L��7LH�����vm���iȜ��t�"ޫ(�9��I`�'�k7�{��n�VD�:7�k �{M��TI�� ��l.�k^�+$�mP�!,බ�&z�^��G�P�}�v�o6�5_���	�Kd$��_2^x��Lo�.��!b�x��� ~�A�M�����=�����4�'.1�?#c`�Q��	��*�s�99�^�)4��e���U��3!�g"O8��(�v�#���7�L!��� �J�=����̅�+dC]j�,�$��!��>��{=F���M�G�֐�[,�6�l�i]�a�#c�]�`��+�_��Ax�S��|��Wiv��݅���< O	40�u�:ͯO�����<�l�>���©���76�7�ٴ�sUo��-y�mԣ<dp��K�b�vc�܀t��1+f��z�b;Ɓ��99��ze�r@Q�/#T:���v'-�Nt��\���A��w�u� e68�֧Hp�o����)m�ɕ�P�'�`PP���l$		`����e�l��]1'�U�|o�(��%J>�%�ך=E|�F�'�oD[T��s���]���*����8��$J+����B:�M͈�vR�my�VƁ`�����ё`_f?��t#������Υ�^Y=C�4#p5�<LF�E���ϕ±�{���&��O4Ԇ�2[ ��ǪVR폛q^7��tR�û�؆T^Ϧhwxp��Sd����,���M�P�6��2�P�*����.%��-Q�=yy�n�{J�f�D]y�ÎƗ��J��GБ'R]i����9��$�8(ʶ�?[�M��m������2g|�i>�!�Y�����l�~�U%���F�o�\g	��BlЧ!�=�Y�;��S�����I4v-?�S`���Uow:rۯ2d�x	�7̳��@V����u�mi���ݴ��p�L<>8rwik�� �.�#������b�����~�[����8���7��rM�.ѕ�31��x��a�*S�zA3��(� ��tR�'(����TC���k�r2ڹ2�/��kH NQ�4Uq�w�:%M�f�3�s�<��;L���Pbo<=<��Ήn�����k�!�r��&!9��0�b�j���0:��e��{�RD��Eݞy�K��˸�.)"��_z׉����wY�c�;�
�	La$��3+��b�
����馢֮ٛ�� �B�q���#s�,����u]��2/���ժ:@'�w/�R��/��X\'�0}��e��*O�o�M��`��WE��̳����k2�=��I>�p��u��ZʡF� �l�/Nh$*���c��,���o�s��_"'_�l�r���&�A6['�Y�Y�m��js��1�)!�����Q�.HO�e�q���&g�t �.:�B��!8���l"c�"3B�(�V~8��TF�Z{(��ZX����@���'�Z���L��SX�iL�eH�}�k�[�?����io3Ez�\3:�,���x�^*�]��V]��'=�<?q���v^�n�H\.���%��E��O��/�]E�	*�r��+[���v��/�s�`�c>��!�k�n�Y6���0�|;"\ҏ�tQ�I��D}I&�p��^����78�]�Mdk l&"�������o�-ü�w�ъP��ҵF�aS�����-08,�65��0�ߦ��ŋj�i�V"��ƶ���Np�&%�;���K-�����Q8�J�-uU�Д�jd�2["��Pm��;�a�+�ĥ}�����g��:�kܕ
����t���Ff�����D���m��$�ʗٽ'O��%��T�l�ʏ�K@"`���L7�?XB���J
�u��~t�{1��;�x+�b\k�OM@����Զ�檥�K�U���������&,��l�!/����
"���6s!G��{\�v���ӶT�RY�\ِA�cÞw+��WoaWO�'����+*T��6ߠԿ�����p�T4|�1�Ld�2�M����\i8���}���7��?(���rO/v26�Ř��ᖌ�����e��	�}c�V�J��r9��$+�!^x���8U+�o�� G�Hξ���3��f`�/��d���F�Զط��8X���3���s�>����G[�B݆����]�"��q�Z#�=����ܒt�F���^�܈��]����؅lEײ�F�����8Z_�E<�"ݓF@3v���:��wD#�'^
�� ��Љ��]�<���t�P���v�Ҏ�	�A�~ ������\���^�_��lׁ�4��?��Y>b�T��.�5�W51zȔ�a�C� �:7�:���%���qX���>X~R�%�nr� ����6�����h"��7�OW��\T��D�%��������ⶶpGB1z�yE1V�;�7�K+��`�	�H*8�&�0~�	���t'$�d]8��Qv��`F����x0.�m��-���v";�u�;I�������Lgo������(����-�Q'`%H~�H�|?����U>V��y&l�1��]6<ʷ��B��4���'������Sy�?r�L~E�GY�ة��� C77�Y�Y�(Y��&X��HJX{V��&z)��2���.�������S>v���\+zF/��x����-�3��A�j�+����dN�T�k ��Fe��j��$?OVp�E���|̳�g�#�:hւDp����vϱ�r�*����nRA�ϱuU� ��O2�~B��jo�|e5�M�~�}��G���pN8F���X9���"�:xQXm1�n=�	CzrD�rXMIs�����u� Leqԩf�U��)̌�"��b���.ؿ�R��a���4&
���}	����$����}�d36E�`@~�#Ơz���M�h)b(]�B6�h�:b��-MJs�!h��6\+��>MO�h9nv��̐�+��۴G0,�c���k�+�/@����h�Ъ�n��gA���@�E�{�s>�}ܒ��-�:���mu!t�����TY�QŀW��
Lr�������iP�H�uBvjb� �tp��I!��I�c�3�P�����֬��GqD��U2)�p�-��vo�<�����c,f�.��M�W;&�x��_j��4g5�t��X��_��J��H��=�?�c�k`���6����Zج����p���:. Z�v�Yu���]��5z��[�L,m
ҙ'M~���o�"�U���Y9H#t�"�+SA:wDɷݵL[vX�,��~ܤdp�>M�-��;�3�To3��#ϢH���������o�3�n�$d�mF��^�[�k`̵j6��Y�G�[گk"�D�޾���3}:�	���}e24L��rڒ��[Z�叛�¼�8�O&�����Oz�S*=�k��?���q��ˤ%B�Lț ׈�V-�K�����z�3LJ��il��2��^��WL_����h�6(#Ӫq�����_�a#�g�Hu��-��=��%�Ĩ��ڳ&�]k!}��n�6��]�6j����+Ĳnf�œ@�Y�������\�yw�59ޛ� ��D��?i
���o�<-�Dګ]���}����M��PL����J�گ5�!a++W����:��1��_�UBF6��)֟��S�W����zlm�>f�����/1�`%�_�2>����_2�R����=�rLq���o�3�� �A|lM@Pғu��"�3�Dc� �Z�k	u%`�����Eoզ9I ѓ��f�#j?��24	�1��R�_��9�+������$��`�z9�xM��`?� �Í����bez�w���ݣL-}YYQ�*�����-tNqo�O���x�Z}H����6��K��6�h�ǅq���wgp�	m�	|�@�~�-`��)N��5���zw�"J�- X��oo6�V��d".�,�Q�w 0������O�����t�l�d���D<��ԋi����lۢLB�s�`�������*P���fU��H� �ZbD����Iu�p��A�{�u��5څ`R�/8W.aW��:���$��[��K����L��{�\:�
���5�]:ە0�62��y�x�@BW$ۓ&�BZ+�PKj@@w��& {�h��	fj��-Ô��itq��y|1�nxHW[0P iR����3X�Kme������e/�b�?�f^d�J�荗�\�>eX�Y�!�� �P�_h�V��9���L��C�$�ϯ��抾j�H<�,]���CD��&J�׶�F��2��,әڃ���Y��V�ֶ݄�;Y+�
+6��#qE�F�z���O�B6�q1��݃�F���x4LE�ǋ㸥*� X�5��Z5��]�8��p �3'fyF��c��AQ�5�����&f�v�`��k 9�,$>ػ�Qh�%	�c ,P�[�[��
��`�f6�݈�à���6Xʏ�O,���Ag�3���&O��u(Yn?A#��31��̢�E~���&#:l�a~���=��[�v�d=���A��P Ϸ���Ψ岠�&?f[q�߅N�����}fn�Q�BOײ,���Y��t<��L^�q���'9�s�_L�@H����I�������~�z�[n�L�t������Ek��zҴ���a%0��_]�t[��m�}[ {�����\�Q�ch̄�
�~1{�B�S��6���tNؕ��z+6�>�SF^z� ��?U�r�\~{�;�����u�͜�w<�wr�����bj����ky�c��*��hŠ��2��@PQw�O|�_�{H�]`-gDGk�Q5�- c(�>G6X���&Ç���d´�'�� �H�XM��}�L!��d  ����*)�=��,�T`���@S�hn�udmY��i�s�Oe����(v�O�c�~r0Mj�α$�`��$>��ga�%/;�]T��\?���;��"��Dd��2�B���:�90�nn�I�T�1�h�n����
��k*</}gd�Oj��@2�+�u��r��4�E}_SN7�QX���� 4ʌ�"��ї�`dV�7Ѽ}+u6j���j��9�3Uf[? �6�4 �O!e�(������_�A�I� �\p�ю�Q�Ji�[�l��:�-l6 �3�s��gT�yM ��]�OTu=��]0 ����&aNRP�������~ �?���嬑L��Z�4]l�{������W �&ehWCH�I�b<%5��F&P��f�8��@�i�N���j���g�k��O� 5�]pIP�޼ �vd���БB�Z)P��@h�B�pt�wl��i�L�9���b�Gj��16��kٶ|`��	��W�B�����k̡�lے�4����cπ�_�0Lx4�7�ܖ�7s������_՞x���3�xQ�4�^.%ZA]�x߾ eZXi�H)�9:	�o��Eʠ��^%�AfwcĄަL�*���y���/�����0RD+4�u݉20�S�^�,�4�!�IKw���1�>T�A"��1_�x7��jW�q�����3�)�)Q���/�#�X�:��ZY�Vx�8��L@�P[���7S����]�M�W��.����^�5��[���=g���+ԡD�Bh��y��ɲ��~,W���a �KN!�c�ξH�
(�\0Cݽ��aƱJk-���9����@K1 � w|zM�u���=t}$��bbA�XM�P��[@Ԉ��U��ז	�X�;���$�Cձ�����AҔ�&
K�\��U�K������2�ܾ��+Pm��3W���V��e�q�N.߷�2�<m&4ſ��-�	��5�b�wz��K��|膬&��E4ko�zzf�Juܛ��4�@O�ɧ�ۯ��M��|	��ڴS�6����=��)�OǼ^A	�	���\V6�����!�HKE� ?��8��:y���{�|�X���ӷ�x�8���@��\���X<���4nH�S�)z&�M�
�f��ʹ��-��{�)I8�R�j�Y����ޱ�j�a��ф��W�'K��i]�Oe��A�l]�M�ɓ��,�B Fq��M{��.E��2)�Q �N5HD�˯C"Zv �:��?���jl�OxKB�ս�n�ʛ����c�Ԅ�'��r;Zo2�E�h5���ؿ��_���` ^�Ԯa�)L������U���� ,����#\�-�o[sS� �n|)���u��0\6��G\�d�����<j���~o�0��2�u�bč��^p�B�	踁���(��N�f�ʺF)�r�X��88�&J~�&�΄��0%�x��|Ig�%�NA��kQ\��P4e���K����P�ˢ >]�V$���
fdp6m�6�<(�0%0zW�����HQ�"pq��p��CbA0��ځ]�������%�H,"Kf�5?І�n�⢋�phvd��e֝}n0�uW���pm��/�:�d@����x���l!e��Lqg�piF�#|��t:��^Mې�bU���G�}�>H�
� l�Δ[�����`�r����bL����/�K����:i���w͂@"��z�5҈TNN�5��ܙ��L�i���=�c���w��N}��|j��^�`�e�}%�UL�ι���W}���Z���1ތ��`�2����:�>P����������@�d��ޞ����)B#��ƌ��o�Ip�Y�#BG �)���b����_��|;g�5��]�m���j�*�����F�T���\��G�@�bƿ����Q���Pj߆#�/aO�������|�3�Ή �]�@JphRc�9�+ mO�_�B�r;^�!��� ���૿���S��ڽ{e��]Y�7�+>򮚽\�S;'
��H��ǝn����h1n$��?!M��t&B�h�6�F��n��P��r� ѣ*�3��Y8y&ހ3��~�׹0�Ғ�`D؄�`�L��w��A/��p�.!�u�,)�ׯ��
I�)ݬ^5�������h�)[����n�Zƣ��T^�H��mx���<(�2�}8���Y7녴��X
D	x:����	�g|6omx��M�D�o� �AYg�zyȜ
�����N�_r� `�1����0�v�����zszɵvYze,���W��4�����GA��,���^A��'��o�0�Y�U�F*�j^f|&4D�wվB/F���=Z�?k�5���vԚ/��t�@�0�-Л�1V�)y3�=�`�tt�i��ؿe�i�t�F�b��DF���%�C+i�H��u�X�xI,�.}�݆5�_�:[��y�xq �7j;�'�kH��g�D��w��͏����1
�l�����'w���4�e�5���{�_�?kNsMx~�rZ2�M��Dk"�8P &��6�-W`$��������] �Q�9�稓.��U"(�_�����u�-�uX���hm��4�f�5Έj�ڃ�>	A��#rcW�}�����k?y�[�d~j�ABm��8(2-?i'�c�DB��قŇ<�D�'R҆($
o�0膖.�
Ԃ��x��t>y�O=��a��櫈4�;@@�Z�ܵ��
���;h���`g�	z��@��I�Zr(�;t���!���)d�З3��+5��Z�8�r�.�*��Ȗ�v�81(��_�:�BV���P�~��	w�Vg��1������++p��|�mbǪ9��d�<�G��ҬZ�ά������Y��L�@C�����qE����ܵl���Xu�o����ڳ��[FS���7噮0�ߋ9��Տ�����\BX���C��E��5�Hf��jj3��;A�?Q#c�C�U�to6<�ܶ˴y`�L����ja��U>$��3��Q���0N>����t���jG
%���2mZ��<NF2�r
4�,�FB��\=<�&]�SW�<h�~��a�8��}����at��e��|���-&��D,Q6/	�J.�e�����6�!1T���XJ��aX�^�x��#A&6�fu)9�â�����'�pFYiˑ��8|��t�&��U�vB�u]�1���/=S0�t&��hf�!'�Eg1�z����hLj�U���r��-�מQ4$�l������P��?Q�P����$C�n;��%s��Z�-=֐ ��N�Gp��[:��0X��56��1"lϵo��7�'�a&�l*w�~�w;>!�"xg�k�I�=����iǺgzF����FPCɊ�]��Ho�9Zo�C&���g���R(�D��f��AJ� ��\��v�� P���(������ip�{W�`{A�t
���j���XUh؀�5á	C���uAp��h�+�&e�W0o2��N��Ձ�����!A��6�믅�N�Si�*���@���,a2���X�TԞ��OҬ�
j�ϥ��#����Vq���peS#T�4�&p�s�H����Rv�k>��1W@������`2H���vN�!��Pzq�5p�5��l1�N����2���F�jT]l&Ks��缗�T�aj�y�M4��b�:�F�Fq:�I���iZ��>|��Vc0H�7G3߱ԅy���\��$H���`D�Be�F%�$g3[O���������C��һ�P&�����<�vJ�IR�<`$&��
k��	9wF:fq�3q�!r�5�DhuT����F�W鎻Z��v2���Z�N�nd)n��yx�Tw��
:�U�ۃP�����vo5R� \Ɩ���a#�b�9�F���A�p"0}@�G��m��x���g�$%�A��l4CWZ�	dX%��B �?�~[�Ƃ�%�[�Gc
K������wS��}�)�PS��ߦr#�c~_���a�N�AB�3�yp�K������Q~���,�)����(S{�`�0���03	Fw?�Hzƻ�A�[n;UT'"8�2?�t�����Q�Tca�h��`^�ji�	�����zH�l��B��2��� ��kΨ:��!��\����!������݁GS,�zD�|��o���_~�3����rs�p��>2���	�s�X���<'����+��40����&�U"�z���	5H�x��l �|:|)�5������9p�Yg@'�� �S���d�f� >b]̚���1������<�����h�̵���͠���V���=��/{�_��F6�W�|��� �S�R�0��+�@�QٿKJ2�
��G�Z����0f���5�d-�Ȩ�+��j�!��cX�G�����S:\*��-䣰��۵>�o�<B7o��)TT�	V���Ԥ�A�5��������\z-���M�y�?+�anGr<yz.��7�F�Yޖ�خ�^75���[�Fs��?��B��TK&��RZ=�d˳yq�2yF��6��QB�j�F�	��(�P`&h1�f̴�i~x��~�_0����'M�}��ۻcv5K�:~}E��.a�/�W S���g2�g;�
AqR�����j�yɿ�@��l8��r�`& ]�49�|���o�:8�-�)z����/�D��I�i'�d�	�Z�`�L�sR$� ,r�SN��]�H�$I7���T�P�|���x
x��г��{ӣ����y7��zE�yO]6�O+^���a������ ?��z��Z"U�I��s���G̀Wd�M����|k���|h�n�o�����E�����;� ����'�f���湂䘈�L������úJ4�/���L��iu%�S᱾���f�^��9Uj{t���K��eT����~˝�z�d�����2�'M�S_������mz��1*�{uT��FM����dF���7,d�f��*�4�S�r��>`E狀�3��PH�2�T�}���M������/���c�1ʊ�CrOB1��+/Ih#l�[8p��Ce+d9J�UP$�ND<���{�%$�<��[�m^��G`���j6҈����=�}�p���ET�T	���~�c��g�K��L�S^ƥ���~06�k�L)X%H��g�6�m]���Jc`��end����!U�ݢ�F
�ŉ�&���q���4�¶'��H�������i֐�a��A���F� V�&�gB��N�`�?f�`}�q���9�/]	y�e�d�]a�1M�Σ�m�wY��JY��x��`�+!��m��B�7_��DTvM7@���P� 0n��L��+��N��7�����>�Ns�KId(��Ց	�A�.�	��\�\�o7��{���|��� >�M���ȉe�ܗ�܎r�����ax���hE�+Cd���
�BI�� �mA�uY��fK}R�)���H�
C�+��]S�5mr?�(�Z���:�љ�� �E��{[�����j���$���Ņ;Jm��i���g��`*gՈ�;�Q��M��ڻ!��j�����$nG2&�L�R倛C:Q�0%� �j�~vl��ڐ�����[�G�LN88D��^$��`�.L˅E���H��oa��]T�y0i����r�8b<�
��v���A�I����V��$�ĩ�J���{�ң�$�K��� f���2�-��1X�/ˢ{�,�K��;_�q`Zۣ��v0�p��%�E�~���E:�7��Ʈ���FTy�`�Q[F��y.��#ƪ)?�U3�g� �g�����MOca��t6����_p@Mz�$�p�����yd�J���R�����KO�P �$e�W�~�̮�Yc*7T�*�p�����M���W�^�4�uV�}h�/�L�>y�-+.�T��[��o�y���r�x��C��39�@��u����+���6���=��~�����d>l�K���?}�`�2�٦���Θ�,z@w���VBV���0׋うn����p��*��J��4������A �S]�~�9��ov;�����}��gw�&�̝������H?0*��ߐ�+�Tz%�v�dU�m��U
� ꈘll�����+��Y3�mQ���[⁚`��8�q���|{c�X�_:Z��J�H�w����N��LE؏jMA���m�v��)�(��|�J~��"��,~}~��|�H�>���P#[	Gs�F��G��:�W�Bk^z��Z��<K�lI�i�
�KO��-RA�0M\R��i\?6`���#�PX�ww��t�9V/:E7R���x�}���{�����@�GjՓ�ۀ�Ż�QG�Kfe=��.��BȊG4S�,&��U��Po�0�C^vbۀ��uT����tL�e"��	3�1Y ����5�e���@R%���!`���0��=`^6aH�wE-��T�{ud���h�z�5l3_�Z$6�������)I"�l �y���@tt^��� .��0Qr �6t��l��h��vy��y�� ���Ҵ4��b� |�z�I@c��|�sn�Xș���3ȭ	���7Լ$�bx�;;6�/�E3�\��84p����\K$\��yS۷_"���皧���S'�*��b�zd�$�lGn�שB?"�����QDU���U��i�SAu㳓|RtS�`w�$�e�\V�XU�D�5E���H� ��t�)]`ߊ����-� ��c�K�)�<���{@�vh�$7l.�@��z��DF�k�k٤���g��j%t��r�!#Z���J�6���X������{w���@d�?�m9#�����ο�N��X"6܂増�����y�5-���C��k8k��Z#�	 �#ᔚU���Tπ���W\,C�9��ko�Sl�S�W M�	���(��I��B�!�J0>�Ե}�Pņ.���xV�+Rx�l��a���6?��9���IRr��r���D2b��}� B��f,���s,�����H��Q����8W��)�a��`�j��:o)��SR�;BT�f]��v�;�a`�!E	���e�M��F#��1g���kH�؃��9}�g�TM�Q���=�X��i*���qϏC]��2�t[\�$}��IίFY�WY=0�SuHe�!B,a%Ӥ���4��Y�AXF��,����D{��̦��ռ�g�d.b;�^ K����ƥn ꧃f'�8�Vt�9`Q��d�Akx������o�����*Zks��Ʋ9��85 0W)ݩ��F��aݺ�v���9��Zu��W��}�sE�^������U��Cj_�^g��Ta�4�+&K�$���r��+�
\����}���J�̗�s�lK��4�.9�$~����d��`4�pux+�
�qv��;�-�+���i?i�ْ��[�u\��*���M9[2���?�.��?7���Lx: ����kA���f��R���_5���jj��!z�a�ǌ��$6��P���r���C�5�W|�_^�#SC[P��(_e���Vd�)�g D�F�Y�gHՊ'��$��n3�Cx�87�*m���f�69Emnv7� �߉;��~�nv����Bhfɵb��)�]���p����ߤ/@�L�=N�S�O�6t���q$L2�-�L��;��^�;�:�{{�H'J\�
'���"��a�ƫ����'a��&gP.O�(U����P��񱶶/u?���=���[���UhS������mHa�7�D��O��]��!��yl6(�n��(���w&���ug��o�\�f.��|����A�P�T�wc[�X;T�v�����!X����sK��߱��kR�ڑ��#̩�y>
�j�m�7'�˖����
�^�O�w��`F�d��k�N�u�{��ذ��x�cԿ mA�WN�uJr�f� �r���{Ʀ�ҀE�L���;�ӿ�E�ӰOa��h~��R��"�Ld����b1å#:b)l��_��Re����	�\�/�x����6��뮚f��D�?6�c���t�VZ���4<6;�� �^�Z��g�A�m�%��Bí��Br� u��4�3����{�]�bN*��
��i(��\|�Hv�� F8���U��;>!#�0Z㪌jT���]�z������xD`S"UW)��BlY�c9�C���~��|]���}�L�d�Ϟ�J�R:�X3�Z'GO�.�ʜT�0/�8���-As�L��@P0L��N�?G�Ii�+����x<p���#�."s�_��,x��_`��_\�75;"��i-W�y��f�{�W�w��A���Rj�l�N�{���������B�@�6������'w���+t�t����<��BGy��,�r5�z"q%���R�qr4�@��Ӛ�����s�C$�N`OF�&E�~L��@��
ƍ�A}:W�2�0���z¨s{z�-x,Rl~��B=2���7z$
�f��p��^M�	��sϜ����r���ܪ�Xy\< ���0b�G_h�,�Q���U�]�a�
X?Xb�w�qK�R��2���b0M�|H���0s?1!>��l]R'�ɂ�|�9M���i�K?o����t,�ņFҽZ�XkϫN��v�d&wT��,Ը4�jFi%S�|��s����j���?�I�pŐ��g��`+ mPq������VWxT%y����F:��ŉ82r�����߻��Q@���gk #_�|�ב�>h�8�FjB�R{|E��c�-�M�A�ί�g=�6��6nu::�����%K<�{^�ɮ���$�K<?!�&�(A)��"�b��P����}�?�i(96����6]:�g�t���Qt��RK:;��IF���˧�k�Z
"{m�)B&����=�_��i��wYY��`�X��2a�{�aɑ6�����:@}�y�	�dy�^� ���4"zmЙ��8V�b�1�͔��B0y
@�M�����I['2{����Gq2���&�KS��-��Dvq�=|�8m�*��D֦!��D�ԋ��	J����+#WpF����<�ч��+X��*T�Ͽ��Hf���Ks����l�Mmt/,�0���~2�/0\\RZ�)��c�A\�'�=%	����F��gF�Hw���!���M4���v���v�b���_����T!�A"+ �D�u�0��\m��y?���'�S@BZ��֖W:I�ޤXR��ٮh4A�4�v���?_\���+dji��Γ�*�����e�⇒&e�Q믎�i��&��փV�2��1p���}�GiV��S\rz�)k�tk�낭��W��gc��"��d@�����6<�������f��9�_�k٧����L�Jl�#��԰ag�_�$E���ʊ\��dZ ��q���~6����	\ͳb�t���<7g�<Q�3�3�������W�'I*��ݸ�_B��|a�,�S歽e�՝�)8�2��{�!����,σ5�<�IQ~U� �n�\�-/H�|�5��"�F�M�n� _��/-g%��	�a�&�"�(�6�\K*k������t<�-h'F�K�ᣥ0B�˦�E�0��e�� ��P��4}2���Y)mB�t����-~ߗC�Z�P3�x�t ���ۥ	�n�!�
�X����JLQ���{7�WPt�rd]ȩ��
������x�{0Q�f��6���R���t�y3����ֹ�3����%�j?�������Je�j��������[�B�B��ت32ͫb�����ɸTT��x��y�"-��
��n^�6}��aV�^_-�^̼r�7��H P�f��뺙�P�@1�������O��fY�t���m�A���={��>�f(�-+��E|ޚu��'�o��;&\L�܇�����0]��+<>��yP�����}���fz �i\�y�.������C���[�:�c�Im
��O�ť_�m�$1�_!:xM��䗙f1T����uUh3����qGAD�����H8/������b�W�:8��H����g��XNN��k�-H��%Fe������#�OV�E�2�z�P��O�M;�Mu�/���th���E�A[K!�C�θ�)�����Ì��5�,���	�R=�^n��nh�ٌ�ϼ�����y��39,�l��%}�x�� �+78�Tٽ�q]僿�o�k&\�Y)��XW1.�	�0���Us6K�2Ҷ�71�,��;�RH�/�$yVr�)2j�>�n�!#C}�d��%d�{3"���o�F�	1�6P��=~9kU��?�)#�Jj�fo9��n�`���S�̀�lv�-`�=����(ևi@��\���_ʣ�<���倳D@4%s�!I;U�C¿%��
�����S	}ݺ��(#i)�ITb�h���=�x���ق�m��4�~��E�9�,Y�z0W�}+}�)H+]%=� ͯ���{px�m�L/\���p��H��(V�n�Es�϶��+�@��8 ��⺮��A	�R׌c;�'�tBT�洟��)�	]�x*��6�e�7p��H�s$�SN�6;n+?M�$SrAoШB	���[r��]���_���+�	������>�E�����������<�ބ*P1]������ V+�|a`mq���#��J�t��o��s��6�݉�q�?�W�g�勍�E�V6G�2�	��G,T2��7����2zqai(�n�yP֋���B~r*�Òץ�0Í!�?G�LC�{�'\?��c����z0`�Jq�2-����mm���5Gv���¹�s�0�9�zQ���yVy^RS���@�<1P�]�ll��3{�A�'�r����{�|՘X@�7tz��͒�oDt��t�����itX���������2}T�d�b���<��tK5>k�䧛^nF�����K��\�d�c7?Q}aq�4�_����rC����4�H�/b �ѕ��Po��;@Z{�+��1��>���롁Zj�ڔ����O��XA&��Su���E���F����:2iAߔ��e�k�}�UO��@®��ҳR��n�M����g�菰�����x��M�k��4s�Hì�c���j���R�)�i�|��2Z:�Ob^�:���n�'���L�����[��x��4����W��b48x�޼�w;�u8\��E:�6�̃�!���{6�w�����&G�f��� ���hmT�I�:t6�4���dN���"i�pe(���3���ׯ)C��@���/��=�2�.� �:��]`�y�E$���������X�cC�u��Q���s���-z#<�e�t�(i�6�輒�)C��,X|�Ip/C��Y��}�$c��Y�g��-A��B]C� x�l|��3UL�6\��%|ogq��g�K�E�_���24l�¤�_Lx���iƦzʾ������NG�i.M
��߁�&��B�ы!}JŐ�C���f��#J����
�m"Ԝ`L�j+F�ID��p�Z/�P�"�#�nUԚd��I�
ƥ	K�m�9K�$��K��aq9ͅ������'�ܐ�6a`�Bj{�sV�ѫ���3�d�2��@�6�wL�Q��%8_ůs�Z��5ʟ�*ɻs����n�}>>���y'�_6�vi�	�&\VE,�$%�M�G�y��e����h�~qաk,UxAhى^B�L��:���g�S��h�������8�k ��S$���+��J���Ҍ[��������y�G���T�M�v�(1+�A�<�&$����m"(��pe�"�/F�YW*�Ƀa
��ܩ�� �lX�`㻾��AgR.dUZ���<&KŲ;�I�"`�D�D�r�׾Ÿ��"@K��%�������e��Z|2g����YX���z4x"�_rdQP�]�eX���͝����-ㆶ�#m;I��U��|�KH�B��_���
Ut6\�X����~�Q��T�Y_��ܹ	�N�u��J�>�����E�^i�@�R1�1\�]UT1�]�} O�%�N�^��49�H�Fq4�$���@�L?Ŵ�����S�������5hm�m�.vK� ����W/Fr|���P�K��M0�t��+����ҕ����j�ڔ/�
��~2��`�ggUI-b�t�}{ ���ތ2�A��ªg�m�oi,�.��,���Ѽ������L)���t���Hj�M��f�ӒR� qH�r�H�l���wf�")M�k�@O�U@Ϙ)�7c"�+?���Fh�ǐ��IoH(��BVD_���jp���%�lmiV5�-��T����Ii�!X��`�8�N�N�<ZbԎ({�� �Yi�.\A��g�+Z�����^�[�_u���bt�^W��ҍ=��ل�:b�p��c���/Ph�	�[L�ft�y�ӬK�k�@a{̟IF���� M?�G���T��Q2�pPߠ��*�<�ip�+���]Zo"Y�j���C�k�VP5��ధx�NA �t���4ȥF}	!e|/V���qںI�0Q[����S'ݵe�9�Ot�p4�b�2}Y�]��V��G�G(�2ʦ�3Vr�f�&R�j�i��;�]Q�gE�x_��h$������{�8S�U�W�Q���D_��T8�����<���O%'�����	o�p��s��y�
���okoTyZ6�������ԆKrH&0�Jl=c �2��:>ER��
k�(SMBq\i�����#�7�<���a9؊���C�e!5����[�׫��~ 4̘*�S-�lʐ��6�.��T�X���+R�~�k�`�9��y��u���M����n�s�Ll� hW�v¤��kX{��i���� l�{�/���[]�h��e�c;�R���v����=��ͧ�	���COgVs��(�!v��Rр�eưݎ�^瘿�e��l��/U����u_���d�?��@<�,�s9�tF����Yj>4�*�� �eB"�ڔ�~Ӛ<�/��������%�Ģ�!@�q�Qf�2�8�5M�7���k��ă�jۚ���xk��W<�g�]s:�����So5�2�ػ�<�k���z2"V"I�@��rj�V+Dtv�ܙ�!$�1A���4eS'y�z�Y9�*��:���o�).�w\�'#�Τ	 Zir�=e��44��W��g��d��wo,��Y�3�UgGp4e{�Lv Sg?�?'-���a-Ly��cO�S*�0��b|X����!��i�gW$?]�0�-�>$�DeM 2s���|�%/�C3�$����xzRgR0ׯi�"�PN*1���e����� ���T!�8є�
���Q�x�	:Wp""�ɝ���&s���a�<�5�ks���xR��!�d_�9��V��5+8JE�f�&��[���6u�~�v*A�͔	 ��8O�;U�7�'�<�w���/�;~tD�.~;2��i�7�l���-�x|��4R"���ҔK$�Oc=U	�q��?zd��9�4q�!��5J	��Ɍ�i*3!�O�P1�@�պ�d!��a��G�(�l��X��^>F$��eԮ	+��O�(g�[nt~�Ic����".�E�߁��YZSRk3@�<�Q~��;L��t_���K�hK��N��XH|��d��eO��/Q�����_�30Aj��7j������A{ Ȭ+Qj�\����C���keo3C�Y�E�A���*��]��
[:������� h����3��WM(�kVm^��؀f���#U�A�t�w ���=�#��YB��D��`Du����[Z���d=�iO\K��jX�)_���]��@}8B�j;OS]�`}S��`x�M����[�`�t*���Z�UUN�ҏ�����?�'bJ�*k�,kΫ�U�/��މ��ް�%��)�3�jJW�� ܕ�6/��c#Oi�8vg�J��F������ǜ���e.��t�V�)��f�|7��3�B}Lo�A���8z���x��$�39b:܉����$�Ewq��v)s�Ŝ �}v�W�O��)�?�����B�U�T�?�?Y�A�"i� 4�����i�3�X��o��rӰ�����@�W}Vp��̅�]J�Iب<�zpE9�p��~H"��.��������WɈ�X7>)���U��<��
7�żꪾJ�!<v/)��*�}��=��%exu�9�.�OߎB�M�X�'��d�_�[�ԈB|�W.{�Z�_
�%��<��@�����S��Q5�f �Ζs�H�C��$�h~�Ea�'iԗͼ����~�.D#�����,&�V��7�+q��ה�۽7tØyx4&~���*8���+?�1�� H�Z/�e�̡J"�%DA � e�#,5c�1�K�hy��S�\�",_��)ڥ�IL���9�jŐ��l����ʒcV���1t���Y;<�	�$�9Z�%����2y���.4z�h�5��0�ɥ¨[5�B�i�k�K��?`.�!��a��H�o��!�
�=�W��9l�9�/���!&FR-X���-ef�k����Q�s���}�dK��Ĺ<59�xѪ;�d'p(L^��0ȴ��*lFR����jB�H�"���.&Q±YV�S�4�/��Óؚ��f�L��%0��GtE��@|$n���[}{��šO��TSc�Z�7���K$�;�9.#�o��0Y��1���]��8ucF�
�(��z>L�b������LSw��`�#^����ā�7�I�����U�m*^�j�����n��l�	�5�[Fn�}�]�&z�a�����s.ǿ��m�Ŏ��$�^�����~����D�|��"�i凝��,XS�v�wߗD2Z�ҫ2�%�eΰ$�Nu��K�B�k�;�q\�D��2'�nS/������j|1.�54�0��Bz��ئ���?���L39ޕ>)����[����]�@j�or�I�V�g����q�X
��K����v��=�%5~�&S�D4Ҹ���O���w�����ڙ,�q>!�0լ��2I�D|jS��#eV��k1F�DxF�����8����,9� W�n�58�l�g�m��k�u<��y���8[�e��hٵ���;��i�L���l$䬑i�ki9�-ύ�x���9߯N�hl)�(�Kp�������l�5,���Ѿ���E�g�*��`�R9�����X���������N�	_��f�G_ϑ�5�(��7���E��*�5���6��p嚞Bq������K~ep��"�Ϸ;��}�x�;��8��5>��=�
8Y=ɫB#´f��V��@r�!� J��,�f�3=_'7�VU�Y�������Ւ�)��z�E+"�٪mJ^�J�Dª���i�nK�{������ˤ}���g�dl���<���5RYLR��Nа��h~}��3�bF�"{�t�nߛE�i��r'��NFQ��T>d17^.�D5Qk2��I��)s�\$�͈�W��Q�V(��7h�Q�Zf$3ChB%sۛD*��g����ypyv�F��+���ua�Q6KJG4Il��;��F=�:����o� ��	�PZLMt]]�y�eR�X�~��j«���F �r��g��h,;���B̚�wn>���ؠ(zDS[�3��T�r��3�O^�u��G���@�х�NC��Q�m�y�Ъ�kh�T#��7p�%��F�S�Ż�K�e&�X
{	���},�e��Z!�=�
gVQ.O���Lg�t�)�~%��ղ�ݡ��=�v�]�ژ��[����:~2��s���g���77���(X��j��Y�?U�U���<�l�A�E��-�6��;�:�]�a�㪑?�U8�k�g�� s���7B���)���J����)X�'�jK>��tp�E5e��৉��o~�5�Ju�&�f&�:��;���W������F����A�a���겻E/��$����=�J��L �۞�f��A����LoWX׌����xx�\}���o��f
�Ӭl*s0%q��N���v�v�V���v���r4�Ǟ�V�^�N/��F9�P��{�� �>A�E�D�K����+v����H�˞��C�F�ڴ���c��{��W�N�R0ڠu�$7a�?�0����C ��_�l!ѫ�ձZ�uo�Z��M1}Q�P+��R�<������"�����Zk����45c���*z�ÿ�u�U3<Q�>@ �f"I�c{�pt�6�y�#�0�Fx��$�5�y#��&�>�m�����0�^��g��-7iuPa.�/�1���FMy��sB5����	W���ˬ�/�ڵ��^����2���q�FKD/ٖ׏n�{��-�Sj�6&W��Ӆ�N���q�Mh~*We7���,o|1��c��Yu�`����tG�VR���������&�Y<h�%�_�"o{�Ӌ불2⩴��k�ƃ����u�Q/y��Q���g [M������=G�{���m֍%����h�T��[.��:�e �p۬��ML���� �=�9z�K\�q�X�Wz.&����t`zvl ��|��n2DG���V7оs��!b��
���ӪM��H���D�)�)��X�>]����m~�J��ld�����6#�taɏ[�`�_꜅�����ϒ��-]2�ꏽƹ"e�P`8��x�~0wX;�з�˅�>%\��*ꛡMKa�f�K5�BR>�3��^�+�e��	��t����ƏhЛ���10A�����ZZV*"��W��p�.s&gG���b+� ���R���N)YD����=,�!$�(���� ��z��{Q�y�$")�����!���c�#c��F �3tr�)��i���o�Q���+o�`�]��'d����Ȑ)��F� ���_}%�7��2��p�-OC )L��)�r	��!R���&��K��'I8\�8 P�8��߷S�&��� �Ĕ��nd��LFe֢;���L��a3n�7S������(m0��?d����v�w�(c���~i.q�����"��X�������4|T?���w�<����������#	��Ic�N�3yl�,��jrOF:��H[�)=u�y��ΰ��m���BQR3S�5f��'��I��
� WwmeOn�<��=6��76�_r	! ��z��1�V{7[���y ��C4�-��x��-ͩ��5B�PAM��B���	&��B�
w���Ƚ��+��y0�����m՝'_T�K��=>x.�w�������������G͎{�,���?k3��>.e
h�|?����
��A}�jI\����U/?3ver�_�?��#8���!G������da�J��x(������?ǲT���r�;�^�߅.g�����[^��S�ǌ�K��Ca�&b���f:�y�����<�&܄���d�B��z_���U���m�,�r�������4Xp��N�7`@G�V2b����	;�e*j�
�F����@��/�<��#��On�p��O��I R��+�Q
���,@ �˚�_/	.W��?���	�-�侪��_C;-�(@��=D�\+OAn�����q�W��%+�#�{w��d�Z5�Ջ�k�q1�쪣�
x9tM�]�[����C/�c"_�rD�����$C��q�f��NTx���2׏XT9~Q)��k��+��V�"Y�1�|��&�����1�N�Ost{m�|�P����Ty�8E�!32�@��|n���������%i�/#D/І�P��Bk�3��l(��=Ģ� �W��u���ƶ�o��$�'}}>b�8�F�PP�Ac�<X�j�������PiWS�sA���}䙯��zo8y�����XG��㷉+LP�H��yr� <�LǙI	J���{�kfo���I������w��,��H�ޣGk]��1g�uM� ��4���^�?f
��GY�2k_�����E'�{e�=����+�7�x FJ��s��cK��;��+F竹��},,d���� �#6a�ߎ���&�}���O���ˌ��6�w����A�B��S�f���2/���D?Q�� ��ݲ�����i�����%�����c<S�C֕�	:�팎Vl��yyڄvA��U;
�؂!ن������3r��3a�c����>>����
7`Yx�TA��\q�h��fk{�^Er lyޠ���gɿ��$ץ�9PI��k�79J|����}������&�!��{QnS+:q�}Ph[L�[S�b2����j�<O17�OQd����N�E�O���Jf���w�x�m]A_NS7dՍ]��>ݳ�f�iz��9�F��W����g<׸��/㧂��(�^����4����o�dg:1HD�i��������N���S�"}M���%FH���0�Xp��<�/�L��M�O�����,�[�_V�@Ry���/<�I����ډH320�j��73Q��i���lIᩒz��iUX� 
�կ��%}�u�&���'�'7|u`��B��t�`YO.,C���<��A1p��f�$��,�u\E6�d��ͭO��ʔ���׾l�KM�9S?�0��O���-:F^A��n�k�u��i���	w�5�u��ƪys��C.��I�a�?�Y9(;ЧU�Q�}�\���џ�`�f��@��ؔ2���!�*�J}��P"m0��\�$ߡ�Yu^�&ܾ�T']�$�JgF|y��H2��-׷V�/�ߐ�
%-��T�r��ўۮҟ_w"��������xT������줕}m�̪���v�Cnk�xn�?mK>:?@Yo�^��yPlTT�Y�:B/%>I���+$l2��s�O>��s+�k�u�mܔ���w�r�[�zܖ�P?�V��NE8����O�`lræX~ت�Al�!a�W�!s��3!E)Z���l�<�!J�5�e�!�Q'ޘ���Mք��ŗ����o����",�i��X 9�J+��V.�,l�p���a,iׁ��6u�<��VfX�@\��$j�����o�܂�6Y$y{���S^�j����M��e��HF�!�/���"z�֗܄���z��SyVHV ah��C���ܛ���/��\�i��C�ﾮ����ɝ?�f2<���5=O�iJ������{	Y�
Gv��t[!�����q-�+քY'z����T��J����.{%f�ƅ�]N�g�U�Q���/���ܜ����zo
���b����O���9���o�Xo��O8��R�4&�w�`���N����2Df���7�x��wB� �j(�W�09n!)��nud��IH���{Q����ETRGue^D�c Q_�gm*D��:�:�S�����l���Z4���Wy՞}�9��(�:�=|]���blw�5}9#�������՛9���Ua�%2�S�KŚ(gWS.j,k������u��Pnh�;������J���j/��{�х1.6��ڟ["�����@s=>�Q[�{ƂV?��h�e��ntkaQ�&�Ґ��g(:��vC��`ϦJ�*��+`��F����n@�w1���CKYe��Y�
���$����	;z�v0Xkh���z0�D�}PZ���,k�ō��|:�"^���ҵS�+=!z ��CA�^����K�N⤤�k8 1g����s�ԓ��^��y'�������\́�;�LQ m׭c�g�4b) ������/ K��X��UC���۩�v��Cv������Q���<A��(d|�MV�0��,� �瘂�Şj�o�ꈜ�!�����Eq���*���w6�C�h��n��G����,tL7�T/�#�D� q�(тm{|Mc�Ǫ4����9�x��u4�a��_�)��t����Hr;w�o��ێ��܁�P���(�����͓���]>�g_�tC,��ߦ�֙����y�DK7��5��B��QoG|&i�0�nQ�K9��H�6�/�geg���x/m}�m8FZe�u���� ��5�Ʌq��	�;,Y�T���c�Cf\��"yTcǗc�&|���k�X�
yh�xt4D�G}Sa��ب��Z����y��(e7�9�Q��W��%	)c�{q�"ȹ�������t�f�N�z��ik��"v��w����Gi�d1��0�O�b)�XТ5�|����f��|!�p�ʄ���D���*e�0
�����l��up��,�U�	,���������z��2\�f��SI+��l��A'�^�h<��H7��NK�Z���D��rn�?qP�Q�T@��k��9��3�k��Nę�5�YN
�e�u0�y�y� l�w�t�� `�X����?���g�N�H���@B�X�5�;���w�V�R��=��A��0@��D����.�aG��~Aߓ�*St9��%u�]�ZXQv�d��Z�Q<�܅UӃ]�s�; ������C�,��_"�M1�)׌�K����;�ﭝK4L�N=�uU`!��QL�LM��iZ��Į��0�����p�JRY�Ju�\�Gc��IY&�F�쁮�[F���?����Z�]���O&�x��d��g����*.ؐ ^��5�d����2"_�A�}>��FJ�A���
�\�+���R��g]���H�+��kg!{�~�c������!��Ǹ#��W�.��bթ&V�'�!�~"E�i���:X���N������!��_ N�y�+�%���2.�+:��.�����\��gaA#���@���k����:�( %~��-�F�w$Y����@^��H���
X`=�4@Idm��Ҿ�{v?�e?����)�%�Aî�ĤV �!��U����Zň����5�4(�=s��ia=�#���yw����4�K�먴|M~0��XO�F
�T(oZ��B��8�L{�Wʾ��ǝ���eS!4E�Y��ƺ��3��oi�0�{�������	�>��>�n#n�"h��*�섅i���n��h��ݳ���8\��-�7�߃�0ȵ+���.��� m��������;�5(xf M��:��I�ː}uU"b�a�Q�h"���L��w^y��h�.=�_6��(�,/�vt�XO�`��p�Z�.�&�=u���w��r��U=)q�5=y��f�Q��i�����O�ZN>�~b
�q��.���0�erK%H�`�.�9zj.�\`3�o�g)q��FXZP������,5�zy�������a��1�z�G�$ ���]5�N��U8��dR���jH|7�z�Q�sjJ#�ce�XX�t�r_U'�]0@z�;��9��Vt�ɾ�b���o-ms3o��$��ʤ,g��� �h�;J��Y��ZW�O��T��w�����������M��&��|�55(��#X��.��JI�.}	�7Lx2@wv��Pܦ�����\��uK%�G \�ґڜ+ސ��Z�Z	��5�+MG]�o!ڢi"4\�ҟ����5p����s>��#=�Y_]��V�t��E�c��#qNn&w��4�V�c�@m)b������0�Y���j�1�#��0C3P�D�w�⩳���n�ɽ��:.r�9��:�Z{B�f��A"}����EL:��p��~��C̤h��@4ӭ
���p-&삨q{�eL�sn�t��c���[u(���h�0�p��:�j��S�m�t!�����`G@t>�E���M�B�6wc�8�T�Շ�T��/�:�>�g��g�#(�S�.�V� _yx�(�g�`1��:��7��Nwr��p���B����Ho��,s;N��{�f���%���sMYFj=�C�"��vz|�NY�Ȥ�j?�)¹��C��O 7�Ce8"H�����|�+p���\9�-�����Exa�h����j�)#�U�y���lb���u϶���#�_��?fb���y����o�K�d!zt�\��2er�;�>Ǎa�]�$��J���[��h�# �t1p�R'۱��'��ی������p����fŤx����K�Q��>w7>�R7��ʃC�����6lThЊ��h���3�kex$+W���o`C�T�Κ��zp0K���?>���$%�xc����B��5�^#%GZ~>�qL�@���.�p�*	aU��h��_�6�����b��q
��Q��D/s)#J�2,��'Y�	H���*^`'fm��@�"�A�eVq��DXf�w߾�"��-}Fv��Åɪ�	��N�Sׅ3w���^k��O�L=���燳�Q쳥CѸ�̎�<0�{�iF$?��x�qn*U��&���� ���%-�Բu�G����nʩH"��|��p�뀌���ɈF-���OuE��Fݾ��Z�W��]ɒ�v�f'a\4M�P�|��T��_�<��z��� �' M�l4zbF������>H�a�ks�(H�����:7RI��rm*�)��d�\�� �%�)�oQ�T����d�>�Gު�<	}�'0���0��G͚�|�_^V�M�C�r�_��Rkl�Ψ�z��Uί|O�P~[��dH�MD�(C��
B�󑃦 W��kdl���n���u�gu��!'#�Y="pN1+X��}6���yo�kbtl2��D?�O��x���j5�>TF�;��>`�����_�lKzB&�)���$4�p��)t��`4�9J{���UM�4�Se6TX���AIr7��M*�
�_4+�nc
?�	��L��?��/%�$��nܜIdn��˳�{�D���g��:���YQ��Ki��n���������Ny6�$�ĉb��1$���]���i>�	��K�1U&�����\���ݛ1��ra���{����NRPj��</i�X/�����������
0�mĭt����~�"D=Q�ß������7���F���F���@}�g�$s����"���gXP��x�.�ke������jmI�J����7�f'���AR��h���V��:{�A��R����vT�(l7Iy�r�H����݅Z��P�p$�W���K� *��+I:˂�*6�	��Ɉ���<��_#�����J+y�?X�v�'�����
�����v��6�v ŗV�i�_+CӚ��dYv��O�%H�Q�woi�>�Ę�BF����Φ> �JQO��]���ئ��6�a����|���`0͒W}�1�Z���#$�#�{�/t �>J�y�O.�.G�7�p0�i;��m=�4�]��n�,��c���<�&ސ���T�c�*Q�G��l#f@qr<�l�f*-�.b�,vtriM3y6�P�&D�f���m�W�$Ō �9�p%mA	�@8s`R2�"����E#~DT���A�6:��9+�ʵ�_J�d��� )������E�X��tXV������5�d��md��뉻"�w����S�֢�jTC{��)�I7D���i���]r���Ew�=��������}BG��ǚ��tk����ϽG�o��&SOH����������p`^������X�||��*�M}�s��ʫ���
���v���^�R����cwa��&]������xl�2k��W�Pn7͵�p~��3D�Y�S���U�Z��R���r�
6F�xTyL�w'�u4�/NlS���\8ɧ����̣ű��C/˴P��_����vޠ	m��Oa��C���a1��|��PT��� S2�~Cy8�/W���GNυ0�L�-��r�@Ң��}&�����Ų�J/{�h���XW �����G1�X�l䎧`>ma�����:�ɬ;sF^U�c����Z������qjЮl<جY��%�'��L@s���f-�(���,qa�h��D<��]�r���C�[X8�u2xZ���c�S�$�G ��(���� re�re���WyxË��y����(Fऄ��'�z��y']����A	�Hx��_-Ю��8�D���#��X�j$��|��^{���W���#,ta���ۋF���T��{.�z���݇��A1�w���7
���w��z(n�"G�<;1y���� �S����i�W�_BE�H���ie�1�|-�,�|�V�!�F��d��h��j���FX����v��|�lw��MMǙk�����Q�.U�� Z�E$>�/z�*�X)��Y_e���
���Zn"Y�LFwȺ]�����x�n���I0E����q+�S*������|D�z{-]�e%�g
�V�Ֆ�a�kB�*؋���,��@�Y.ks�{�։��@���}�rD���Љ3y_�F��􃃨p�U����A.R���@����=�/�����"#7�s�p;Y;��z�����\�.xr����Ad����M���e^r�8��Xr�~pD�ac
H�z;_�8?�e�
��iz+�Zh�QV����Q�k��w|Sp��n���r��1�m*#v�sSF��ha��Ƈn(:P�شbb>�9�OdR ~��[k(Q���dX�q�o����o2-{��K�a���EJ�ɡ�OS����v�9:���ksi;6
W,�6Y����QcjG���,�0�ۮ�����n���4�W�5 �����ϊ)����kA�������-����!���O?@�Ur�(BB\,u�WzE�� ՂX�g����2<==�>���J��Vc�9e����g!�Ei� �t�|��^���=C����Ӎ�B�z�k�w�����+*\>�O\:T��%ALx�Tp�S=
�x�y7w�(ؤ�9�x�>\�8X�y�8j'|(���O�o��z�	)��Ѧ���1���I�~��0��D�g�$G� ��vU�4f�0�ܨ�����#�X���?(]&ŉ��'�m��s���L�T|?&N��{5nՈ�Arc~�z�`~�o{�>�q8C�x�� �m��a��7��D��߽�3m��O���H<f����	�·���#ƿ�®�k��a�Ǆ�{����J��P���ޟ`��9�~��Vm�bW!=�%���AK
�� �3�\�,�)\��mM	�ky:������5Ľ����gM�l3��9�ѹt�Ľ�鱾:Ks5��[�S�bA;hO�SO	�GT6ꍒ���өF��J��-3�p������Du|A��Y�'����TcF�>#3�,�6qy^s��(ˎ2�S�#,,0ğ4d(� ���]F����?�����a�8���ٯ���d1�:��WhJ�|%�y��L+�쐰�	t.��k����9��@PasDa�	V�f�-C�`���ZKH%N�c��PZ��<�|��� �/�����kÚ�R³ֶ���ue}�W��y�A�^�/�}L�V���p+&��~²��·��[�
�Z�e�g~��%	膀�����WlJ�z X���bE���bN�w`{�ޖt��e���<費\�����)��9�[��fOڢ:_��@;��Ҥcu�I��4�T��?y��Zv�-��=�.��sn�b���mtg�PVNm�6p�v]��Ͽ�)P�h
ʉa�QF\��,��c\j��<�n��8�˒x����F�s#;��RѶ�a!��0^�'�6�h��-9L׃o�*�#{+2-���k��&��`��t%�%/���)���{(�N�7ealށm����B߹w�0�Iy��V�{b8�����ʦ�}~y^{t�� ek&5�R���i%[%P��>��̫�D�`0=�KTG���u*җ��"�xE�G���H3FQR�\�^�f�U����
�`,�2G��q�}G8��hf4?,wf��?��X������>�`ٞ1�.� hWT�\kx��L�.�Pҥ�p`�#U-h����������<����T��}����[�� ;9P��VL�D�/���EI7��)�2��Z]����n�@Mf `��rMa�\P�]��@QF�m���f��P�U?��r�yYT��A���wT��gpJ ȨAWXN���ʟ�V�a Om0(۠�-��.��Y��D~�D~��Y���@��8Q��)� ��9���)UC��d��%�� �ۂ�� n�d:�2�,��<?���}�����9��A-��gK��RƜ�і}�l׏�)�z7h�8�p�P�bӚ�b��Z����BGw�y%����@j��yK�ھ_��^B���=q9.T���5Љ]G�c/@#�����V`�Rj|���|��9�S�9$�-�a���Sl����\� r�$Z���-�AM3����=�H��*�(��2��[�z�Zg��O�d�̀77
��>�	�	��?w��7y���||��yT��Q��H"������\��/�!�xh��=��C!���X6�nͩ�O�^�PG0g)�:l4\l�W��/��/������$QӐ�N�h���P��{�wF�]��l<�K���H��4�'90I5��A��0D�Bk���B��nf)������.޲��]dcF�2X��6m�h}S�.�����c����6�B���^H����ØB^c҆M2$/�銭&\�Z�t��qt;`̛��7�E=K�đ��Q�b�uE��_��J���qj��D}R@x��1r|(�=��{6�z�i@��,���J@<����}g��ݹ)V$r$n��BH�RF>?�@*��U\:�\ξ�?)3`e]�t���C�~���Ryї�ԑ؝N������®�!}�߈֐������X~���P&�,]�������BgV� �U�W2�R�����3�T�CF3�}��eդ�#�@C�C\���U��i9��c,(�5�Z�Ȩ#���P�v��|�=m����(J�<�i+'�Xڱ�9�V���>o�"H
�]�xϢ�ϲ{{�90��Q� B{�B"+���K�!A'	!�aA�Khj̷���%�*xe8z`A���B_�#㦮>��1����%��E��P�L�>��ÒӨ�������e=�õ$9��9]��6@�+��+jh1>���Lȗ� �E^�l��׈����˰B��rh1�������{G�@�S9j�gށטkH�a���lqA}>����a��Z�.ͻ�x~t�>g��%�0/W|����N=��n��QO��fU ���".��\���vv�4a�_���#"'�Λ�@�G�-�xTc[�Haĕ*�P��>�ʽ:�v�\b�1�Řx�q�����7ܠ�8K�K�&G
�xm>��:j�{��z�>��l A���w�N������ٕ���9Q���gH�)�	�~����_B?I���dk�nR����$�IA(QTVvQ�Y�S���x��N$������ғ�"�3P���Mh���uK˴FLc�ԭgmw�y�[Mq�剅2�ś\/�q��s��۵H�b�f��ۨQ�4I�1�((���>���
+�d6�a�*�AHz���㲜���=ԧ�EXT�ۂ3\���j�����ocH��'��&�w�F�%�
F�ރM�0��֍�=���g�Z:E��Ƈ ߒ\B8}]^z�JT�${8N�R*�M�]�ȃXb���G.3�Y\�t���;�q��q��%s��{2��d _�ݍP<�e ���bWnL��kh��B��?�g������k����Kmj��B$�C�H�zbv;3C�����2�$��x��$�w(���f�8[�:������eQ�7��'oe����:���)�c�E�X���b�Rc�5�EsT�� ;{�g�|�>Pv�<������\�F�	r��uh�X�YNج�~�7��~�z7
*';�7Gk�Zke��]y�R�R�e^��d��t;z�	 �_I�/+��F�G43t�&�	���f'�"����~����+�y���|���ٺ"����������tLx����ԙf!J��(�Ki�b>^�sV��^��7����%�j��k�%�V�#������(��;"VA�r0�L��e���Wւ�Ɋ9"Yt[����u�K����mO�����T�&�
-L��&��G�<����f"��d�oXFB��]�ߗ�4_D����m^�8�؅�!��}O�j�c�,��e����XA�QP�i�.����r��/�z�����&�	��tB��ĸ���_�B ���C&@!��{��ŘW��5���uH<�v��L�W�7�Ly��˵�bpK��`ݏ�u�M��ԑ���@rP'���Yg3.%s�~s/A7ӆWg��4?�LY�����f���%����-{vȀh �ߦ��7ܴ�t�r���7e��ɕ)2��x}%+���:O�l�,��x��!-s��Mħ���b͉��,�|�f��a��$���1�ˣ%�d���CQ��	���p��#D@7X{,���'XK��6~�W�ud�b���L޳�y�[NI^������8Gk��=�"5���;�7P� �� �������yϬ����W^}2j���:�q��P�r޽z%�ˇ�����Ӭ�T[9��ql��x���(�_��7"�}�5�$\v�n���/��E�80!M��+�M�P�VR�4��0�����l8X�� on��e�zY�b��Y��<63�Z�fI��d��96�X��^G=��I1��Ґ,�՞x���!���ȱ��q�0�*�����o��f���"��Y�r�C�ϙ�V9�g?[�B����/\jWC�C��wfd���fg�xbK��R�e�����W�&��*6N'#���jd�Aq�R�C[$^� N�=��]���OW.M.z�[��0V�\�I��lC^��(q���
�濮(4lO�3sUq���1����I�m�&��7����AUI��n~V�2�J�kŅBSW9S��sV�&�0�'"��5Ӫ��qѝ~����ؤ$���?��VXV\4��UWo���8[,���7P��լO&0��U�s݇b��g�2�(�4�KVo`<d$�$86��<�[��^�c�|K%�0��x�י�A����̥<b�wb v��@_�F��.��*��J4��r��V�f�>P&A�ɩ��tF�[,HU����l [�;w,�q�N���!�~���h�����zN\w�I:clw����=V�wZ
7^ �� �ㆬ�B���F�O����fS��m�#F�[K:T���ғ�����q���w^,zG�T_����<L��uh�=�3YG���s�e� w������|�v��\�뀧�q��t���������i/2���� ��Z�Vh\�f�P�UEX���]�n,���K9���j���&̔`�Dc�2#=��0*خ+�w��qӬ4e3qp��*r
�?��:Zӡ\3B�6+	�B��A�ER`������U2�i�k0d�Ի����/�?~}*������
���F�ģ��k,�l'>�-S��S�NP��i{��R6��`z����F�rᵭ���:9e�[c��	�Y$Qد��6砡s�j�{�r�x�:Zg�LE�e�c��/$���Yx%@�'.�2�{+�|��e���P2Ә�Fr{q)�o�u��!�q�kS�'��n?�=c���W�N���E�O��*RD�$R�,�2{��ʗ��Z�`�!C�V~�U�
}('�坥�:
�I��Z��;��ސ��I�o�Ow�c�52Z�o�m�!�Yp�ފIT,�:����M�����ݽ�B����^�A9fF�a��kO�j6҆ ��H����ǗpI�l-�m���@����]]�@��[,�AN���1�5�o��z�r7�i����{$��G�ƻ*��b��"wI��ھA���J^�S6c���PLs�ʈ�C���`�9���=؛�o�5|�f�t�9��m�'_�Yy��%���_�"�`�\̠�4q����Ԋq_�1%� ���&m��-�+�8�<O"�m*�k�Csۍ�{�-�h��}ܱV��'�$��IT*=�������T$�
�!H��Լ^ȑo�a�
��"Ţ3�1r�Qe���(�}�@�������R�l�\��V<9�8��b���ؘ�q}"_0h�_�g����1�4%���}g+�m�2�HhONpĞ8}�*u[|�!����ǝ�*��P)O��5
���uc(ʻ���Q����� dAI�����1ˋsN��O�0L&�@�y5L(Ѣ��Cf�� ��8��z���'��������]�֤���oS�l�����Q��/n�UL�p �͞ N1c"�Y͇kw�в�h��ӐL@����E����-�U��S_�
�?�kr�5�x��h��p�4N��{%
�����w��ϟ�
���L���J��x}t���jU���W�q/�{У�}������|���N������;l*Mi�4��G���ǆ�U�Ο�Uzjr�Z��N�L:�19jm���9��SV+̟ION=�u�Ju��+����_C�!t�\&��+���Δ5_d{uW�"0�|5����L����[��`�G)��)�U�0����ķq���S��r��R�|q<�dV7�NV1��}�R�(4��:Vìzo/��`��@�0�&;���μ.'���|q�X�p�cg�������+�S��ܳZG�#さ��9hk�Tމ�����<��N
t�V �׉�
xPx����4Í@�C�"N�L3�c���J1J�I��?�t�j\��E<C�s����^��m8�I��d��~�l/����&�Kt�T�Yп�(���\g�@�Eِ���V����tȍ����x���t�|����!�t��� ��9��������dF�hC��v`u$���ο��h�� �jE�������B��8�u���@.��mE@y��u�\�v��$\��Vh����} L�gl3��c��,S���]�݊Z�M���кyRH�-2( Lw�~؁^�E�{��P^T��LT������
�Y�P�J2ʐa'��#�q��,a7r�
h		�v,3d,74�.9ς����M.�[�e�O�e���: �G��<���y3��gM��g�̈&�@f�WqĪO��j�X���������G�bW�@�9�q(�0t+�L��{V��62�i�(�x}�v}� �<2�L�h	w���E����L��Y�Uy�R�>���/�Os��
[�ʆ^�b�J�;$⣟E��$�&�������|���j���5�V�.b�[=<r���j�@mܺI�b�H��������Y������6�+���?��0�,!�qQ#�őϹ�g��׹�`�J�k��<ER��Ge=�.9q�����V��BC8+%]�Ϥ�v�b�A�I%\���P{���C�U�_c�T?pC��Փ�[g��莉(�;2���O@2�x@�UR�Dh���4܇>>:�~�g۵�8����>_�X�.�(vǓ�_���+��Cg yg~2�tg���3���%Jgh3�V����i�uŬ`�#q���	��5w�O�#�Xl��=�D�fv_��S�!R�~kn`FY���Jh3.#b M�ɥ���B[��p�F��C��+�OlDk�Wi�.�&I�&E��A&��j0K�u�?A��tF�+���8�	zZN�����և�C�J�VEn d}������\��6<<�^���0���������������Sp�阢�-�G�S8v#�����r��k*]��s�p(P�(�~x��?�⃩~�We\�z��
�0��f���4TwW\x�;ӓT
. �
q�+�ɓ�����W�k��b���y���s5�XQԽ�I/S>�3A����X�C(��wWK�)��q)���j���ѹ�[�߳(�lQuM�D�B�B���Gqr�۫����B7ġx�J�I0�Av����|�?]��������n ����}�-�2���25�!{�F�`Kc�ۤ��L�b\^4&G����`$�����k�|�n����k����ZmC*`3gdH��AHn#K<�8� ��3�̹9�}�m��ț=Vt�9@!D9�L�|�!dm+|���߽��C��F8���:�-��h�};7�=���%0����n`�a:/���iP�z���z�l�J@�`��0"�����h���x��ԇ
��~���(!e����jb7�pLO����ʼ6���P�g����hb��ɳ3�@���x[Xx��k�1{�4�b�U��aU�{ ���Ѯ�����,�ET�7���M��W���L���H�71�2�k)��/&&���Z�4�i��h��Q�_z[�uOQ�D�Pc!���	��N5�=1	�_ݻ�6��Le��x\��sG��*w����Ր��J�^��?۲����/	����d�������H�̚Eu�h�W ��HS�I�J��4l��|z��JF��
(?.�Ā�8:�unZ�����Jwg_2ơ*��W+��4�����
#�'�$�D�[�����&' �e��I�}4��|i��k�0=\X,�8���ݪ_�*�W�[�h�C�9�ҝ�� �j�&��Mt%�X(�@R�ȠPtC�%�b��%æV�dW�l�`��g}��DzGp�ø�y�鰖���m�vI�oCo�"w� �:��?b ��3Ĵ��+�b	��ãB�¡�kc�^Z8���b�C�Ŕ�ǽ�=c@���X��7����?[G�J�!a�>��L�����)���#��<�ȗo���R��pI�M��J6�f%"G�/A���b��1�����C�q�R��o�f�d}p�@�����5G�֊��2+��Y�aw�<b��l�Ox "mu�_?R=��5[Ȯ%�m��%�lv��`Rm��U��j, 	���鯭������n�w�|Z|�Qɡ0�]��AN��`w[g�j�A5U�u	�yd��6dQ��A�/e��Q�0-T��A��ux"�8i���.�Ϝ�Z�v<`@3�{|�'�Ix�tR���iYK"t�QKT���z�t,qX3ϧv�RR0I�������0����A�g����_j�q#ŵ~����r�p#&�h��-'E瓊�����fjP��ݸ��  _�v��,�M�p�vV��u�,dTn&��f0���*)r�l���z��]�T楑w�����A-4��x�#�i@\�;tz�A\��$�F~��)
C���
N�;	!	�S�!2SjZ47�,"E(��H�A������D��l���=iF'���_���t]���rW�ُ���~��o��rG;�WV-�Z1��hy�Ho��5������F������נ]���!�A꜇Z�X���s�Ѝ�$4@t�J;2s?�����B�X�w��A|\XR-g8��u���a�@:Ȓ�<���Xe�����_�=}Wn��WD��S�W��h\RS
iRd~�Y�������G�Lm���+�6!�֦l�%0���R����kl����R�I�V?̠Bt��p��<u�\��I�(�Wmmr����P�u:1-�����<��[H��
[/|g6��6m�m{��w�a�㚁�� VK���q��ۙ7LʮmP�� }�P7 ����5�R9�V$k�y;~�H���X[�ѫ�ܽ�-�R��j W
��1�}����^�=gv';ԃMs�A>�Kܙ�W9E1��J�~�a
G� �
��Td�0,:��2@Bz_����L/�z?�_���W�ְ��>h���/|�O"-e�S,]c�p%���`d䩎�`��Vmk���cz.����9��6˦��"�'yI�7q�ܨK��"�϶鹛s�ǚ���IV#ls)<�� ���?�����F?(GN�?g�_�0w��Y(b���:�ޘ��5Ix�x����L������	5���|��a/<�9l�5�ǫ�S�-z�K3�]��Փ}� ��
yD�UGH�Z&��f��,eh'.,
�!��b<ϔÖ֩6�\O$��&�q(��j��Z���m�D8
R9�W��3=�/���ȺE�R|N�O��[�| ���sT�����q��g�ˤ܅�����P�����]%^�2A5��C��?���ـ&���"t	��\�Ǿ���������<V<�"��qNci	��d8m���k.��w#RZ$[4�Z���]z�:�p�yGQ@(�����^2�?����E]p��Q��(����\4�6�F٩�Z�|����F(�����bD��9��q���GR��b��C�J&����v���nL��
P��]����@�X��5&����e�� �G!��c�/��cg������na�3�R�	�.՟�c������i�`U� �o��g�Պ��2@�f�Tp��e�D� ��h��J�f�n=3�܆�]��������Enu�lk��b���PKv�Z�f<:�B�a?4������4GI�o���n!��Zg�@�Q|<a�wod�\�#Y���d1}���0�6�ȵ�%���e�nHd��Pg��{ͺ�p��;�75�u��r�!<�6V�%jOL+����Q���5�����|Ȅhe8ӼM#q�]j���0֟`��*#}�<Ǒ���i�;o��5mS.}�N��M9V���Ta�)X�]�f/��x�j���zKdMM��X�^��mz��١W=ۧ����թ=ZO��.�y�.<=���τiD��rG9��q[� �d��rt��{F.M��kcRx� o�� ���y9����Ї��9�3��%W͊��G�w�/��7�yv�˟���_oV�Ed0Z���VvK�D�Cyb�N�����{=ec�bI���u�>TU��TH�P=���]=qҗ��,�Y곃�Y����1��P�kl�������Ă�pd5�[$���Ig?V������s��K٣�ro�8.<gk)}����[�������� ���V@��=��*�Q�/Ӕs�s�����QY�
ɇP猑�ِR�^	�n��K�H�j̵*�����ÏJL#��Y�fo�'�ƥ�t�ᮈ�w>�*�+�����j�j� ��j�$
OS%9��l�ց��(���D����,���(�SB������uϊQ���z!^?K��=�K���7���6r���%k)���>!��@���x}K=� ]-K�!u�S7Oq��IX�]_�"I>;��\Cp�U�����z2P�t<�� �G��Ln�w�	�S#{L�lE��P�g�q��R/�DM�ms�Q %�(�S�ޮޖ���<F������|�(����c�dO7��02�p�.�Ocq������|X�FM˞VE�p�L�dUL�� ��aM�^��	N�֠:����J���OC���g����*p�р��9ɛ��b&��ܦ�TE�%��R��DN����q�F�g���2( �kZ��@�Yp �w{K�K�p#�H&�F�j[�N`y����*��5�D&�q�Dx�ӛ�[�@�޺����1�G�M�zh�|�*����p��ca�L#ͷ�9�֬"W�;"+��x���a���1���q�����������՛�k���p�t5F$�ݭ���L���7���"Ee��Ε,7o��}.z}Q�ǵ��i�C^Sd�D���h��j�" $�h���ս�
K��G���������K���K����\�#�&�Y��Gz�0�e����CɁ/q7?�����g���r<n�iZ��JJ�3�9]�fI�HG�*�̬:$�O��� n7M�!S�T��:�ωY���@u���k_ǩ�šr0���RZ������]���(2�=$��1�[[�t�7JGR4�<�%i���&�����T��9��q� d�(Ҽ���8��=Yyt8����� y�i<w/w3P���.����Z�"6*�O�����d~���0�&x���P.QS�Y��F�f�c4o�g��6.�y2�S9��%�k��d����%��2Fa���+�]�	?7��UMJ��s���O�t^�)c��#P�~����p��]��] r] 5�����Jf�6w�7�����Xb���R����Ǧ��h�O8��A3qW�>���-e_}�~�v��2^9�����ʗ�*�=��n�F�GI9"*�*)��p�^�
Т��! s�!,�:}�J=Q�dY74R��$��OޕW`0@ۊ���{1H�5��h=���{`lEn��Ц�Lf$�=����OF��+|��nZ��VQJqkɖg5)޺"�v��)�����t��ڈyYi�'a����ID���S�5����(_�gP=E-@�v*���kR�%���D�cK�UG�Q? M0��m �`��y�k ʧ�]��3b<�vk.�?{�X�g䩹u^ M���X�HdD�q�\�'�.�8�S� ګ~�d4 �g3��.>�~HD���5)�O�/�A�,v&����A�L��皓�J�j�@�2�\n��ΰ}a�n��h����a��wqR8y��hu ��R3[rL��Z��*��v�)����gC�/M�4/l�+&Z��>2�4���#��[�d��� O ��lۋ��W�D=�(��YE�t�y�2��D@��(�К����<��n{?��=�R����T��d�M���Ok��EvG�<�q�R>�s�W�Eg�rQ�6Թ�Ź� ��e����HtH��s=�q���÷sW+�����.�H��*�Ts�ׇڑ098���G�����:�e��E��T��M��Dv�����Y�x���Y�o���] ��<����������	�������)&��*g�!�j5�]���-Q&�eQڠB4�ɰ��uq_�-�t��G@<̫�����������k�ޣ������Zމ3DD�N���v�
�M[� ��w*�􅐾���r/��7�\���@��W�B��Ҽ�W��Y���ی��VN��r�z�W|��9�a$��G���d"xk�J2��P�Pɏ�g�9�b5>���G�b�inTW���o�^�w%�mey��2^fU�@���Q%,�����@"��ݞ�A��b2أ\�|�0���$�đC�J'�-��v�8������D��t�{"Uq9j��Y��j�.�Y2���G�?"e�e�*��>3������������Ϥ8^f,;������Zv3]�;����bf��& 	�op�mo��գ��׮[=mmjڧ�r XU����W�I������w��uG_�;�q��OJ]m�I�$I����qe���Y=����\��`n��ܜFZ�U첟7���h�~��W]�`[I�/O��LB�S�4R}
���h��I�"�pēU���;�M r�����ݾ�M#�&�ޚ>g/�Fj���۟�Q���b(\,����w����X�ږ��.��ΑUq���3I�>����I���B��oA�ؗ$��D=h���*:��u~��òs�R���c����i9���<�n��g���������xߔX��q�A��?%Y�:8��w�ᨵ*�ߋd�I� ��	����ﴯ{�j,�@�z�lQ���ޜ��`F˜�i��ZaRo\|�~۱n�^k=�~���噎`����RS>.hX#���:�vd"!)<��ڷ�m�����������>���`���uזCA'tAo� ��p�}����V7����G��a �$T�Y�� �3P:W�����8Lq�?�8`�{�0'�|�n_�"P�d�	�?��vqg��	����QS�钬O������O�M��Ѳ�]�A��ah��yV��Kg/݉�'��δS�&߾��l����<�c	����yp�`iK�$��p��%2jBty�����,��M�AL�9#���?��X��~�A�U����JElk]��A�пM��N,��F���bo�8}X�af�y#���ondM����q���m���z#B?�<�vq˞���M^��}DOM�O�W�U���Ç4}�8 �:�j&6��g&��sa��b�E%9IB�IKV7�F}�R$pB
Uܦ��Jۓ����&/��tZ�i�}E�Z�����i	�r��AE�	j	��L����f�����kn��z��3����K��T��$:� ������Y��]�@[�C���ͳJ/���"�e1�
�s�.��鏴��u�y=\�YР���fL�+�dۅw�DYi�m|��/7�? f�;�q]�u>m��Ъ��x�T�`8��ɵ��A�@���҂{����ݽ�ͩ	o\m���{F�n�����mR&�0^O�m`�s�Ey�Բ�����!Ւ��<]�8-/��mB��ݨ����ڧg� �"�5��]s��B�F�%=>���TKЇn�{߿������4V�X�'h,EH�׮!��&ڨ~���1����_d���( �`K);�����wR��^����=F�;k�4n�*�����G�7��)�������M8ᾍRhI�-��L��Z!}]�[m�C󬈡mzr����}��`Ϛ���M�K��NWm����u6�V�z-�t�j���A�o����z$��U
�Vʸ�y���sb8�M]�_���Q��V�=�!�p}1	y�1����BxS �f}�ɉjFjęqlTb�z�������|���9c̜D�:�*�^���C�+Xw��W��C�������f��w�Jʝ�s2R�Ƹ҆�n}e�}�E�<�$���񵳼
�' %�x`X"[�~�ʌS&W�}e(<���Cq����_/_���w>:�u,	�A�MQ
sq��H5�p��W=����W�>=��^��#��CF8��'^M	tX�V6E�x}��Ώ��L�u�b|~k�������qaO��-�Rx��d��P�9�-����H�O-z!cZ��t������;~��Bsj3��J�� Yx��n�d��k��+�&����C�|��36��/�� 4��4ob5Nye@5��7W���y�l��A�G$��_�=I&xD
�|-s�6���f�?����1W��6�|%v�]6�K��XL	����t���՛;�U*�M��lKtg*��/����鈾\d������x�+)U���B)SFQ\F*2@Q���3�T�sHW�A
_����eݾm��\)��a�Ҧ�(����B��y���(Mր'�oN�|}_"1�T��r �T6>�qN%C�l;�G�ݝ+��B�^���}pZ�%X���$"�4����0��| ��ʁ]�*Tg��&MF\��!Ԍ ����y�N�C%��ړ�ܵ&��o���sh �q�35#��Rd|@*�c��P�K����5M�Lo�J���u�2S]�w$z�:�h��L|+�;���*_l��5�YJ����/��_�!ގ�5��`��$5!G�+A�a/�	��I�7B�B�rup�V��@�_>G�.~�C�%bM򍯝3�P��w�:9������?��?��8U�۴f���9Z�Hzy+K�J�8��L=]^ 
дk���\�,��ͲL�pZ=��K-��Geh��@{7�mi�Nj�ݬf��5�����P������KОьo���,�s�WcҰi#Ѥqr���c�4Y�`�����{����7]�옱��)��4{h��yښ��;^Er\Au����Y�/�7	�YbQ����6�I��̵�#t@�M�JP1J�D4M*���?�wS��SX��qi���m�?�|��Jm�d�wr���P %���ǿ�Z�M�IՊL4��_��bs��YF�Nw�T%���4�(|��|ܓ1ݗ�ak�p��;b��z��ڸ塮�,����#;1ne7�:���Gn����?��+R���#Zi��J������;��M�08�����h9�T�P��G���>�q"���t����5K��t*\�ՠF<."�7-���d ���O?��%r�0��A�F�����B�&V'ڶ��BR?Qb%���%!�������9���PwVvFCa��׺��FN�#�����Wd��l�8�[����f���C�(!��Ɏ���-Q����-��P3��8�91�@��0_�Qh0���5�t"�Q���C��w]��C�wۢ�dTr�<�O햸��2W#+'��0ؔ1�m��kg�&='�����R��K�L�$�Lh�W�Hd���6���F��K����s4?OBQpb�~�Q�p��&�t��9Lڧ�G��]�g��f4rծ�C�!���/�2�C4�X�{��!�M��'�a�L�B�.��`�!J!(�2��`��\-�;�Y�A��=�O\�/<V�g@��U��<B,����O����-�os���&��2�4�N6POUWr�n9�~� �����X9U_O����m��S���\�R៖ZQ��a{�ړ����I������U��� Y�^���G5%�,�� ��D�]�é��1�����l0��V���B�F�3�z�m���=uq���cf�����4�������Kcla��=D���8�y˛�O�_������8
9pN�TJ*�26���Sz׷g�H HQ�S�zhY�b��+i#���~�+��"7(4�J�xQ�-T7QH8��5_x�'������3�)�{����FO��Ix$M�@#D�ӗ�X����I��<��՚��3Έ�:�v�e֝�js��7��"�+��t�R�U�(�w�׍zr�`r��>����u�A?���
W�#��}���r���;����7�C \<�9h2�&r���X&#�^�Vq��xG�6���w�4����#����zO$��[5Vz5��!���[c�ȸ[�p������86���Wd< ��Vp`zh���$J�����y߁�l�	U�q$-n�d��Zh8�_����#,PJ=O���?/!�k�_��]8���d����u�I��hXD9'�ev�d���)�مꁼR~�"�>�'��E���n��~ �u���Պ��R�Ac}�4��M��Z�')p�=x��Mq��)��'��։=v~�L��6�G��<(P#��U�d�������i��Ɯ�4��KE�0���>��n��bs�a�:�\_�p�q�B)�]��)p\���*��3ק֦�"Z@]F&��qs�!/�+LvP��#U�r_#��?�'�1xQ�O_�$s�9%z�XD8	R�E��!B�kN���~ր��SQ�A��?@�f<�C��Y`W���_icο�b�~�X}�DZ�H��K���.��#��U1�Pa|3�rLSB��l��*?��S��C!�`'�3uD���d�gU��dI­^�f�2��n�h[]���F�x�ґ]���M_~:���뜦���h#�ǖ>� $y4;ӓ�����
*���V��ۉЊ��>�5�NXJU�D
���U��%[��Z;�;J�l�)�������x�g5���u}�"��V�k	bE�,�6ߧ��k��Ϲ�����&�C&;�\	,:��������E����2����:�S~�<S�O����L��2$2����T��)��j=��T[O9(�����J�$����Z�p��%���ְ} K��Zf�AC��d�N9VY�>Ȇ1��X��f����F�F��̈́��!>%oX��C�I܇n��4�S�0�U<�B�L�H�V)@^j�=�����n�!5��%@L)T\U�0���$la�H�W��$�:�0����CA~0L���on��Y@�s��7��ɍ�|�Q��S$ȉڶQ7`;���`~[�7h�p�`9=�Xo��dx���H{�8Ӭ��ai�B�<:�e5����,h� �W�-f�tB� v5T&CU���,A��@;���:3$�a7.�����%fb���^4[��Z��}�L`K��в0�����x�G��H��bءZ�[���V�9����@��⣍r�Ӥ�B�; 0�KaY�1�i�{W�jЅo���=�!����Z�m�}��[-��������`��m�!��f�R,P<S;:���{W-��oE���F-n�����NBE�M3�^�T2#�o(M��/�Q��%t���NN1�ު3�� ��Hj�R��8�����~��]l�s��)E����.ftј���*m{w�:m��T��G}��p{{��2��{_W�I�|�5]�=L�a��//�����C�M����29*A���tݕ:v�v�}ڦu([QT�jJ�����n�Q�� _�c,C^Q�tz�(.ZB�S����sq�}�<p���v� }�=D�����o���y�-����_LWC���Cxd,cL�&*|�d�\Ѝ{�v�p>Ho'Nl5���Q�U4l�%]�k̳�_���i�U[���m����)]��9��&oVɏ
Q#�.���[/�����'$惄�W��tv/���
 
�3-���*D�����+N�Y�����|]T;(~ɎF��OG�[��+�5G4�%��`ˏ:��w�D^��h�O,NW0�?�[�Խ���]z,���i7�b�yn̋ܘ0Wܶ��s�\���x�H@t#��V4�~��]=7
/5��w㚭� mL�9�Př�b���жMt�&��'�)��v�����g��eU��F�87�N���Q�7/HB\���q8.���6LWn��܏/-��)8p�0�QG�l ۺ�zd�F'����R8Q�u�)cH�
�䱘+�.[�p>�{#��҂	e��H�~;�q�Ϗ�`"c6�Ku�qᷞ�j��O�^� �i���6�0����.,|�r�Uq3NAF�͹��,��w���]("�\�.o�J��-�� a 3@�d��㉂&�BF��
�ȥ��&�י��֞^\E�����&Y������ib"GO��u�JūZ���Y}�,���u���{�
��mt���ђ�)�r���XCo���m�f�|��\�p�-|B�vZ�y�z��2��A��o���b�r������1pQJ��>1�$������K��Iv�|���PH��E�MW�N�� ��dρ�i~��U���\�����,�7gr�b���s���l*5Ґ�M�$�X����_�+��?I�*m�a����B�_���C�̭���.�J	��g���XゅcK9�;Ϋ	L;��h�u��a{;�@_��Xm�%-�8]��]��F�4��U�"����2"(~�0F)��}P?W&��ܕ��,V�'w�+烫_u���r�/� 2�����(�ԏ�&�mP�NS��2J��"��U����r{cq�n��%П$��8\o��4����}4v�mV斈��W�p���ƞ����'��~-^�ї�oV��e��v["�C{���ʄ��}O�q�;��]��+K�*���ḃ`�T?�@
n�bg�_Dɞa�������8j%(*%�A�C�û�r
{�C�ixd���O��UuO*9��%�%Wm��D7J�{ �>�]�Wq��J������{�����Iy!Ы_~>���;\Mk��9�nY�I(a�"E#��1��5��f���@_��9��$}���߳/"��]�i;1���+�eb�Ո`i"L�"���	\�3���T}�l��e������N� ����7ly<�I�����l'U��Ż�eT�n��iu���d��%����F��T�M.M~h��C�����[�S(��?�V|�VNi��GjkWAL���e�$�:�&�,A��Q�.�hy���:7=P��y��^tL�pY܉��J�4��Ѣ٢8�y�{1��"f���Je!$X��m 􂸟�'���|�ex@�s4��Ŕ^�}%�}�z���).�<��*a���M;�7e���qlVh�C'9�������r�s�X�e��Q[b۵b�w��9�%�����ݡ�zߔ�<�����5UkNfG���@�����$F����;�ޯ�Q+�����t⿇!㐖N��TuD�ި���[Z�wJ٤��TT7R0=�޸��Yj�=�������w�Z��`?}���ɕ������Cz>r����u���Zvf�{���������ص���]�->�v�6�������$J����$=?���A�{&{�"�iN	yM{��l��ͺi��df>��zU�o'ڵ��4UJ�D-�Z�O�ve!y!�Ƥ��o���j�G���ۂ�mI�
j���Ӟ�����ca�"$�Ot����Si>��i�e�2N>.?��A�wSG|3��io�W:M�?��֎�՞�y�H��	��6qM��%/�E�g3؎7���%(��N5j�.%���#�%�r�=C�����?��%�K2'���H�*#rTơ�/���z4G�r�A\מ���F�Q<\�Z�p0&^�ru��lVRq;/����U�%%	��~�]s�MM7�"����X�+���� {���ʊ�R׶��(�~���jR5�F�O��X!��%,[W�8N��2J�S��>jŕ�NV[�r�J�Aq��3/F��O�G�6����:ġ���束��6B����?�����$�"��3�}�Q�_�1Cb����z�k��{�c���Ҭ�eeQ��5�Cȓ�	�٤�z<�TM���z6A��u�Y��h�v9���㳰����B�}�,P�e�0�X��=j�4. n��O�ujQ6U݁��2v�7�S^�0	�,��3�%�� !0�mBLS�~S�+�U��Δ����J|:�f����x�(ZVC�l��k��z��@��hc�ə*�5?�~s�N�P�$�OvY�׹?sr%ǔ���~�R3KL��O?�[&�p�������2* �岃t�����%�v`I0�l�7��@}YLbx��ӔH��MO6��(��;M�廞����!���l�E�������-��ѯz��K!:���=̕}��L:���(tߊm�"�=�� g�Ō�����	��I� y�{Ů�����pi��7%�/���5 �v�a!,��"���k1p� c��5z��̉�����B���>�+�=�	�}ִ�1W�A���[��=#[�sDÉټ:Ν���:��Z�W�4 ���	:��Q1�z�y'�����G�"K	U�p"���Uޗ�4,����/�b����Ac<�Y3���ھ`���~��|y�!��?Y���u`6�j�=��,�h�;f���R>��/�ust��W��M��3��]_M�5Q�i�m*���Xxc`$������05��&�N!��Wֱ��p��Hr��3��?*��(��q��K�ϑ�T���Т��n����ˋh�]�^�;�0�����ȗ�%��P�2�F�9��x�;Ϧ�F�D'�%�"�K��GM[Cf�~VTh�?M�9� *��S���*���I�{q�>'У���mu��k��h��UV��(]mB���<:�^I�ErS_�C�v����>qk�m��N���Q���aG�`��Jc׼��>n�%s�_�Zd�-u�|����'̔����
-�X�.~~��#���O�p/l��f�61ݭ����A��L_dC�SM��?g2��;��^2#��1}3�y�*witV��Q����+����I���m��ͧH�	���x4|�INz;�UG5�T#�eyxՋ������\uvp��3���w�я�XQ@�itz��zz��%��h|�9��,�`�v���%��8z�(����b��Uj{���(��aYB�����E�6.�q�
Y)�A��n��5��Qef��kQ��^j7���9�QڴL�|@���T6u�Fd3ym�+�=��)�Ur����w��%�z|��[{[�V[�gƧ�G)�:m;KcjY$3�۬�� [U�U*�%�������K����߸�5�����^2��?�"Ϳe���RX��S��-z���>���5®��`�gaJj�����v�Y�B����Xo�ꌐh�����G��3点�N�J�6��v�5a0�$c��	
�T�Q�Ԍ�t�h��rF��n�Is�+-�܊ˢ�7�0�}��1���۶Vǃ&荱�����f�<�k�5�)������O(�P�6��d��=�|u.⮑%g	#KM.X�-�b�*8�rG���]���UhB���L���
�M�o�U���������!%��������e�mn~_��"�L�����!�lp�#cp;Hh�ђ|#u~���"������É���a��?4ڄRȔx�O��,o샧m���೛4�
����p�7�|A�Ӎ��_�3��n�i���.�Ď���!d܅�����'�w��2Q�sML^B�(M�/�_H�&n{�JA�س�B|������G&��9�5��z�(a����	��VK:��j�hȒ�N�Io�%��qVދ��>	�������,�P���_;��P�:�$G�7�� �|M0���e�p�K��16۩ ���"3q�Q��RQ��Hl���|,���z�G�쁰��9���� �!�X*EԳ1z�H�5�?����鈴���-*�kB5V��8���	؅?65�,�E��wqƞ�G �����	g%(�"�*7���V���ֵ��~��;g~���.^!��z屇�s�F�82m���k�9d�N7E�-;7�[���?c�o����#X
*�� Ѕ�z��:�לcS�*,��?A��F��c�����bwk�E��H�>��@*�$W�y4���+��d�l��o8BqnJ��n@Y��AO�LE��]��,HU�AN���|=�bVj�)�R��8n�jn�9� x�q�nV{���B�?���v{y}�77��+�Y
���������{S�`)*�^ۘf��0"U�:N@�F�
^�֛P%7���a�\�0��b�+k	����'�v����&(����.�����K/Y��9�%��{_��c���Ơ�r�2A�ִ�����]�I"�(��� �T�g"��/�N@�^�2�햪D�{�k����;=�t��0M����`�?V��gh�$y�Y0}�K"�H�e�V�/`�JYS�����;��b�P��۞PA���l�%#�[,�+i��H�����\�F�b��R��|���&s5��Y�Zh��Y�\&�B���}���5���x���Q���~���s4sć�6u�x�Bx}�/�Y�S[�,(�K�qZ���2�k8T��/�o�*�n�w����	�~8������a�{І���#6o��*������*��o�t�B�2�x�Q��\v��%'�e'�X�epA5-)	��J�a�8Y������-�\������x��D�5��ƩV���9
��}J���.V�u	<�."]U���Z��T�D(ҊS"�|�sy�8P����l��QT���Dc:܆s6��`>ZU���?tB8XƓ;�?\p0���M%��h)}�V�!y����Kh�&��F1��o��O���
�̠���S���'g[�)<P��=�P���w,�$,x���+Ԋ3���A�7�q|
RP뎲�RE�f�dgM&�$(�)�f'-"5����>g��8���XW���[2�A3�L���!��7Io���~r�l���&���e�m`�Ѭ��|�9�#-���ˠh���a�_�ѡFi���&N��I�G�O�&���o�WEm]��G���l�V��G���������Oխa>�a����L���/��+�)��|t�=x�;�?(��P^ê��ȲQ��҉h�"f7��%��u�.ǟlc7Q7^� RO�z���i�'�����/,j�(l J��Y��#{���b(�l~�w��Eob;��9c�g��J|	�j$��CZ^O��C/?����m[Ke5�X����MMݦ�4�£������i6ڊ0^t����؇gҵQ�߰��v��V�������<Wf}��;��0���w]b��.�n�䔆����_���GI����@�Ld��.�ɵ"�׭f�0Ѻ�HV�j����x�k��"�I�����{<3��XzzQ���
?�Bg*h���SO��g-&�U�b$J�|�N�3'<��_�a/���𻍀�z��/�f�Z.���b��-�!+�6Q���śREX�۸M2� e�͟�ٜ~XG��i��f
�nD޼,��KЯ!�s6 !�n5���9��.���\)	��u�߳w����m�9#���.F�Ǯ���$h�I ^���m�!6E��*\�����k:x�,*_c����#�+��{�V���Iҡ��18�p���Wf}����U-�p����6�L�fJ��D|��?��ڴ7�jū����r�E.���&�3b�;vjÒ�z2�S���Q1�\�E���Wj�/�\�A�,�(�_���ŏ����q4N��q�2��>��F�Zȷ1�(yy�k0K}6|f�Ш�z��5M�9�ʃȟ��}�#��ٲ��<�NKj��!>��Y����{Ama� ءpW �Q�"q�ГyA�ګ�z�ax�H6F����������1����tNOv%�2�` �N�`���2e��T��DNAfm��x��ܥ�6�:�ݬ+޼�Q����H�����ہ�i׀v+�s���Ww�}	FEg۟퀩��!m�-����T�&��ϡ�aU!X>ґ�Y0��C�P/��*�r���B��qQoUI�z��G�I���h=����Y��D�R_��c��hd��ZQ��j�R�(�4 Tj��IBy��U�DE�i
���0�>�|N��|��O>b��ۮ�-NP(�T�.�x�yk���R��lS���B�Q�ke���F����L%�u�u2�'�� ��Fa�1�9vSA�P]�d�~��>h�(��#�Zw��}�t�G�]$ib��2`�$��vF�Ć�qx�q`��)8���-���q�k�@YG�	�5=H�`Q��;��[��%�����N��o�?�o0Í韺b�Fg���.���و�,�0O�'�a�b�_Zy�2e%e���vR�����(cp�,�%+F�!�K�3k��A��+����aCd_%$\�M���O�l.�����@�1V2;	 Vf���{���*���V��K&�S��@7�M�_��z��L�˨� |�m�謨*��������D���(E�Ӭ>ֆ<�"�F��+�r��<j�k?�S%�b�+A�Si~�_"ڼ�}���9Ȧ���0�P2�\+��|�}�\�qg#xc_�P������иk1N��`~�Kv^E�����@i��`nn6f����_|��"p;�n�VY~���m��{�`�}$�tG;٦���(�<$�8��;d3��أ����i����G��,���C�OK01��8^+��!?�"�,�G�L��=���kX�k/Ǻ���}5e�Y�B�M�տ��>E�"o�!�� �U�>�����m(&�2����qwA-vH���|��±,���H�^@%&���m��3�nk]��nW��ٶ�'�t�,Ox�� D��?o���
��a���&I�g�C��/�l��i����
���E�rѩ��x��mR�)�޸Ψ�,��Q4���tR�7���	��	|���E'��\����$I�d�ac�7�N��<����S����9J 4k�K·��(C����ǐ笾�!@۳��~Q�f�^�C�J��� �{ G@s4�NDllh�Ӯ��0ˊ?~����su}E���ؼ�������y6|�>�$���hT���\�_P�Sd�sKQ�Rޜ����㰃9��W��"�]�+$���Ճ*/Y���#`����$Cy� x�$��-3LT�:an�\�&8�$|��%���,Q���K��/��uw,��.|��#ka"p,�r}��l{��[��^y�r��&BI���'�N�$C���;��ʍ�3eo�l.� M;��%{'�s�"':2��'n�w���R$�y����u{�м=+�
b��_�����[�6K�'��(�L��ٮA>�Tj��3F����;B�CS1�����܈�R,ת�6���P7�oiY�]��ºG-"MP�%&l3�cF,3��3�I�,D$�����)��TM!�5�UgÌ��G�.�b��M�]�I��	�gr�;���={仁P�Bty���܀瑦1���9~[�G!�V�;��Td�Z�i7�K�%lW�ە�*w~3K`�F�k��G��Ju��O�0zz'iS�v�������u1_��)��Ɇ��,q��=�1m���Ő�h��B����Y*c���l;}���;r -�V��F���Χ���%u��U�')�((gA����T�ЛtCw5���+�V��Q?�?�����%®H�c���D!>���y[_��w;>^b��	B�',yk�#;_�}]1���tT�"Ց|�����^@B� D��>�0�b�?��J�7X���j�f�/�����P�g���YIw�1��Z�J�J� �h�3}	j�&�J?��u�uh(q9	�����٧ ��ɗ�!k�XxjU )n�*;B�ry��UK�3�|�p�ݞ�C1 *:�g�f!���$��~2�]��XǕ�ĝ軅:>���d	�}\[	��j�-4f��ɿՠ���V�tWv�L�s'E�y���\*���LЛC�ᅻ�o/�'+�l *��ܾ؄)���aS^��0�ޙ�9��R��P!�Qmh}�	ǗQ>9ig�~j 1	Uu�B�&��+ףƲ�=�1݌��,���R1��)+;A�ÿr�*�ǘ>&�V�Z43��<b����)۔�aI	\ќ�o!"��=|#�
?D��;�Cc�=�Ӓ��y�򱟌�o�8�(y[���N^$��/�}��Ԣ�� t����J�?�ݒ�1p��6���K俞�{P!P5�8Ƕ��䪴��W&�t���Au�:�P;6�zS�)L:�Ege���ր�4.�D%A�"$x!�_/�42#aFY�VF^0ʏ7b�h{n�C�D5:0sW���^.qs��RAaǞS���k�I�i���󦑭��@�($ ޟa@	sD8h�MQ��d���#�K�/\P���P$KiQ��|��E�彫˝b�&�� �̛���G�	�%�Q���fiv�.y�e-��{�i>�y�~����Q�%�����5� ņ�n��A� /.�B�P2J65����G�`�8)4 `�2�hP���Ld���r/3dJy��w����n��+҅'+R��	}$\�	�3����_XC?��E�3kMmM�<+�Y>��э��1C�yt����|��z��)� AQp���kN�З�����!Q���d,��:��f�m��V_��Pq��D@��D��8Q���%�����Q����1J�����)-���(He�(�Z�nX1�o�l�\�W:�Gľ3ܸd����N�GժnC!�2˝�&��N��گ��ڱ���c�X�f���h��O�h�2L���ҍ(�A��Ű9	]������)$o�3�1Y�1�İ�����\�@6N�����ilz�Gٵ�j��J�Ƅ
��48{&��������Ka����w:#�sG*vh�wB;��y��%�hU"�oZ�ߣ;���w�o�e�����j�&q�A��]_jRf�A.aev���A��4�[Q���U+m�1V��zӅ�V���v���u�&Ƒ.�\Q	�T��OŚk���c�"��^� Gc>5绌��������%�ݼm�;늶=���p��?1��w��w��	]��F�=�"���r.���M��OM�fe�<v/�̴�����)p�C��QH�]8�̚�1~���m�hi���SSVz��7�IɊ��� Uj�_�s��`��\k7�����d�_�љ~D�;+)�0���K��&ik���IJ[ h�v���(é�>���,9Y�&�|��S�B�&���x�/b�)fI�ԑ�nUߖ1i��`x�ƾ�A��v����k}�T�����.�f~�gV~7�T����Y2x���NXG2Q����&��|f��
Xl�~%���#^hVժ�#Z�y.9��~�b�B�F�c� �ϱ�6#�L���Ei����8I�#��y����R�<�J������xpk�sQN2��~��x��T���~�IJwήg�U����悓o�m��;4�Z��G��pX���^<T�L�����\�ߦ�\Vĭts�)]0�$	�� ��Ӣ����d�i�< �z�s�"]`xa�ꋐ[��dn�fDQ�&趌�~�8$ל���w��^l��R�
��wBLA�/w�kl�p�����J�V�┧�_ �'[�
!Mn��n�]9h�����Z��l����O.�e���*�V��Ś�ݹ�J`�K+��Ř4g���o6��(\tJ���-������<�?�N����a���I1��I&3���w=8�Q�^�f�:�q�?����fk��u��3R�1y�`����z�𡩺#h,k(��f.U�\Z�g���'OyDw]�t`$[�s�bw��<�s+�9�0��;J�?�c>q]�7O:0�Ju�m�ظ���]��"�먟���k�.?�#����L"��S1����Y�\�Cf�˃1լ�hu�$ՙ3��^8S
�P���֧�<��[*a����n�h���jy�L��ӝ���OW�N�A$�t�<��	�9�����A�|�&G��$9��,܎��J��Ouc"T��R�h�ܧӄ��פ1?�^D�`�?��ֳ{�.�Ӿ���^�B�XMK��_Ga�ˊd9yްbJ�Q��sy!8{�^
u�sɎ�����h짪i>x A��磩�o��<ѩ�=X�em���o8��0?G��sS��/��LG��r�3w|&�퓒j�$���0U��H�q�1����~%[�V������Q��E}��AA?S�~1�M���o��?�6�M}�f&A�Ok,dz����B�*y�&���=��m�<8d�����r��_E�E��/��k,lx�ΐ�����Y*W�R����-�f-�����@a���1��)��Y�l/ҳle��ɱ����5g���A���P��B��jq]Em;W��E�X^�=Q�0�"��i�9Bk�:����b�Uq�܁x{�o��g'��i�6[���2\z�)z�!z|�9,d����Ӵ�Y�������,?���4���j��R<�T�S�p��~�����Q9њ����'�+\F�[����fz�:or���b�@d�&�w�!Dr_(�t*��!7� p �{�iV�ϴ.1�.*'^�L%(�~A�hz��!0��1�Rb.�.x8��y-��_$'��#�ZvHX	9���EK��~>:D���w�5�}���>xUb��̈́�3�;r��u�߉�25͑�z��t܊0�[TYN��g�|����6��I�x�6� �U*-6i�h������/��'>�Zi�XQP5�6.2��£�!��� ǳ�i-{P8�)!�����yC��-�RE��r$�Ө����[�I�n�B0m߮'Y��Ӛ7��}�&|��~�R;�_�V(b�����e���W��w^Pv������z��
��o���_ۚ��"i�%+��T�3�A�\�빈��a2u��5]�J6*��Y�ۤ5�D� ޮ��s�}��p�����;�S.}%JY��]�� �.>ݍ
@޳0���/���oZ'��.>0}28z�Xs@�4佔����V>��*�JWsEx���36!� ��F�](=K
!&_��������p������\�32�b������:�I(T�[��W^������VԠ|���h��_I��n�薰ʗZ�Eb�s��Y{g������5�QPǾP>y�N6��N�0�X)�-�c؏�\���K5:�]����{��N�B���]��R�\�SR}�J�$g(dj9�5�Ƀ����k1��w��wm�"��
H�Χe�_3��+5ssg�cO��2Yq���v��̥�΋��� b�yS��z�i<޾�g��˵����k�;���V���:�ά�w�ϰ����jk͵�sg��$��
H��˴H/�1���U#�=�(�{þrmج�|� �~;�*K����Du5��xӯbR����0 �fO��^�L�<��͟�����V�� ��Y��TU/Zrt�?n���WgG�M,��E�qQ>X��-�?�zN�*X��a�岼�$�i�Q�b��|����tg8]?�wa����O��Hx֣<���[�Y��L����wu��ȵ��7V#
>c�XR�	⑅���	g]��4	�d;�{>�C�@���m\t=
p��7�)]-��ᐆ�8�
�>�KU���Q[\`a�C�rkT>���ТF����ѷ�%���<�z�<}�SFb����w��(�'�,1_~�J*p��ݹ�:[�Y�A��N�T���Dp��l��.ғ�!�"[�<������Hz�aA�Y� =x�2��6��=Q����T� �Uݭ�2�{53���DNZ��NAH8������t�IY
\9\e46���K�Q��,�2��2<�B�tlOX�=i��ϯ��[�E)���DM ֺ�?��-D�O�3-�!NM~fl��Vv|�l�ڬ[��qѪ��8��D���C�, QU^���.�E�&�1���(:��3[�N繪��%It�Ǽ��` �	���S6L�M��շ-7>�hhe}�ߐ��CG�᧨my^%%�P_�&�� ��o�qWR�ǌ�~8��w),_�75�1P�����߂��8I�L����;�s����;q��cnM[ȍ{�Bw2��wX��� @�G�#��e�%���%:]pg� 1�!�4����k��婥�#��=!\����q�&~�_/s��;��*Ą� z���>�xCy�X	m=�$eÉ8��=ԫ�N+2�2����b�nQ�=:���z��W�L#?��Z��;��P�mΚ�P� ���g�y�I��6��Dhq&y�W�D
*�7?}�5Jx��!�澊�&�dYV+�fB#�����%�S��w���.��$��q�Y���}J�w�8�RT���"W����p���X2��V���޶!G��l����f ���J��O��d���b2�T��d{lv[��4~�;ֶ1&�G4MQ^N�\�-	�:�q��w:xdu�3v�4@T&�!��]�&}I�}��d�oa��[o�����;`�Md���䜉id޻�Y�̢���j��qf�\�yn�gO���ܠ8�ʃ�]�k4-�Œ��ve6�a.G�^o�o�D�� �г���.Z��ވ!�c^�!��.�VDvb�M�����Pp����W{zi��m[�&k�P���r9�:���p.�ս1j�NYM	H�^[��O�hJ_��fJ
�O{F��d\"�Ҟ�5k����8~k�F�����1��Kģ���M�: �$�o�T��+��s+�kq�Zj_-Q:*�����q�4��+��9��_L���%���Jz�?	Ǉ���kI���m
N,n"hߎo���Uo%V�l�1����TJ���3us�EJ�|�6� �R*|�[b�t"c� �'�	��I�p~ݢ�nk��Y�R�* Z/���j�R}�9��N���QO�mkS���[	VuFܖ\��%�B6�]u˰V��|v[�O� ����Z��:�2MP����h\��%��������S�<�����$l��'�`(j9A0��.t̪�{7�NU�W�.�R��O��Jg6�yK��b=zao����_3B�S@i���:��)��<�tOZ?d�_l{��8���-�w��l:LaEo2�l�-���(�됉��_Y��#�}��@`��p+/��m�����g��A��u]�M8��ـcW���kt�[A��J��ќZe ����KA�u�����CΐF��w����&�TA.cw���\;��K�tҫ���-��
��L3o��c�t���i3e0~�
�� ߞ�z����boļ�����"J�ã��d�K9���j�����ry$ۢnΤ�D�.C Qe1ڋʭ�߄��ʄ��QGuwݛ7��%��9K�/��Qc�m`|�Q�h7y���4NC���k�AϜ�bN�Ǫ�~J�b�w�G��H<S"�z����8��Z���BA�7�U��r���L,�0=!ث��*߶v��Y��OKhwIN��J��
��>����G%� �W�`	���E�6O��z��|��z��NL.�e���m�!�0�(=�����@Fe�_��wpz�3�J��k�#X@+�/ke�n�bc`�:�j`}?���ƄbzCi���|2a^K���6�G��?����DVn��#�fw�-��	�'��?Z!�����K��"�4Ǹ2O2��[&�b@u���O������>d֡�='�L�!�h��3����sSҗ�SQY��%0��qoܵ/����I� b��^@AH@\�+u��D�z#��?ig�{��B�������$��.J*�~�Mf".\��-������u$)���-�ԑ��<2�$��F$�:ZH��@f�������;3Q�Rڈ_�J�s1ʠ҂�5g��2�r�9�Bl#o�k�d@,������sw�VH|Re�1.�^���J�p��Џ�f,��1��@��[w���]	�.�\���H!E����� ��K����`����X+D�1����P��4�r) ��"��r����k[:ГH3j�#�-���=�M���|���v�����@�mF$Pg-<�B�K����<�_�t�;�Q�=$���4���8���jzV��ɭ؅�L%�sAf���5�Zm�w���b��&p�7*h=͎ɶ�U���`N�vG�-�To ���Y�Ǉm�����%P\��n�1��5�]8�:���-���Lj��	J��z�Si�nl	i��fS�O+�nό�2m:L��̔�����"���G��PͲ������E��!zo�g�q5�eC�!����8F��N'�7���R�`-M���AM��dd6��@��4S}=�*ݹ�bA�d�6���?I88�����D�@��3P}��f�%��=�i�,a5��Ў��F:4er���T��_=��џO�ݩ7@��8핗4�,d�b.��,��&RH�/H��O����~�U�؅���N�-jf�h��]9��V��W��a�G���4���}?*�=U��1z��)u=sn��A*4�3�Dіw�Z u��Z,T\�+��-���T|7��iK��?��CZtXPn�B��Գ���Ti!I��Cs�Ň®<�8{K�;�����4��:�}�v�#`�ѣg'>Z�<�Iw��6�����|�}���G,���	�ϱ��7�R+Y��d�C�񢪏.*�U�d-/�	qq,�),�`9�}��ӟ�<n3�/���Ռ�m+�.\9��fs�mH��IZ]��]��\�V��\8�C�d\�8�n`�h˹Rv 8mU��4C��e]S,}�8N�e���pu�ǳ];{<�۴����7�����g3��S�=���ε�O��]�����s�M�{M1�|���ʄ�G�T�S_���~WmI�G��p�q�~ñEJ~,�ئ'�ғ�>��I�.!�%e��dH���L�IZd��I ķ&��B$Ԭ7�h�8f�#��X$��!g%�8�* `�����e�!�{����G�0�j� �&�Po�O/$��C�☀$Ƨ.;���ճ�>ܰ5Fqx~�E��e�s��k�x�"��4�)�/rhX��_�yE%	TDQ��k�U��0�[;�FB'�P"s�������^n�rV_8���%�ʶ��.?�9~t�:�_�;�g���5�J�Bm?r���%����0l%�y���QhHlcBxR�Ǳ�cmB����=��5�8[�=*u�G�:H�R��,vJ�ɷҡ�@��U s�֐�Y�-hD���sؾ�WjI-
q�$KV�&�}:���1��,\&O%�BF �u��ܼ0v&A?`��U?��+�"vW�DS�#Yj����pSg�%^I��l��L?��E�k������=i� {�B����!�um�B�����x
�����|Hej0���i�V�,�3�j���ϫ>��j���L�H�F%�Ҫ��e�I�|6_�(��u������/Y� u�'7�{+,��Р8&}Vygf�������ŵ�O4�k�z��A瀥G�caI�\]����J�a���rJT=0t'h����"nU[��	��Er&ٻ`}��m�G+*��qb�����x7��w!�H��I���$�}pJ#Mca^��X��������q����!��������퉓b|��]i�<������fH���c�lU�@�\V��	:U�B*b]9;�8� �*���E鏚�nq�}�� ��gR��4�a�TM�:;#R#�[��9� }��7Co'*W.l�./s�Uhw��{Sߍ]"g����z�:&�0-���ެH���)6}ʹ�C�N�K4]�W�6���X�TU�Pp�8C�s�K��|��Ť�^�i�3���W��I�V���k4�H0>!ށ؊P>�/ ��Q�o�� �u��q�_�T�db��AI ����^�QY���Ͷ<ծ�,���F��"N�a�L��.�^��Fi�~~A.���"v���~��H��W��aD���3�HtJW��NI��Yjw�_o�%Z�u|6GD��:7��q� ��8��WH��~�em��E�\j�S -�)��*/sm��\�ƨ�δ4��a j�a���?��!3��v�9�Y�^���"���Lc��/؈�Q����$V:]]�?>6�H��-�_)���߬��,��Q��͚Gϑ���n@��f�p�H�$'Y@�!\�h�];��ե&|�����G��L�SOU6߫����3VA-���V[���P���`���sZw-�����W��D�����E���1�Gyu�3��x�e'P��1(�nP
��A	ή�
�0uQi	o�К��JLB���V�2�rZ%�ɽJh#��� ��}m� XK��NXa���&ϒ�p��u��o��5�lx<�%ੳ��V�B'jl�N��b0��8��I傒�fM�C���I���ڢ�V"��(��5$?b��5/��X��`X���O4�-��s��"ŗ���2B2����#\���M�i���_�4!8�(3��ȯ��q�)�D��_���6]��������>�HS�ip�w,�كu��y}�=�k���D�Z"E��U��V��:�h��2�	��hk"Z3��q��%��)�\��RF�az+�g����u���xz||�X�F6���(��$�(�d���^�f29�皩�oq[�N�0��ֵ�핝�bS˯0�s�۴�9^ĉ#l:5���f��C<o���x,����B`S�E��Y�q�m�#� -F�ŞK�����īP�!D�9�x<5�:�b�6�)S����zYke4�G�B@�k��qi��$|��֪a��%�QȎ���똂�[������0��qB�~�2x��5���t�l��f}<��<�\ B��S�8��(���IGN���OF&���V��L���͕�3"j�1��	km�������]��W�OS���U�c���_A�d�����4�TB���{�A�����d�5���鷍͊�i��ʁ�H[�����lv�a��+�d�����f�,����f���;�=�MK��������إ*���7���h�P+$0�|m�ztIG�(��}YX��3���1+�0��?�W�&�7H0d/�����;��b���3k2gD�C�"^2��o��.�qzr��^=���Η�.�)�[hh@�,�(B@�KO���M���_�ek��i�uzgl�
�+*�����Q�|JJ1A�S��쀌�z�H=�Dd�L�^�+ 4�Ӫ��t,�p��,bU]�7�^�?���w� m��ɥ`��DN|�Y��B�V4��9Hn8���z��r5�m�	���O�gnbEXJc�C���u�紫��Iܦ�I ZLh�5��&65��>t�6��,o/�ũĀ*�e�Zs� �pY�.���;�ɝ� "�@��ZJ��" ��p�H {��J�� 
#i�S�;�~cc݂��K=M�7��cg���ԓ,��QPm���ν���H����6���2Ye�ZN�P6���Ɓz�q;]u��	5�����x�#X�7�FEq%>���Zb����HȂ6q�y�}�DdP:�1�l.���U�X������&�������+;� yə"�����S:�R\�Eh�"�s�j��^�� ��lls�N� &�x�^OV4s��y�g!��9
�=BG�%[ 到��]-8���t��L��̖��?d'���E�t&��]��ω�vb�U͍,B���Qc�N B�|_�%�܌�J�妸�4���[u��h�oI��(���Бc�6���7����v���\Ʉ]��ٸ ��_�<eLNF���1��%�/=w"';�M�?�9B�y����DA������0�y��s��'i-�,z �(�c*��5=0(ۗ;e���C���-Q��1��=Jt��&'��ߦ������+���*�ITw+�!O~����VM��ɟ+��(t���+@�@#dJ3w0��t����+����dp�8Vz��Q�3Ⱦx(ۥ��kR`u���7��ԯ>��EG�O��T��
�&Gṭ����?Y5<F,���e��+|�{l�S��.�OB�7:�(Jb#�G�������tv~��,�E��=�`p�0\���h@�V��,�{##2y� H�ҋ�Яh_`�䵃*a�T�[�:���,`C����-����3
�9~R��?Na?�[ؼ�_z1�!偧N<,T[���α��r��";��$�[�#2G��ص\4�	��	߿C}��Q���0��»lH4��B)��h�Z�j�K�qf��:n�˜���]K ����T��T|�p��iyEZO:!��9i�����mky�N��qf���t�[Dy�QU����§'K�h�oc��'uL�u�~��c�o�A��S/@T?�m��T��)<F1yH���]��j��@"`�l+�	����҇[�\ܢm=�RLR�O�k���p����~�ϫ��t>�ߡ8|8b�!4E��CG��9+7�2��r�=;h��R~��,rU�˳8�t�Ã�]��*��SZ5����cЦgf��0
�l�>�G�̓��f�הR�1�@���i-�K}�k�<�s=��@)<�A��M�T�����^��CN�	�Ψr�Ɗ�W��=���}�2;-T�ґ�D�.�A�5�gݮ�l�������"�>Dd�aj���j��U�_0�!h���oț���x:n|q=(��N�
ӊ)�v�?1@.������i
���sp�!�r|j�N��DZ!�>�'[P�R�E �@wP�������:@��T�ث��V�H3<�p�C��S<X0 �(�����*��Y�a�������r�Z����x���sf�����}�\�i�w�nUH��3���J��N�C(���iG&���U�>)��3�����,/^4�ٷ~`��d�S���͇����-���X�R=$i��Q�<�2v�9@����'[�@�뎂KK�����1]g��ŞR$��C���c�� �\D�ߛ�dev�]��h��`�W4��-�� 
LТXo�F�K�%���`�r�C� 2�������Ow�졖�K�Ϫ|�͙^8Pf�o�7�d��i-��;M�nW���HR� (���O��wZs5��p⹽=>]��0�u��0E�n�ڷ������8[���̑����4t#�&][/胮=����1L��愽��b:u��Լh��ëdx�_RYs�.��~<>z��sz��`I�_���b��ʿ&U,?�	\��]���Z�ר!��\���EY�pRyuL��L'�Q��.�̚�󍃸��N�A�F���]#y׬p�0u�Ť��$�CAg��#~k��!<��D��<�%3���ǿ?A�Q��Z^K�z"������Րy���ݴ��ק�I��Ӽ0�X�#�w�. +��tl�l�č��xNGp��=M���A�Od?){n����b���Dll7#+��ң���8݈1����t������g?cWJѴ���y1J�M�|�������.Ǌz�&�3�p���~qW���Gb��x�C�1��&�;�#��^���gT��+Q����2�n�Yn�O����^E���S�ݵ\i:��%�����C�L+����R�r��Υ�Ɲe���<��cp7GE��zU�+r������]L/b���91^:�-p:�ߕGM����G��KlOzW����kB�����!̕�j"nlڒާ�ǪVF`N%L�����	ʇZ�s��9�-s�bbf^���d�HN�Js��D�(���&���?*�g��^ &"#�W�c����u�I�ܖ>~�8ҫ��o���|B!���� �%۴�n%��(�;E_��d�UU��㲣�+lȃA��$�x����_�	 ��#�g��2�����S}�G_Y��Y�;TW�A\đ�������]� 1�� �J3���C�:���8|4XK��5	�/��]O�.���Oy,�'��*kb��u�ح��O��0C��hVdt�!ii��U��ϳ�ӐT���A��0��3,�"y܆��6?��nV_�a��E�-nDN=��ve� oO�{_���Z�`��m����t��}�Wj��t���_
H#G�@8Kx3*�|<5������9-�փE"^���-�b�|�����/�b2N ��a�8j�{H�8}KR�/���]���'�f��#&�)��8vB���:�ey\�?J�ZHAϻ�F(|9 ��ψф��D�L�S���&���h<�=��M�>����[ihf\�s�O�_���������)'�˷���c�ld�nA$��lII�hW���C4S���B. ��@I(���R�/3B�TȂ�> ж֕�S����P�z<��f��q^r$C�l4!�c�E?Z�<;<�g�_j�
��!����/�o��]T�a:�P;dI����g���%��o�q�V�����% %��V�C}�Pk3�0i��QK}�]r����Ɨ�Gޏ��4��J�)Y�1��-f �/X�7;��v����� �?P%!/=������T�{>|94A���σ�(�v��Ɍv�w'-��Ȳ�R>t�MV��c
L����'�o�Jv��vޟ'��~�榫�'��I���#彉g�7��ЪW^Q��uL(v��G�����c��&�*�e_�$	s�Y6^
��ĥi�8sJ3�,3��#5b����������ǠCm8BH�9��^�mD`�s9�1	�c�C=ǥue�	��[�vsZ�,����5i.4ݽ���k�W:S��n����,��� �Ο8��M I)�;�8B&�Ip�]?Ou��1O����n6_Yk�=�IӻzT��V�-����q�1I��5w�W���r�=�?P1�!�i>g�1n�I��bW?'�OV\�
\���t��.��ήCX+!K��Y�j�Ǩ��K��9 �z7/$�<�u����\��%g�f��ثE*�{�.귷[�a�����C�]�^$:�_�`�6~
f�pŽ�Cx����RL�uC'��� n)qM���r*d5�9a��My?�Ή[ZY@�$�mM@�JuZ)�t'9���{���e�҅Ԅ[���;'��m?��A�]5uZ���5�1��Y��y��8�̲��
�o��w���F�CoM\?.�ۺ����C-���b:"m�\���4��#
�+Ey��k_ġ�*)�k%��qT�xt����-of{ų��T%wMU4W�p3�k�]X}����]t	}l4-���,W�C�К��a�fã�:���F�R$({�-/n!�G�Obݏ9}�,���R@���dM?S�C�k<i)W��_�GI��N�/��^����X������5U���؂ذFk|���2� erW&D�~��������Y%��y�As�ȋ���"I��,.5#/��;�*{�z=�=T�ۯ�K���B�Ys����;���E�Z;E$��b�k����ͯ�{ �7I���A�2���ʬ��Ԁ/'���OV;!˻�����՟�=;k\�vh�r�
@��wC:�>} �o<��Tq�ڤG~�U� K�Č�Q9WH��hx�'x�I�U�Y��I.�c��e�=�^�Fzj�^a�Dd�#�F �E�m���H����F�?�\�"�/:d7\9Jlpz頞�L����ա+���L��D�����l;D��mrjY��_�g�N�lnBJb5xi���Ϝ��������-�@�#}����D��M>�ۆ������M>���7�?:8�%�[Q�R&� X���w�m!1Ԉ�>]]c�}dk���UX)�)ɬ�������/h�L��,v���1(��&�zl���79ѳ1�m�j�M����x�W��{Ω\���yǍ"�F2��`�>V\�/b��֠QK�ț(
 -~�ݦ���;���ª�|��U/Pgf��1�� ~����nw'mKv�>�*�7�}lm�&&�v�¦��u��������i�߿ ���tM�J�5ϼ�|:����"L7��	�ʸ`h��E�De��	���i����7�����L2mYP�HlY�a"�@ I��;AR��qzٛ}�Ds���V�!�	 :Ҥ�si&-Ce��d�V���CP�p^��-/���Le����?F�`����NN64໼]sƨ�4��/�߸��q��?������$���9h�`�F7�&�j�c���Xuҟ��Q9�f�1��E#4l��0���?Hq:���p�]V�I*o5ݞ�~�y����F���D�	��iN%>�ZU�;t��.F��GE�'���l���'{�~���7�Ζ����V�ͽ�A �{SM���_�fI����p��8Պ��bM�1��o���h��*�h��.�Ļ��.ܿ���+2̀�q(܊`H틊�I��'z�m��,�o����1��<������(�O�pS�n]{���C/���x�={l�/J79N�cHk����n�����7⊧ �!�㫤zˋ�c��ʓ��`��6W$��[�{���I��qO�Ҿ��#M��9�d��xS�>/���Ŵ�]A!���&Ga�W�]��>���)_��e'�u�.{�<��L�c���7�mq@f��(�0d88�⻫�7$�� �B��8�iY�Ƅu�� ��;c8ƽ�.^��HY�a*�Ll_Y��2�Y��R�wt��7e�;+��k��*4
��������Э_V�\z��p���?�������A=0���o�3S��<9�[H�t�jΟ9cғ���ū^��r�gC�� ���i�\�7T�&��}��U�^�d�r���c�A����9�b�)j?>$��~e�;
��*��)�������GE���/T�f���"�p�ɗ�4?���i�����c�T�;�/���*j$c-4)�Tױ���P0e�����*�Q�"�o�DG�ZnqX��ś@Dv^&�[���#W�pR�����#��*oȘ���z+r�<�?SS#�X��3'?�wݰ^u�<��~_�"Cǃ���-�܇��6���`%
��E�3�V 4��𾪝|���|���9̌�5�݊{��XJ0�"��}�fӀ��/�}��)�k�H��5k�x��l�ߡ�����=6�K�4$)��{{&��1z�jC��*Ђ��e��&x�o�2�fc��j,&1�&�mn�2@`�Y�~��G��mI������d�h��=#�cuFC.`�����{��ҸP�&�a
�B�vM �e�Va���jaP@:4�]U�����e/С����o-���Ա6��b����Q_>۴�Y���e��6}3"�7��'�S���u�����>k�[3���U�<(=��fxl��8E��:�H���mD<� �Q��^8��Z�@`Q[Nغ��˸+�:a��k��
,��u��a_��	���B���Vf̶nwm���AӇ�a�ˆJ�	�������;�6u��k�?�Pq���X����a������V =o/����ѫ�w�Ĵ��/ȼ}wpi���S�ک�[c�K�eq��$�]���#�7m� H}�s[��72(k�#Ự���D���R�R��2�,�zbk-k��<~��|�1�'�1LG���w:E�u���J�S�O�; 9���a->��ͭ�X�[g���?��J����mzB&����Y
�vm�����3,,i(i5Bo:���oV�a�i��-S�m�~������(	�&�ka X�yUw�(����d�S�r�f�k^�D�/"-�!(�o�ٺ}�:��gd��.y@GO��p_�лfEJ5 �5�X-㧉R�Fb�.�z:^�C��KW ����Rp'��vO�l����f��D�/_D�]�	���9�4��z���O)�[�T�B��G������-��x�ѤLG'}v�C!�Ҭ�o�%.�W(3m$0P���&X��>;ǈ����Uܼ��I0�O�Q�W��ͭ׋c^ը޽7��VA����c8e�#�.���~.S:"���ɟ[���@/q��a��D_!�W���P�YO~��gW�c�b���1������ce��ؖ�T��vr�Z_�1Xc�um�V>i��^Y1�%x���Fg����aK|�&�]�C4������jG�^-v�s}�l���Y��)�8��'fuE��Vܮ�Uj��A�e�1fұ�������>�(&��ޕ,|�}��&t�����>���F/���J�#�f�S��(gK&������w�G�Aq,��U��@�@72�e�*��,X\u#�G��`.&��5ӴV;��W�C�f�����Vnɜ�+= �� -��?O�� n!�W/�e��.jPh�2��jp�
j�m�HE���\�I��B�͇��\{n�����ka���t];���V]����W� n���Ϝ!Hg��ٻ�]ڪ ��9��r餣�1�f�	Ηk]����+v��G6[�®���6zq�������ޥ.�ظRs����H���pDի�3�^;��#�q`e3{�!��B&J��:�BE<��!tDHtdb��@Fݛ��y�6b�t1���#����1H����Ȭ�&��w�,a! r�T�YY32���Mfq�?��P0��e�g��C���Rv3~��/��Үw�+�Y��U��G��1(���U����ě!�X.��xE��\�_�4�JjD������(�t^��gz�����3_�|�#�f���s%�����xV$â�"����c���=�	�,|��թ��@��M���p��Id�ԝFSU8ziDم���u%?dn�n�� <������-�;�|^���àX�vQƽz�J�8 D�DR4GM��٢�kw�+�r&.�NeV� x8Z�4_߂���+5�A[2� Tm�)�xr��+��Ӂ��"���$`����j���۬?Զ�C�PIc]�-'�#a���6yZg�����7�gV���А������^�!����0�؉[�$��{1�*����;�K���<=������u6���~s����V-�Ƒ�^#g}�s���A
+��"����q��F�z�i� �#V��n�LA�!��˳�D�����0��aW\�rb���<[���<8�W�%6G�#i3k�nW��QW���sjt����HdB(�n�#38��-�O04�ׄ���:TJ"^eƚ:�+���ص�ȸ'{_x"����-��X���h���ۑ@AKl��O�P�3�1X���� �mbtm�	j��^�@���ҁi)�N��t��c}�2�lU���q%XU�c�>�jG�L����?C�� ���:�GOq�!�3��$Y�q����m���!�YW%!]EC2�ԵL�A�J�`���!C5nQi�Fk�D�"i�8�i�^���Y��6	�vq������ߓ�\(��ag��ne$4�%�����&�/�J;�Y!%�ហ�q\p���]K떪���}�]��~�
�\bM�"@�7&�����h��::Q����x�U�eo�;�/T%��&��8ik���oE�w����� xF���e���D ���O�K�������eV��t�KBYT�݇���L�n)�W�@ˌ�c#p�U}�#~U�����V���.U{��8vs�7��(X^F�ʤ��)���1	�6N>�mJ�p.ڼ���(a���>�3PH��	VU��oW�f�֟".��	�]&4 �_�:�j�]�g�8�iF�<ۼ��O����f��]�3�f��耎2��tr�Ka�	K��5����ŗ�%4<�Er��3�r��u��O�L^�!}Y����Sq�%�R�&]��컪@ЫWw���tه�U@v�6YS(��&�����j��n�l�f�50n���dy���jp��I�t�n�G �뎭3N<>k�!w��MG/gjKsS�)���	UGt�N��7�h�x� �BKJv��N7M��AXx� ��l��)�.���
UK5>1�FޞNnSǚ�S{����j����9�x�]�|"*�2�IF[����.X S>�H�b�����n2>�6%l�Π(C��Vuec�W����� ��2�'Tկ*sL���E����kJ�cnٟ��� �v5�������{����N���K�oi���;���kH���)>j��j�Zw|��_'��frS|��/$�"�w�%6���[2m��i�Y�|
KS��V:1�0��Iuٲ	��d~���w2[�^���c�"���̶�жB�{�� ��wXn������wz���\i��p贶�>�C��wZv��$}�;�Y�e�)����ԩ��ܰ?�}�@;��_ ��Rr7}z[�5�!,�* ��[T��Ja"�ՅH�;0���f���~|q�8�/R�'���g��i����Y�r
�s����&�#7�RF6�2pՌX"~e?�z�+�z�[�}��Еk����Tʪ�7�nί�}�EV�?.<!t���y��?:�7X�8���{���X��%T{Y9	?��-^��]<G����TnfӊR�!��hd��TY���t�w.��ƅq�y�G��M1$5˶���4@����ȡ������:n3!��� �$��q�n'�$�`IM�ݯC�?˞��'�ߚI���P
E@���W�E��-ý�w��w)�C�W����D�W�}���2�vbL��<B��6��t��"��~��/���\N�̠7��� �}LHn�<B�d/O��#u� #O"%�ȟ$"Ky�m��m^�hh^�$\:��ݭ�h�y����d|���9�5���鹪Y�O�`����?���q$���gC�yY�e�Nc_՚�,^�����'1����$����L�|�A+Cd�|	Nl�n��ʽ�ó6x�����V?�Y�T<*{��`(L�o;|�����biy�L��vڭ�������߄P��>>�_J����Kx��Tt��<�loF�v����q6{S1�����Z�K�4�-�~I	�)�-8�F���|u��Y���S0zC�&)������2�^��ٺ;���
�屹�7���Q�O��ۖ��K�s����ZIV`C�Ц�@��d,CT�����$~O�@|��=-GxY`�ϑ�Mj̙��o7}T�'�Aze6�����,B��
A��E���||��_E[���B���[}�PbO����=�# �?{s}�l�qʿ�薛��ʊ8[)o�I��� r�Ѷs?�h�K&?�K6�Dg�9Dj���h锶z���so T�ZS����x+�?!�{!��Kz�{�(
�u��<�*��Z�Ka4y�~�����fO�v�X����İ#�J���!�І*و�&P�z���(�Kb)�)t�N�Y��Bo3�o�r��N@4|��-M+�'-�<�m?qT<U�Q��l�7u)�Ɉ!̻�5¡䩲Y�{ ��y�znaG6	�qP�~Xh���6u�;W螘��A6S$�l=�B�o�-S���<�Wr��̚[� �$hh�א�5:&���<w�A�$�>I~�)g�:Ȅ쿝t�}؈h�f��w��P�<��I�2��3|�*!ǥ��� ���L���x��ё-�tb�鍄��P8Y96�< V�]�*A)/g�IiL{�N���ht �]�� Ш��Lx̪�1�٫l�M��<�y�D��7�x(�城��h��$��C4:���~�4����
��Z��T�l������{#2i*x�8��P��	��M�ys�Hj/����7ۗ�Gڕ�O���,T0/�$�L�֬��zd�XX�]�Z�S�������HK=��?�E�������;#�o�r��N���Ә�/2��4�y���� (���ظc�$`�ژc9�;��?�WB��6|�oΆ�KAb��}~ш�X+T�E�%Y���B��7rc�yp�Xp/���Ab�{�[�w>�L��k9Y�R�K[�lH *Z�ܛ{�7T�x�(�E�<^'A�k���.�ח��DDi0���3�}H\TûݍrnK>�j޳.a�@Ex����)�e?5>ռǻ�6�T�Z�d�����6d�*kS�Ps�.��L�"����S��SLO��l@��dwT����e�����{)i'�hC��Q�YP8N�)?y������P#`i����������͹i`_�(m%*���!���N@�|f�o�Q���/�U WIjeS+�ֵ4g$�n(E��RJ���3�*�?���y�����_�P�lh٤8x4�wܓY��-���h=��p,
�b�-��d��:f��:�B�	,�j�^v9`��(1׈���Z��{V7 ��9l��m��ӍsI�V
��!�;�\�T��ޕ!f��'O����I�<V���6��p%��(Y7d�,d��O�6�׸��Գ��7��TS�5\��_�t'�o}�F�m��?���U�o���h�R�\��y?_�3E
��І�)�^��Ҳ���q$�+�@�.��[*��oZ.b;��ч����y��x
�~0���o�v�Fww��'pT��c�ʶ�Xx�X_�xĥ=�N�(\��(y=cD ����	�v[�n�W�F���J̩1a�gi��)�S�7�Fw����Fv�)�R[����p݅�xN�z"����0£�D�W~�m�DJ<�V�� 3Y�U�H.�s����	~?�kTZt������p����c,�$:��nJ��I�z%�o��v| ��p_ӹɍ
ľ�u�����r��)�R��//t$�,5�?������0���A�.�H��vd��v���H��)D�½I�������7�o��n$X�*Jc�C>�O�S��^�G����O��o��4y�L������sA�����q��F�5�bG���~\�I����V�>���!�U$�͜��iq�Kg{��7�pAq�����u��'Fu:A���c�q�8��j��-��>;�"jLxH�G= �Yn˜�4q `���-�0(8��ۦr��F>S�Ȗ;C������W�����@Ï ҒD���Ő�Ь
���;;M�MM���*���
Dx���Ame�A���LM�Rq!.���9N���o;l��e�P�r�Jݳ:�Y}�Y\ܑ�|h��#[�d�H38��ّ��0�뺏J�>GGq����?4"|�j\�"�ҸLƌZ��n�F��n'.<[1���j�2���s�� ����;���t�˷���2cv��L�/ʅ�ZIe1�����/\�CEݫZ$�I�1`��A�w�ݶ׋'�i4t���f���BD,��f��(c�pb��N֏L��'�T���Uq-�W�&уPW���v�)W�:v٤A�`�1v�,`�*0s�ļVC:f�8L�Z#O����ε�����	���$B/�{I�����Z�QTz6]�o6z�]�5B�V�G�q;""�L�)B�2s�o��U�X�s���K�j�c��
�N��18 �OU���~ܽF��0���(��]���͆�M��]��u=a�Jy���`qҕ��{Ӫ!������z�؃��u,�W��	��BvK�Ʌ�M��z�Čޏ<�����Y���<��'C��_�y��tn�+{�cS�V���q�(qj�sv#Ѿ���x+��a�Ɓ߶���ѳ�C��Hk�T6� �U�����#���7jDsĲ��1&�.��}R8��g�є��/���|�����P����cp^g����azMF��I	D,�Ai�{�s�7OA�x���
�M2Y��ϓ�X����|�)��x�t_�l��?�'	��
q�N+8��ߚz��)���gU�p�'C�,�GW���i:�0S�����r��.��Q� �_��(����Y�7_�d���Es�W9Čᨐ�2�%[נ�	"f)��N��i����ծ���@u@֚.0˹I�+j��� ^�<HO�+P�����WlwCA��y�k,�@y@�k��UI{��f�X^�
�vaK��>!�A�u�vA�%]V��w�"���ǀ{.�k�?��XE�A�q�g"�p��5 ��j�����(�.��QW=�F��!���k�7
�ϵ����j|���ޥ�A4��
���x��b�<�Zʸ[[\!W C�#���$(�`c�����	��\�vg�h��i�� ��tA"��0�g������*��ƽ���N(
��Nf�X�{7k��Ey8#~T��c%+��`k�xĜ��Ϥփp���
:'b��)����Wk<%V���u���ND�CE~���?K�%��&P?X�Yh�[�Q�B�>��%Țx�6����<uz=��{f��*��Fz��)��S����y��W���<2-�1���A�-31 �<Ӑ[_�b���YV5�ȡS�h��{��e�w>P%YqkS��Tզj�j90��Z��/&�K�&܀�~�1G��_�����P�Ns ���m�ڈ=j���fDz#��$����p�t �?���=��@�5/���X�;)�n+Zӆ�,�Zn ��n��X}Fz�C�	�#�L-:�θ[>F� ��5�#�~��y9J���r�cn�9@����7TA1P�����8�f�2sܣb��J�o��?�5^���b���;����<ٙ�@�T�謓C���:�J�Fv�9"��y.��uwBcw���B�V�x�
hhմ���.l�y�]B���y>��<�6���6z��1�y��.�*�}P���	��Q�S�����.�m���<�'�\X���՝t���;m��ngE��m()Ū�H`�����!�K)�Y�w�xU�IKג^H��bRS��Lj��5��g�3bH�S[�U9֟�6��6���s����6��"5��LT��a	3M�*a���\M�-�Y���h�?���
j%Q�-�$� 5��n�f������q�K���Ӎ�QW⹚f�i������z�Q@}��B��b�n�A$��׍)�ހ��-a���^��?���W��&����BzCHF`y���=f)�y�kq*��|Y�ԍ{��!c��m�y8�l��%V�w;P��TD��7��-��f���OL��g�����(��[ǩ&�s5(-]g8 F}Y��-w��v�E��GF7��G��e�q�7��n;���h!9h�#���w�U↞��USRz� �M����]<���Up���5K�9"� ��)��-���<p�7�X�ڗL�~-�5I&?��	�9ڦ�w����C�u}TW�ɏՙ��a͆?�=��U�*�B��0���?d	�Ȏ�`uf�;:�!5��3M|�T���Wc]֏4�}�-��[�o!A��Ba���ݜ*����XEd;�A6�����r�jwX���^ҷ���i�x*i�?kA��wg�A��
�%.��N^����H���%]��3�!`�F���w=�u5v{�����N��{��䒠?�a�G/q��B�nt6��^�k���cV�~"�L?�rnZQ��I2R>��I��Mxz�#�Z��=�\�U����ӓ9A��^�����H�>�|s�0+��oJ�O*w~�[�b����lԛj�E���6*�ŸIf�V��,i2�*����Ek�z�e�ЗAU�k�k6~� <-���)Ok���+UM�!9�muf����Q،�%K���K�@�0ŧ|����D�/�j7�&g� uIv=�d�M�X8)9���jJü�l=Lr)ɽ���WS�e���^w�x�D���\2��}�4֣�����
�� �{ϓ=�?�&Һ(c[]��jk�/�+s ��^[
��[5�w����"d�~�U�<���P��O]ׂ�����(@�̎�t�RT ����f��'��)̟��80���A)�������5�ˠ��^Q1�|��>$� ��<��x�0�X�*�v�6�I�F��*É��/���1,�p���<�&t1�L�~"�m��~h�$���Z ��$�̶����p��������v+tKQa�=�Q�p��Se�
� ���ATq�4��O/�K�HQ�&�L�N�_ru���@�7\��_9w�}��d����/>����OY;̿�b��4iW5'!^y����)i�ߗp%׉y��+*���]-9Z��`�Q�'���K��P��i+E<�u�n��+�i%,�-��0
I!��5k�'f��%���Oȑ�7���3"�� eן�틭����!R�����	o	zk�%ƩA�x�mD�x�v�鉋|썂��[
���vˁ3
��C!���i|��[�Sx�e�ΡD���QxU�e8�����(o�`���ë��ر4������m�-���"�	� j��P�71'x�(�?��%�KcsR߉Q@�<TW�q$��}}�i�eK8W�V���%uy ��n��m���CHzo���g��w5�R�gAa���ҪxrRn��eې�n�<�j���
$��ߗ��_=� ���a�D7.��mZBE�
V�N����s�hm��o[��|����e$^R7���@��Qv�:���5�(p����0��n!f��[OPY������$4���袋�8�bB�|����U�Y��m�����"��Gc}�Є1ǩ��y�����/x��#�<�"�dA�/919��@݄&n&)��J�$��!B��@�Aa9��8^(��b��(	!O�`n?���3�]�Q�2����H��"+TY̮"|�j?�0��w�{���9��,��~��X�P4(���dG	q���?�U�\p�C�3J��a��Gʾ�>u.A.�-��>F���h���&�c�"sY����d`�g`�3�<�I��׽Qb`�$',�����މ��y��{�����#�����ݛ�OeT�揯g�)�(��{G��︗��V���Rw���AS�}g,7���˾��v������Z���6$I���IV�ۥu��.9gU�VS~�����t�j鶍�ثF ��s{�����f>�ŀ�R���@vB��}ҡF��Rh������ж���GFiH{����l�Xb�͏�i��a�LVP6�QB�	��&�W�s�����9��`Α�I�|�~ 0%��e���
s
/������Os鐚�9�j��$�	���q�k_udW���v�0�⭜~�ܢ�٧&of� ݟ���(z���l�qy���	hQ��B�E�D���mK�ɧ�
f�U�:2`�2�� �"��j�k��g0:�k4\v���o"mZzx*%�ۿ'p FE�����|=�+-C�"�q5�Y�QV��`
��˩�l>nE�ɨ�Ƽ �-��d_���}7�&zR�Jy�@	ȱ�~�����zkH�QLL������	<$S�C��,�3�N��y���IP���!�5�i\g�������3�p�X��X�!�#`s�o���R��L��,�s��-(�4���m)�Ĺ�M��Q3�A��Aޯ��&��>2H7�`��<i���!u���|��{�"i.cr)*����-j1&iZ���-��>�l�y� @H�(�ٌ�a���q`��[q����+�6�m�M�컩�;�a�kz���lTu���ג�\�R`�����q��Js���|�{�)�d<�3����뺩i`Qv��{�ǝD�<�r��W�Ն�Sε���ib���:$T����C|�~��F�M�򷋽��ؗH_��9����M��5#�[G�ywj�>��F�8��G�t?�U,�g��4@���XA�
-�!�qH��&��P5��pÍ����"��3�8�t:�>El���e��������Yf]��f[����F��z���� QdȜ4E�b�b���ϰM�s��N�<�:e� /H���ZH���z� �܉*j���Fm���$,�[ȼ�� �.#���n���{���H��P����Ez|��`��|�7�D��%��+�d�7]�\�0�
������@�	t�5��2J{ӷ��t �e)k��H���ӏ��W�j0<D>`�^�o'���h[	��{�	>mL��Ļ;�^A�q15�kS��#�`������MO���+�Өw��=S��r�g���)wۃ����k�
�����(��z�g��tA��r��� ���#�?�/��i
~e�d��w)4�e�?s��x�Zy�*m�l�g"m�H�ˇ�kNyON�B�^��/��(��ED�'}t ߯-ZRI�F�L�4hф"ڸ���n�K��	���}�A��J�|���*	saDL'N��B8�f0QQ�(HЛ�g���{-Y:�v�	�w%b��M���
����_��4 ���}3��t������u�n͚�����KH6�Th�L��� �`�:�EE�f� �uw.wn�e��q�X|KUZ����M��|�p�6"x�]���x�u1��iT�ߑ���"祥Fp	e4��>@?��A��$���!����ЭL$-s[�������� �I_TDb��-����x��ų1�x��ן@ދ��K��Z���E�%R�@���2	��A[�}���5�x2�� Aṯ�V/?З�NX���O�j%JiU=���5��~	2Q���+��?u���h(��"�\��|E���bc��1��U,#�@����TJ�,��4`�������b�p�Y08"H���$E�������O�FV�䧴��8����f�Ao_��&�p����%O� 󐌢��F��	�(⼶;[:��4%�k���a����Iç����NZ�qU��]����卶?��=�=���t����KaRP�/S��Ga	����i/����k芵818��zh��nW�>Ѭ2��]�6?:Iw�Yxn!�g]��	�="�q�"�U*�?��,��/�_�Sj�%�$x�[׉1W��n�嫥�΄[�E>$8�S���������@&ofZ��1�nN�g����s����`A�܌=+GK�|��#���.h�Dܺ͊�4��N�E�#Mar���T2�S���7�(�H0P��A�4���z�F�[���j�����$'�O"��ň2�a���?���˰ �>�$U�ȯDO�{*�^�aL6�"i�r������0�3�k"ؼ�u	� ����`!�cj�F�/uy�D���d�Z=ܝQ�U���(Ѩݦy��������փ|�-�!�xo��O�z �Qo۬���n�Z@�b���'R�Q��
)<���I�?�-9@J�Z=�K EKV�_y�=U>�2�nh�r$,V{�s���
z��= $�$j�J�<�Ht�g�-V[��֋�-��u	@<fR+D�n"V9��60����}�i����N�^(�ۚ����3�-ET,��&ָ�d��s�˲��/H���Ng]�W]o�r�
��wa��,|ϱ�ck��E#��&ن��w�QV��q� �j�Fm�C$��,���WI��ԙ}�L� �S�ְ�$t�,�_��DÃ�O�tb�OujL��Ii-�n��t���zT�4R �Ҵ;r����Yv�9Phǫ��z_�����V�Ƚ������#Û�/_-�7My�0؆�(%��?�.`��lw����>4��?4�$A��W� �?�Ny��9�� ��^���7;�_-���˔��?����!�$��'��aޑ�#�����2
�~PW^�e���&�a!��qmy��f��Qwl��ݥ ѶRf�L9���3���A!sW����Y.���0	�E����Z�f�X�و�D�l�+�E�k���U\��9,���-�*ȉH}<�M�2�����8u�q����v���헤L��8Nk9��3�-�bm��R��@��֛S�/�v��o�ۭg�ע��:b����Y[��<rq���h��s}��@	e��&�?�u5jA�F�j z�0��)���gvZ��Y�2#
����T�'�ѫ�K��V�;��|��mE):CҰ� X�mo v 
��|d®-&�缀ĔS��7�[Ui�U�ѿHȷoĸ[E��u�רZS�U�'2!I)��(������E<�T��HAVC��[����y��^���`������U0�_�,�-��)��r@��s}X�t���z�d~�<����L~��>��k�J"���ݘO�u�!�&D���dږ#�c"ɵ��u?�+�
\�r/�;���pkEvԬO��0�EeN���c[��O���ɱb���7�}ۻ�	�,.'sI�c�G$��!��Xm�!���]-U	��8�K�{Ԩ�N��ۏ &����U������ﯨ�?�Å�p����z%~j���}�l�#?�dա���i�+����?�X
0|>���9ڪYnr�<s皷5iM�Y����֪�s�y`�o�K��3��l��bn\�ʪ!&؁gl��ڽ���;���O�y��A� N���+�b�	�`���5�:��>��<h��,���꣞Z��B*�瓺u�q�ACRiuA%�%ٗ󔞦�����-j0C,ft�2�#�!x��Y*u�nF )�QnKt�9���Ќ��*�f�Q�Z����������hYv7F�ټ���T���O�K�mt�����K��q>�L������/0=N����+����nd$j�ӵ�0�#4E�L�8C#�9DM�k�D���&��E��2�+J��RDs��"nl���J�u�y�q+�]�\]��H��卶�V�i�.s�<1r���"��t�f?*\ ڳc����9-�>����[�hQ|���1��V��<�D�_o�h˅-o�ǂ.�U6�2i.�g��
	�ڹ��:�=+>�+�qa�����f$O��7�0�sM�7������j���v��p}p�H��0��'#3K��`1�/d'fzQCv	�@�4���&v�v?��4�w+wQ����h�ż�r�Ёe���#:���tA���|����n�� �6����yi��X[~���f�x"ij����z4�iR��m9�ð�O�X�?�M��a�ч����fd���W����L �����ŊM��2�����Sߍ�B5il.��0�5�_�=F�vE� `z�2C��Z0�A�X�:U1��^�����Xc�>أU�vƣ>/��>�7yZ=C���/�&/���]l
�F�)��Mw�8us���j�#�ρ)��_c��k�'���vCE\�~�X��i��i�`�^"s�
Q�:9�忿͔���o<O�v�������V�Y+2|��>Ot�(!+�Kǿ���n�r������R^[�~ȌvY	���4��L�k�q먉��$V_�a�Q�T�+n�E'�cl�T�]�4s�e����(�nN�"�W�\I���O> I�a���Ȉt���m�0?�l� 8Jӈ0�Jm[�+Un��{�lM�ށ7��8���V5f:2��=TRyd���#�E��Sr� �/4�^�c"�� "Ҟ�ݗ;O�h���
���B�7��dݘ�\i����N1�e�
�S��79<x��������a �`.�/�2�mY���J<���B3m���Tz�sT�{Z���Y�F�ÿ��ȳ����ST|!����<bv�,NJAq�*Gc����$�z�wb	.�X�PI��pe7t"h��	b��!ǂWsr�����'���}�CYǬ]�Ӿe:W��ч�@p�t�!U�DE����|o���	5țI��m��wD�UU鞍!j����@#�Oo��)�&6�\�{��-��L� m���7�H���<1���>���7n����/�|S_Qh ��I4�̩��}��/`	V\g{��L7����c���³=l`��^����&7�i�␭8��)R̜<BY��EI�vSfn����"	9�.��?�feB~AT�>�n�L�n_�;G��	2\�`{���K�syż����9$�����icP6��!l��1P���̰�ʌt���y�+���٠�q� y���Bg�-!w��5���s��cf*t�	��ē�HX�^Z֏�l�bm�	"1Q���>w�af,=tAHq�����ނaX�0me<"#���i���b%��$�6�2�X�"�o
f�EG���s2#M�[��j������w��g�"�/�=~�~]L_c��ez���SV��a��x0u3�1W�+�=e�̋�-n��)�5�RW�2W]��`F�S��ЉTu�Q�A&�����d�p�<�L�����Ó���|;�8���T�>ZT8?�d����w�>�.CnT�z>��<S��<�Gq�F�(�h���j�ki�ȋR��m��	�ɽm��>�&��:��(M9B�sHW&l�z���ͺ��� XUA�&^DZz�آ���2���Kl�M� �Q��d
���l�l�̝)��`����uޮ��L�	mU��4�����	�3	�h>�c�֍��I�Z�lzK5���>n@���zBUЃ05ȦX�1��Ģ�I����3��9���{��^�-��y\~2�_��\T�&@�R�)��2�8�C�f�쵬eHuPc����[:����nMg��TJm~Q����,W�!X-y2���P�W9|����`��g��b�`�[p2\�����Fr}����Ҳ�s �f�Č�h��v�S�x?o�W�pk�>��R��b��~$��B`�З��4�B:�i���GQ ���l�p*R�#�kt����>LH� �Q�I��cj!tf�7�(�~�פּR�꿢�$R`��*GܴC_��e�Hb���R�-�LW<Z���J�Κ#��{��:!��'�s�F6���	�n�aA��m2��]��9;y(�W���ϯ� o'����s��!�����*c�u�hR^��.�����R\w��ϗjs��{A��������G��"F�	���yO�x�նr��VDN*U�@��d�C�e�bIԞt�w¦�Fp'l�y��G�~ٴ�{�V֠w:C�U}����$�Ȃ��x�8`fh�ҏI،8?d]�zK�G0M���Y����eup����k������J3����*�&VH_��L|�W%�m@M�ŏ^<�]H�1�P�d�"Հˬk3�l��HZI�q�I*&���H|U�uA>m��7���]�r?���YWB�Z�M�o��gH���l@��U���aF�P��1�2�x�X�Y@�ˇG��x����bQt�#'�����"ʿ�@�����埣�Q)OR>EԊ
��S�E�5�''��Vuş2Qp����R������I }�����b)��\R-���[ձ�.�i�ǁ��q�&� ���Ӱ�)H?$@z����/�S�e#j���J�H��Hk��c"�W"��ۓ���pHd�z�+�m�,0�Z�׀AGt�kǎJUz��4a�zi��{����� ����E�Z총ߏ�^944�X��l�k[ ����9�zC9ܫ��݈lg����rv��H�������Zt��х�	���)hyj-�:���TĎ^�5�<Q��D�a) �ۿ�0�rִ!��⡴�>�G.n�0Zk���%Fj.U� ��1:���w��۸�hf��FP��ȰÎ9���q?�h5��原j�I��8�˫Q���t��T_Dc�틞�Urf=��گ�9��i&��E�E�w8�����ձ�����rF��ϡ��p�Έp��v�Г��'n�J;��Yz�g8���c��H�����.@����5H���z���i����W��\�R!��m�҇�@v΢���a����:Sy.���$/0N�7rf!d�1�=bx3����B��L�7�#"קK��D\8zg�/�m�Q{��4G�O����05���PM_'+�1� �W��a���3�1{e�F?���N�)h	p2�*�Dm�W@�������)".���v|�D�f,�3.܇���'���`u�����7`D�y�w>� 9m��6�G��\Pxʐ�S��b�L�(*TlX���]�BA�Do*�Z�<�'
�Ke�ozgۦ]�N�#�=��4�#���t�x�a����'o�TTf�P-�;�rD�STo(����ecA'$m]*?���i|���f۱|�~�.���U?VS%���m�9��U,��}�A5�]�1IQ�
���B��)/I]�E�Q�J�}���	��W8��N{re󧱩��|\��A�T�B��@r/�m�]�ٟym]h��Y�m�[W]���0�zt���`��*�����#У�-��o��U^Y����+r���o:��[Od��pGN����f��ϥ�4d��Aʴ��{��*r*����U��7�Vùi���[) 3t=�H����L��!.�����	S��i���s
�+�E̰%\~jOC9Gw6s�+�_�8���4|b�=�ިD��Y�6!b,+}��?��� g�D,*YE�!��E.����q��1	�ZQ�p#v"�*N\��zܼ�7�f"Y���� ��e���[검S�瑒+�nz����8`7�S��(�"�Y]�C�_�$�/9p��W��0�L�áp��߉"E�����VO@���'t�:���>�|k�q�4��1#D4d�
Z)(�nڏ!̀C����v�zgZ�X���ϩ�ۗ�<��U��_��Õ!;�p�n����-�$f�b׆Z����4M��^���ZEv!�R�R��T���T��N�e��1�?7���K y�u�M/Bտ:	�ڔ]Q/�	j��T_�X�eJ`u�40>;��d�j
�m�L ��<�.�gyLȍ{��6q�`q�J]��¹�'j��q9�lWª �0����-�:�p�r꽽M���u+���q��<��jK��Q� �\~�}� ��_j�O�]�63�0�2΅0�A5�� ��Dw�>�;���[+mw�������68�@	�l�� ��u�1=@59�g�|9s^�r�k��	��`?�W5�]T����K�SPz�;kQ���K&���Y��N\|W��}-2{����k�g$�嘊��aͩv�e�A�%y�(62�l��ю�4��L�6(��H���I�L��m��������As��;1���9��`	�G���m컭֮@�R�����IN�am�}ˌ�To��F3��"5%�A��w�p+��A������m��nՆ��x=y`t*�ƀ 	�U@j<㾘`u*�튶BbN��σ��R1�dٝD �2�u�� )6(��
:�
�T̽�t�E�H`d�lM���J��_�iMl��7�:ż5ѳ��>��#��Q���r���G0��h����`��!�s��4�9�#����̫�z`�G��l��p��̆�q ���?a��� ��}Zk������>�)U��O4������|�I�8�)�3�I�paj�c���O�z���m-=G���ݛ��N|K�HO��7�B!/�A�G$2ۂ��?JZkM���9���9���b7�ui,nĨ}c��0J�ΡE����g$��n ߯)������T�1���
���>��0~����jt6���ޟ�3��s��]�qP�F�D�<�E�U���𠘘.��Nr>�O����$>��2��s녻���H�/4��&�>�<���+s���s�j��b�l�}��x�~��.i0 ��ƍOo&^ٙWv��ʇ��5����]L��pU���a�)E�P'�*�����G��̄�\�q�-gv��.��������� l�8��*iH�k�RU�b׾�-'%��8� \B�z���*�@,  7��l�U^M��JkV|Ϛ3����{�2�¯�
�������^.�8/?���D�t�́��Vr�Fr&�E�����OꊮC��h�;߳tN� �=�@�)��;eJ���Ã�9���>_I��<�/I}-�FCU�[ʍ�[�^�d��nh�(a��fc���|F>��HXMr�H;��f�j�t��]�XY`�����=�$�5�<�H��6}��X�� Yo�3E�5�p�N|8��x��T�*p|��L�8~�����/�b��p7��E�d͎�;y��F�k�t?�U��\Zy�x��FM�a�'�~�v��v��:���I�k����y�5%B��ᚁ("<<{x��()Uy�ˍ� ��}��4�3aM"��N�@��]ٛ0M�������9�/B����c*'�S��^��zPf9��|��1���ψ���,=��V�xU���V�o��O)A<��KJ�f�������m���_����W�O��:�&��������-W`^q[���!�w�j»�2F� q��wX�X�Oݠ"�_�^N=,l}����b&x�p'��ԕ�K�T`j5�]�ƪ����v�V�T�^�W� �ώZgtI3y��8�.�1����pN�?��|q-�UG��uH`Yƣ ��}I!|�G�Jwfw�wԑ�,��y��s��%�ۮ%rG�.��rj&�	���K"`]<)G������#�EWx	��|��f�1���q�}�t7�K��1)�)'��ro�y������҂�k�M���l�9�t��$���w\��D���8uvH�mPS\w�lE����Ĵ��]ML���EzZ�ݑ6�o{2v��VS��u�VO_�y)U����;�.c ���{ב�=b��l%��ED�;��dw�wt���sm�R�߫�z����Bƚ�iC�j�*X�J�GW���ӜK-*��hRs#�郅��^�H3p8�J�.��Ň���̒P?�2��b�������_R��=���_m2�D��-Eg�+7�����O@���HH��_���io!�)[&���F-��8�_�RY����Y�����+�tɤ�A�-wn�SùH���c�I5�2����c�	_�݊��2>�XR���^��.Q`�}m=}>���;�����׶t:�����2��?\�1���3�a�-�������H�z!6XW4���%�I`x�Gcф�kb�3
ߐ�4�1��ȃ('�%�0A���;}�e�D�W�(�.%�9�QR�sKG!5�;��"�ђ.����`��{���[|� 2�y�$����D.�z�k y_��a3�̌S)ȅ�F��s[�VE����8���0�Q����i)��8�ˌ91)���F�P��%]t��(���ج"PP6�~O��U�T=VL0��ߪޖ���t��V|����'�<�@�r Lю��� K^ZpHHc��8kwƴ�'-�d?v�c�S9�ڠ�0W��5oO�	���'���ԯ9���*�B��f��ȵj\;�� �1e�ˢR�Ө@�e�-��ۍG���6����#�R�U�fk�I�:6�`�Zn��6��2�lR-�ݔ�����S�Rr��m<��$��,u|d҇Fҽ^	1knj�(W{fbF�%�C���k�Rs%Z���}Sв�~q%G�Zw���e�u1��(=S�ߠ���HNU�����_0( ��-$~���r19B�����X}b��ͧ����:��b�6�Տkݚ��?2 W���>n!V�.;�a{��j��&|�.��`��f8�̔��)�~�`$��~*��9��
dq�w�g�!P�^ j�<�;�ҙTƹ��@آGz�)Ɲ饱nR�˃c���j2�����T1Ǵ����AbCzux�� *U�|(�I�.�wQ^��c�Y�Y�� ����l�8sO�v]�v7@�U#v=W)�`��Pu���n��5Y,6�0z�옘{�2:p&�sWBu(��5>��J���	�|{��ˠT<�?��)DE������.�+P����6��<J��o%��.ǯ*�d��c�;x�G�MծI>�#\��>25���!x�-ӆ���_9����3����>G#��
ٕ�q9��[^��:����(���6�
�(b����A\�����Cݓ���0�C�Ff�Ql�6q� uu�<���{w��%�+of���J V�A@&�C�j+�D���`M$	�=�"'�԰�<V��\>*ѡõ�!�1n��F�!��n>=�!Հk�w�-ˌ߇*Q�}(2܂�����fS�C�"o��YEq8]���7)�uG� pw�8��)'##2G���^�e���J��:��\��������?\�gr���M�1��B�KhuSD��X�򩬼Ju���kP݉��ap�ѓ��5+c��8��{B�>,.*�B�����ߗ�{Lr`��/:��������݋*-«�\� D2�P���a���$lO���Zݑ���P%)�U��yݞ����u�c���\����KR�R�Mu��Ҏ�VGcw��9����$6�>��,���=�`}������q��t�Y��5%L��+�}��7g��X ,s"K��d�۹�A���(C@B�� �;�&�q�_�Ix�Y��u� ��\�P8r�P}t&��8ӗ��������K%02�D����a�;�Wx�)�q�4�����pT���v��[�VS��,���]4�Y^䗏ۍ��ARy_)h�ć:A"咍֔��9n��v}�ߎ���!�%��C���Z4������M�e��OSu�o���u"��1��մ�!�6��оwP�����!�;��0*�L�zѠF���Lb�$NT3J�_x����f}��oV�cI�I٭��qPŃch�`jg��Fs`����a��>���bZ���IK���&X�"�%
N���D��zt7����x�)&��P72�
�U����^�|���,RΪ@c������Q�\���>��;�ì�DV�i~����44���%�=(N1�ք:f<1���uLکFJ��<���&��W�g�΅O�XOk�s��Xe\���=���qB��w��;g�L���,c|@��.�N��oׂbG�R���"���lv��u�~_�+�z���Ïyo��TH���	�b��h���r%�9R~���p����Л�)�΂.�^�=q�Z��W,��z3u�Ⱑ��nS �Ͼ�08��x�ߗ�ȥ%��z��%`%2l��U8֍�7iL <�.����B����ܟ�|��jua�S�ڒ�m}�o�����V�\I{KK��Po&z���K�<�q�aN�G�G�Y+�~����[F�tk	92AK՛��ty�)��Q�p��Jp��HX]$F��`-���7In�\���d�g��V��H�R۽Q=\f9���r����D��k�y7��N
�}��rE��p��(b�����2d�X+4�o�f�AmM0Whܪw{�0^.�+��,�9��{EO_VC��ٗE5�H�Pe��� (���Fx�u^��k��{�d��^h��)����H8��{�l�ͧ�A���kQ$n��Uj���ժ�鱵�'�i�Q��}��邷���/E;`�U����\���t3�#�Mi�n���Zؖti�Ns��}�Q�վ�.:jI�bYKA
�%��>�mF����K�恳�����h���@� =a=
��M�)��=cY"S���)�Ăʟ'6�f��߼�<̔)�𸹅��5���bId������KG��yI��3t�sx��ϵ�5���f�#�㵝��A�� @8N��M��e�@��խy-G��v�˷�}%�'��xY8l�l�Icu6� ص��R�6!��
%O�`��&-8�=��>��*v��a�V��|����/�9wl�;�`J�#!������(WrK�U��푆)A����SH�Yc��x���A��s�=�%��(�uς/���=;���R5�6,�{��`d��j���*@�!�8���5<����@|�W3�;[`�_qQ/��;�|ڎ��EQ(,fm/�R�D|
�<���%���o0"�� OG�I�=�#v�^"�'R��{=/L�Ͳ��`���}n�ia\�)�B���%�}�lx�����{b����Q���n�:�s�¨PX���Gj
 >O��R� �:��߄f �v����:cs��^��)�����A����y����R����ʐ�
+|>�[�7�)�=���va&Z����|����:L���~=��Z>}K�B��p��]n�$���C>2ao4M�l���pC¤�9/C�q�_�G�ڊx��Q�~���I�Lݴ%N �z1��8c���e��x�R)��'Q$�E쑗�rJ5Rg���������p���t�6�N�S����y�KX�@��(E7.D0���K�rZ�5��Z�^��SE����Me�-l�1-�����}�]WP��7��_����B4�+���.D��Q_�'%�d����"4�Xoϙ7D��v�����0��}O=Č}3C<�/�(�;3BrP?�ξ��b9�J����cXQ�������x��d�E��"��h$�x�y���@Р6��<��~��!���A�Ʀ¿&�qu�NDV=Ձ������%�? n�� j�D��.��=��ʱ<��`�ĦV(FZ�a\�������ai��M ����w?�a�����? �̀������8��ږ�"�_�o
%Ä���W���+������i!�@�2^��X���$��Bn�}E]�
��ь��I�����: ��V��0�����7����ލ�kHXė��v	���"��8��cL۔`3m�&����ZየWcT��X:��?shc-{��s����-��;(\�h8��qT���`i"w5pb:��i�ٜ\Tv���.$�p��NO�x
4?�%"�yneӪ0@�V��,���^FQ�p����������LK��b�'��Av�#����HL�ǃ��X8���߷;�l�yK�zR�b8U��ׄ��s�����d3
���ۮ���l4��B<�~��U�Yja�{/l�e:���[k!uth�W+�w��	��?	���R^ܫm:�T��Lp�"��&�]������x�3���@�<zD��6z gSG�#،�b��)�h�P6�b�����վ�� Ou%:gWE��:���0v+���� ���ކ�bQ{E��Z����CX 	&��H���p!��#��ꪋK���ߧi��{tCؔD��U���E�_{�Sn��&���z���R�ƄW�'u�<�u�p��zC��Ҷ��ŝ;�恼ܮ���l��6�:�O���L�j�v!��г,�2HÅ�����(z�"�]؉�\6[�{Q��N��6#F(��=YQ 	A�D�;���!�V�55�{��6j�L�r�sG�՛�逍_�ܴ���۾�8�`�ݭ�G;a�d;�^)
��b��Q�uc���Y`����f���#*��шP�kD�h񘰉��V������O�����-g�.��#Y�d����~X���*nt�ukI��_tG=/�j�D�^�ù�Z���pɹ�=�N�Rʽ�9�P��������2�+Wvi�7����i�O	[��0vZ�p!B>ɳzK��O�"�Z��5���.=w��.,���Q�1�T��xa(�j��t��:�1�D�&_d���w�{�G����~1i1�'��D^ou'�QU�>�D �~�K�vL�)�.����ߍA����ց��q�� �&hL�z��r��]����e��g���TЉ��=���7�������m�[b�4sS8��PN�0�=�$�g�:��o�I=$�Z� Ŧ,u.D��M�6B�1Sv�A�����)3�x�	�����Sᖠ�7?�]�d�s��}P��DSXl=�?�v��.�5�e�D�z�1t ��a�`kЯ� U��0�}eO�2��$���n��%V,�}�)ZAҥ�����búk�A] �,�"L��P-�{�|���$AS�AЗ���-O_�r?j�ݿ�&�Q�]B�	���5@q'�xջ�kX���C�x,��"D
�͞p���6��?���b=��G���,+N"ie������;Ȗb��Q��xKnQ���0{�-t	��޺�����y������w�Z�m�h�b�i�;nW'�&JS�aMb�S�؛�{
�u�gN�?�#�m��w��}f4��9JS�K���+�V����dށ��͖E�d�J���hӈ������@�Ktз�&���(�{q�޸�Gz�Yz/d�6V��t�{�V&�h�53f3�O�%��|bC��.<�1G|O�~E�xȾ�� آ��z��[5Z�B+���z����d��Z/���b��x�|]�u�����YwC�(p���ZA����x���Ѐ��I��՚b�8�Q`�22���Rs��!�6���$�]��U�%{I�w�7#�r����b�2�5�h/v�h��S��E/�K�S��_z��6}�3�T�c����
>� .�d��wU��[wr��6SA>Ha.��~�U�&���ن>��6��M����g�(u`-��v�a���|��2�r�������ـ[��&�44r�荇$��:ds�rG�]�*�>Sa��Ƙ�uS�8�EE͈�,n̋�Y�8T���j³%9�٬��_�6Б8�D6P?�x�� ��<XH9[7���g��G?0֑�ْ.]a���.6���FI~��!����k]�h���11M:��kgd7�cz���k��a�ݓ�� ɼ{G���j_��x4��8�=yf�����t��c9����>+�73b�!�N,]M��G�a�ggz�8�ؠ�宀d�&�_e��֓~�9�Z��Q�C�4��!B�Z$�� g��5+;t�ϣAe���?����:蟭OS�(B^�γ��'��i�I�0�q�!V]��mi��M�����}7/�d�����p}�<=��n7����]r�
�4�P����cK��l�Q*h���"�Z5��`�twQGVz��#=]��&��}&�����L�p����v	8?��N#{S+�$o�d�N7ѣ��y����[�Ԏ�7��v��n�e���nS��z�)pM�s�S�T�= ������s8��X0:�a��=�$<pp؆rOVc�Ph$H��8�@�lQ�Sa�WiP� 1��Y5u�$���p�ψ����u�(���2�$#,;s��@�u;Ԧ�Ka�%@��n���DE�@��A(Bhx�Z�pdk8�Ef�-*��Q�9 ҂�Hn.5A
P�+ȓ�ֽ�jr!FZc�"�'�:�'��BȈ��8��|�-?��o	ݯ�j��/��|��&�ܥ��c�Mrf��-C��Pt������˫���G/
kf�@�W��g�@�E�35�)}�Me��}��B���K��)����j75s"Ct�g�L����_�3oH�,��:rm8�M�"�{/<�qje���l�F��	Br7��V꽥�������T�*d�����E�+�e��ϫ���rWA�Q(�|\ء�.[���$κ�4J��FP�����y�.�Ԗ��L|�4F���,Y3�ġ����! ��xA|�ex=򄙜{���/k]Sc;-�h�i!��W�u���o�שwwW������+[�l/�d�Fr����H���i�
��?Q��/��fD�g��:KL�2��qYE;(���2����߶C9Z��F�ӿ����<Q� ��a���Xl������Z�O�oOE��/���\	�N�	9O3¤�[��.��-�شq�8p������y^_qn{���$�߮2�����Þ<~��=!��&)�c\��iM�R������x�+�lx��,B���E�&�{������j�$7�9̜.��=�m
ΏcҊާ��W�K�Hꍞ/����rr������Z <��B�����[�w�@	JF=Q[`��Ґ���V��.@8�\����"l�L����MM�K���ַYdh�90��fe�3e�iנ���i������L=c%�=P�o�@Ok��#���Y��\+�O�N�#Xj%��T+e�7�/�&S��|8ddօ�x�gq�wz��`/0���䉩��0Xf�Z<9 �l�y��a���-�UQ�&�;�\_��W�`�S��-����w�P���p@���g�K��Y�h�����YBL��~�:�q�0�|ǎ�9p3���%�������_ђAK1L<'�m~Nj6���+�7vM:��P!̲']����^0�՗�H�<ai�L��,y�����r1f�����u��Ҧ6�b�P��cGk��6�[�S���((Iw����2�~�]tTدc��=�_B��0-(���v�H"}����e�I@mӘ��i���R��� �t�y �C+�+NP4U%�5�t��IF����q�6��_g�{��qy������ç�J/���^��@��M`�a<G#� �騥kptB�"'GT����j��/��pі�'�pYuY�!���	4�� !�ɥ�e0���ߺ�mѪ������e�b0�I4�^jy2>%㘟����]w���{��}藋���b���_ym,�$ѩ?
�f:'�E�Sh�3��Nǁ�� Yz��To�6A�,v���P�S��*v�Ds7�w-){3,X�Ջ�����3��;���{ʣ)nl����;�q��X*d<�$�Ƽۗ<��r,(2�v��T� eb}VqB2=�4?�Dw�z_xൌm��f��vb�����1�u��&�bd��gq>h���e�D�r(Q��&=�	/CI�$Er�yM}�bl�Cl�л¦�(�<ygF;6@�a�+��ʤAf[>�>25C%�p�(wh�,?����<���LT�������R`�lv�,�� ��TJ�Z�gi�r��
RC�R����:Gܵ��U^n��L�3gb�KH
�_R{�Cj���$��gu\�{��iB�r|/A�#W���_w,�-@���y��S����uxj\�l��{��+A\lI���.k$*���9�!!H�3s�^K� ��E�b �$�d�<���0	5���(�`�{n�ʚ�Μ���M�a�8	)yb���ON��޾6�O��M�����e���
����%�C��ʪ�8D�6�]B�6�ZFlU�
�@��t�q�'�	2�zPʮ&[�j�����^Ҁ:��Km�8�̴����k2R���3�>rF��k T��v�~r�.Ω/q.k�?Y�JC�H*�u��H�������<D@��#���}`��y2ƺ��	��d���~	�$�P�5�8��]��ӂ�6�D�2���-%55w
��n���
҇O�.Q��`��^���z��`ꗑx:!4|�ļ[h����]�">�e�8z,�,���I�z1)i����.�:f=�����y�iՇN~���V����L���Qpy��s��F��I�ѯ��5�MÁ
��&Ģ���Vzɟ�.���̚��ؠ��fl�����N��؅o�.��G7UV�_h�p�B�%@����m�c�\{��< �X�`fz"`�1��x�eF��&��h��#�=�[�?��'}.	�-K��Y֯����c��u��X2ukJn����������a��;��S�n���UOC���	R?�p��ؕfy'�n�gr4g��G��2��A��R��XF�|����xxz����B�����oĸ��~�[lh�o�)�;�J��ݐ��������'�*�r��jxa�����i�2ʹߘ3�R3�Q�v�#5��G$���G���C~�����\#F�������k�??�l����*��h����!rb87��2�j߃���*�&6�^pd�����>������eHy}¡���9�־���>��cV}���zQ�-�M�z��$-8k�0�4�>@�5TzH�F@�|��t"z�"\��e`c�>{�
�3�	7. �UX'��ZmG�vV �/����r�d�0�l�DD;���j&wƶÑ.j�����r�=o��>��M>�S7�������{�EXvW�K�L�]�(3?����'�K�=�&I�$�39v&���(����F}Cv%�������Kj~�X0��wU�[n:��:�Y�P
/6yZ��^|���������c�o`��(^�O&�:�ǻwA�7�gz�Ci��%��a�J�P��{!C��W'�f S `�N�I��^?A�R8��7�C�-�ѻF�#�N��o��-��e{�A�-���}PO�;"oA�Z���e,߰J�а�u�3� {O���U���+�SvZ�D����P�κ1_��l�PB�W�-�ɅG���H���Vv�`�<	�,���o�kf_����31*s��Ӕ�HFʎ�VO�2mWj8_�G�c� v�HQ�K����Y��}9����bH����2�[ANpru����&��6��)�!,w�6)��N��M��]f0�o��s����V����Mjv��s����행�W$1H�� q���Օqկ��҇���MyµW�B�y�(��o0�{1��;�!^hz�f��4�k�����}�lJ����	�n7'it?��Hpjj�}�� VUqJjFG�qD��j/@n�L�4Z�w�7�Rw���u3�g��s�V�@}1���f��ojܓ5؟B,!���|�e���)�W�?~BL��ǈ��y���A��v�e_��GZ�	�!$%��z���<�5�s?{�G��KSS����e� .�q��@?D�h(!���_�7�d-\-��5�+Aat�8�¿6V����	�ϣ���@T��i7�q�LtG�$JV�*��rỖ���'���Rtn�(��x(����ǭ�"�͢�Ѧ�b�+�n�b��n�}aF�D���;6N]
R���cnl@���I����@ta{S2vwǗv���_���$%�����AUW��!	|��9��N.'	����"Wt��v���U�)����9#Q��@�Gu��"�%�s�eO{c��_s�)ӊl���$��R�do��h��Y/���y^���Q�Cr0�\�:u��Z��y<a�#%�(^T��dKcS�Ql^\��{�K�tv�kv�|a�.<n������z7Km 1ݜ+�ՊD��U��"K|��E�AV����5��-���5�0kr��"�v����ۘ����?��^xj����6�}���1q����x�|�!�O�� Ub�ȸ��!/	*x�.����_P�&��dq鱼� C���4�\��y�f��I���G��i�዁���D����D��%ꀼ�_S:{����`.O�u�0HvC���C�E_'He	)2�bZo��9�r�Եk9�w=�n�ϴ!w8��c�g��1,5Q洤�N]"\���+�M�Nƥ�tǷ
<щq��bJ��|:K1�3�2��>O�'¸R����E=�`7�{��-�Z��jq(��A6;H�T�p.�Ǥ���g�kd|���jI-n���H#՗'��Qy+�np�,{L9��S}f,�oG5�WՍbrV����y�n�e �3��=5ь�}��zC_u]�nxn�O6PD֖��s���p�g�@�b��"C��v_����3�C�\��ԃ�����ҏ��3������L�b���ymM�|�i�>~
�=��8�����,�M鈡=N9�I���'lu�&�f~N�ɀ�ڡ��a�F�w�ݟS3V�5�6�������{J��mX�	��	h���5m��Ojg^W�-<a���dq'�!�O9�/RH�t�.���O�m	�#���,�f�����B�W�	4�ds k��ؖy��`k���Ό���.&^�y}�r��������xw�xN��y���L�Sj�B�6<��H��2N�NG��P� Vm�
�o��\,
=�����\jo�������!�Yt�\��ſx��{�3X���mNe5��(L�����e�f[Z���S`Eꤔ!�U�vI���N�\}�
�����˥�OB��!����j.��ܺp-���n[)���:����vXn(�d���@�TA�O=x2���������-�H������"�`$����s®7AI�!����`H_����9�ņ�:�&B���Qx�e n^��.�%i���SݍCkg#S|��dwL*+m��<d���R(hXA45��h�	/��J�^�}�E����f�����Q�jB��#T��	A/ق�{Z9��(�7�O.�F#B� �F�{L)p�4[��G��*��s��%�RB����V�G�i�a�LӼs����i��(�}	���{q�ʦ��s=t^w4-_D�T|�
��Q���F��I�؆1�@Z��O�� G���Os87vgMRG�n�)�2��J��P;-kL�	0��(��vZM#�H�$�����!Mt��izJ��$Љ]�.+�<)�Y���Mw�v_�����T�ԫ؝:�o4�����_����� u��}�����O����;�N�C��\���S�1�!���ܨe��qP����_鯍;n�U�N���%=��X~��2n�rR�{*�Y��=#�k�ɬ�,sU��E�)6q�u[�\s(��R$�|FO�6
�%��m?�Z�^ԫ^��a ��M"� F"��szF���B�-��{ ���?��.�3������(�˭�F��=O�W	�L����ވ:�9��2�(W�{���m/P�A�VRy���Mm�ح���)�Jjw���@ ���$�B]�+��R����N������Q���7�R��{�Oa����C�g�0��)�k���p&��R�ON��Ԛ~<�z���uq0Z{��	t
�+>���7�{Un����`�O���Sy6�l��������w�T��j��S�J�`s��b�`{��Vk	����Tь�@C1q8��w�c�W-�fo�K OP�$+��7�� �;\�����ӻ�Ml�4J��(:��McĬMy���|:e��ưcz���e�3�kLr	&h
��JN{Y��!�'3D`�4�|X�$}܌����_lU$ͨ�����P��8ݕ1r�0탒2���6��7QAm2�����	�-t>CU��[Œ��FR6%f�ɢ�I�W(={���-(y��lo���D�����(רF0���"��z_��!|o�׊;k��þ�<;"���e��\"/�cVyck(���=��k���F13�����w՞g�j]��d,f]�'_
0���}�����{.�|���x�0B*�^��~.rő��э�;�AZ�ot�W��,�W��쩨���H��_0v�#����6aD?7�m>�i}=�k�x��8��NJ�U�5��~+�X�M}_����%��S��D�i����@%��c?�d��t_���A�3b&7Fu�"_v9[�|q�`ocU���l���4�C�7���R��ȌS	�F9ǹ����������K�x��՘"A�z@�\|K.�#��� �=��Q�s1%B�殟���=I�2�{[�^?v�tj�iR�-R��΀H�W�R��q��A1uގ������k�*]����� z@n* d�c��"�˻4�a��;�o@k�83�D�a4��ADh���e#�˸P�n�އu��94j��0J%���Y�KzVݻ�6z�V�����������A|��r� �R���
�_� ��k�)�v�tidޘ-��4T�,�ž���)�3,��Nf��,�
ZD�s2�����Y�*��6��� ��V�0-T�d�Z�8"���W��[]|�F�ҽ����&�B	�����?$����V�n�\*'g�QL��.Sۚ+y�v��3���^
�S�U �脙¿�v��OUKfw��x����щ�G8���\2G�s�t���f�� �QA�/���K=�o��"[�k�� ��}Vr#�����*�[�m�7Au1&"��t��»��N���Qx�9>�E���K������E��Z����_�W�B�
��ϕ5��bR%�e��]�H�$گcrodA�d_6u���'f`�l�tÕ���R.R�拡Bkp���}Ҷ��X�
?�@����r�}�d���3�k�ڤ�gE7�h�gv��͚s�E�޿�e�����!	��W���*��k)��^(`��q�HK���xM��3z��gʼ٫$]m��GO�p�-���>�+�#����]H�z0}<`l�C�޽֛u�"�E<��/V�M|`D��8�rN:�0�>XS�+���Y�QL��a��6`���X���D9�3�(*-�"����D� ��� �Ij&(�a��L.J�̩�"xS돹 _���h�޳Ba�|��Ї�݂���	@�d鬄b<��ĕ�-�������*/�{��͸�4~�9g�yl9w�5D���$�0�֠�[2�<1L�ۋ���AS��Q�x��b��G�l?PJ��]~Y��}ɝ��9�mƯ�ѕ��sȝx�����]��x���!2�#��Kx�r�sg���6s�m2�\��|[�΃=y���"��e���{NTZ=]����f��J;��u�)Y~�z�����!����3dPQ�|=�˨Z9wу�����R�[���x�a*9;x4qX���I�2�z��q~�A�ZE�ppWkp���9W��o@��p�y��y �@� � �<���Q7׾��VM�$ޘ�"�;�O�*���H���}ݟ�x�g�H��R\O�
(����B?5�y��f��%���b�S�7@�[8�g\x�	�x����䎏�3*��j+k0.q��o�Z
��tEU��H��m�a#�����C���.�(�Ap�Cf;�QJ3�԰��1�Xz�B�`I��o�^/�,�_�K��-�"��}߇�e
!\������Dy\�g�ę<�:��L	h�F������D�����]������!<��3��EJ�&�^U��s��o5�[�e���+o��P�I��2]-x��eJ��J�U����.�?�*�W��ҁ�N(�������h�;p[/@�K��j�7u�y��	N�j���f|FA�o�NqGgQ��nZ����fBl��G�?��@L�/s)�!����(�kl�t��UWO�R,2n,��GmY���Ǖo�0,^�^X���֣�q&)"�(r^2�c�1��'�ׯHI"�Sh�%�0�oc/E��������d��/w�=8���kRu#W[���������8���8���산�9ޏ���v=֖�f�=T�4���N��S��tj��寐V�<��D4�l�UR���-��g�kP��#��Z����~k��#ēU�L�4�8�/G�8}�Nh���](\G(����KOQ�|�P�R
Wżv�����0$��,������m�:��:uh����d$���?���f�An��EE@P�i!�b}�.�z�!�u ��V���Ғ� y�GM�%Za/2Dc����(�ha��3��yv@t�� ��aC3�j��}V�ǣ���#���Yl)��y0V��b2��O<�V��$,�և橑��z_�.�٘u��eN�f���M�L��3���^��� ��#-�KO��\^�;Z����ޘd����^�a����i���z���9ag�۶ Y����j�#��D�m��<�dI��t�?H�-��{��x#����<��)N҈��nn ����αI�P�M��>'�7�c��O/�0,�k��A��U$u4��U�4̟�&i�o=�5���^6�*�R���r--�K1rчC���vg�͇�V�dg�d���E*�*��?}m7� %��P�������B��d<�a�DW�33����N��K����J�,>�q��_���Ǎʈ7�v�ަT%�ޑ�.3w���OJ��'�av��-�Pݤi���x��:�߳3�ܭ�-\��2��}X�=���������p=��O�L���˄�����<[�V��#M�Y��|�k| �k/E�Ѓ]9��9�7��i�y_0���)fZ�g`Ow���dG�XH���VJ6�]�}K_���r�J�L>�Ŝ$�������p�U���#�����?|�-�i2�]���HY��)�|�WB�:�.g�j!�Vs�����3fF|Mvo,IH��BV��
P}z}�r8�Ū2�N��͊Uf��x`����6��v���4�H�z�Ů`��R!�����(Y1܉iѦH���,)��	��N>U�_Ƥ�3Y8�?�|G�D�F��k�;5�L=� ����9.�ܣ�s��Gy�����S��8Q�۠}��E�{��vm��w�<c>��-M���\A`�������~Ql�J��c�3��O(�-z���}�^Nxf�l���E���,8ɔ��e(>�a&�ZyLZ.���Ƿ*�s�0�����*�<炭'���m~^�ز�Mb��D�˛��BU�$^�ZN#���vc7��n��l@�>�"�Bv�)��u��� ���2�L ���G� '+Z'Z�7�� J W�Px)��*�)2S�X`���]j�p`i���k��#Ղ5��?�͑���v�c5bc���WhA�&�&H߳���3�H�<�ƗѾ�%ڃO{�/���9.��)��S�Ѓ����]Ĵ�~��� ��0uľ#�J>��9v�y:Dd�'Gw�?d-,Y���9���6���=�ـT��$9�d]�8�5��A��/p��4�(T�(�J���֐Ҩi*������hS
����-�~���0-7|3om��H���_�H���6|������+2�4e��#d��9\��'���H�:�r��O�-���/:Ӌb��X�+�ؐz�̵x*"��C��^�0��VT�vl�����qq�Qµ�Kdg���`*�/��x��k��.۽ u�c���|sآ�י�G����4�4j��%]��/��M��e�n�F�q
�� X<�DN�1U%��j�(������d�wu���Z��m
濍Mh���B�ܟK8�j2d�,��ɴb�Dj��L�q�0�o�뼴F��>E�#`�j�����5~�Ⱥ\���9�(�ݮy1��>�t,�p��DB�ћ��$-���P�b�~���=���\��>�����C�D�x؍�
�ɷ��I�_�wB$*���� ��ۣeD�CB�wB�̲E�m�XQ��Nv�����Sc �K*�ۈ��Ҋ���"�6%�I#�'�^�=\3b��Z��g��?�P�ۜ�}�A}�f���A( cgY�����p��#;JqsA ��w��
�b��d�R���z~�Fۋ�<���O$�ch��h���7z�ɬئc�l���̔!�&T1���!O���~�f¯(��%_�DK������e�%�E�5���T`$ �)���������jR���/��XEYW��9���0�x`�g})�? },m��j����S�V-��rL,��>8d"�F�P�4镔~�Ki��"��P�1�����YN8��xЛ6�3z�bY[I��.�JQ�k��\}%�9ߤ)�,�)��0�vkm"�m��&�Z�|�nr2�Ԧ��Rᄏg׹�2�5uxHp���%��$���#���V��W��T�`X}��B�֋����G��JGm��_�m%8)���h�J��$�W6�Q��v1����5����/�7{���HY�zC0�qI
/m����$6ZV���n��Yw��Ӡ����c��mzӞR%�o g��;��3*3�H�a"�D�#� �,��BZcA\/�� �I�O,��f�>��m\�?HH�ϗ�)T��4Z��E�U!�5�8���t�σ#��]��}�+؟�T��ڹ�=��p�;�)�ZjM�s�G�SDB.��ݎ��Xய	��� �N��E{1��3��Q7A�2�d��q�-AAê^�����(,���vV��܋�ZeFQ�.sO�6Je[��dڭ�X�²Ĺ-`���yu /�����(��Q�Y3���!\1Js����4�Ǯ���f��=���dL�o�Tt�&��1H�����p�UT��]UUn	/��B_b��
�����q��z�N��N�'��px
!ώx����aS�#� CY��/��W�v�$1�?�,�[�㯰P�k2�u��Al/p�z���Dp���n�XQ78�C��c��mgv�Cl=�����R��������>�[3�`��s_xa۳W�7{(9{
��	h�����GR'�R��E,�Fl�?��%�vw�mT�4@"P�?Tt(�I�|�5&�6_0	��C�ZÒ��}�5�폳���8w@�x�ѱ#��������- m�a�_�Zh��,�+hL�Pf��c�M�gj�p�%$�"�<P��U�7�}
+�Σ���W-آ �\&����V�Q&ed�ȟ>3�sw����T���]�|K�շ
�Cނ���c��AH��������k!N['�?W��ݸŜU�|���g���(�XC�, H&,GZ���7�u��6�]�7( �B��ͅ�)����%N�n7�&�V_��+�1v���<A3~/��;�F��hB !�:����@:�RU�iz���i,bcho R�Q��������E��-G�����V6�I�-�#|Ta©+���6�n��3�'kU���{�y܇~�1�٨i��0�?�3��a�ۦ���t��g���%��p|�K�%f���C�����0*70P,Ϙ����~h��5�S���5�+w{����hҴQ��ъ�?�Ł�����zP��d�QI�L!(,�0i�s�tYm�,,��.)�q5�`A.���K�"�0�O��9Bh<����be���H����T��6,Ʉ�{�kޞ����	�p��d�;��׈�>��r( �,^���~�l{ѾV�2�C�쭵�`mh�K���x�)��W81�p��v: 	>���Rex�٦!���%��� '�(n�8��\�X+��W����}�
��X	^zFt8lr�rf}U�hN��^���<|UJ+���U������w�2<(t���Mu��\�% �A��٠���+gĶ)�7bfӐl�5,�p9Y����a솠��xV�J��K��06�s��0e�yq�n��K��gj�z�3�>���������#d;1BsZ�5���	�7� �2�d_�����5D��Og*�95� �s�>z��0ta��r��.�ی*
�:RN1=.�PuV�^շZ7[@�9�mZ�/���SH��(ydI�-Ez���j�8\#�V�I�Ka"w����2BUz�%����GPڬ��Ɓ��c�$J�,Uc�k��?i7({��f��k������άh<Ҍ��[9���Sz?��ar�0�����K�.��^�3	��=����?��+��bO����G���#� ���Lδ\���C��<n�a��O.M�^�]�e�m�,1�{�}1���%�M��A��oE��K͊0Ԅ��[`3a�V��P��"�G�*����WɃo�U-�cΤD#\�uz��$]�~�^�5�R^�}l
�l��l�Y�<�N:�h�j �C}��vu�P/�y��O6MG�h�)�]}��tQ��5�p���O�L��h���� ��f�^�\�ȳk&d~Ԧ�Wu.�!��Z]R�-��Բ���!�v)gF.rz|/��. $}��W�U���ԁF�q~�0�A�B�j��Cx��^ɾ�J�S��
�_������*B�k�AVH�:���+Z�j"��z�!f���-D�`��Et�iJ0<���5i{��L�gW����m�y+18˝�z��o�ЗT�� ��{�"����ۈ`n���XcłU�f%�����ؐM!�!���������B�q�/��yO��鼟��=��l�H�Os���F#��&�v�Nqǿ��� �g=�Z��a�1'5�/#t^�<�x��ef��Onְylghp��ۓpoPaq~ދ���Ȭf���x��M���Ckm��O4E�X�gj�c�.�;�.�X�0y+rY�gGfn����M�7�[�ʃ0R��z`zd�:��|~�5�2��
��߿5����7������.�N�ePj�G���A����Te[o�3���ٚ~m�c�u-iC��h��?Ԍ����"m�O�%�>a(Nq�.;Ij�2ۣ��]�ݱ���-0�E��+�� �!z��yö"���`Ɋ
٦���غVv���#r%���i���و���$=�kc�`:u�o��R5ݟ^L������Z74�3��
�b�g��"O�pP��̉[�+�����ryA��@Sq�\�lcd�;`��D�<�h:���]٨����ۄ>���!��{��X҉�SЈ"WD	��VwC/��@x˭�4����T���>R�FB� ��Y�V�4X�%U{5c/SԄ/���s,C��@�K��=����2�62�q�������ƾŝ���I�
5vy�j*��h��L��ӦS8R�j��l��Mb=��|d#c$&)���2�,^i��M��\�KM��Li}s��\y�1@e+��E�׬�4�xNX�,R4�F��s=�D���}ֲ\/!��W�c�RВ_��w!KFY�s^��=�X^yW���M4��uTo0�de�;������t �bR0똄��z��� o~���3��Ӄ���8
��"9?��b<q0t�BGW����u�W*�FO�Lhn��k!Xj���=����ڛ�c�c�1���1�mwp�����E�y��Q\��\JW�Fb��8}.�ۡ����l<��연�@�e �b�	��E��%YU����%�K��s���)W�L#L��eC�z����H��d��evz!�?�k�j	{ض�f-�aFI�D43ē�T��"������ձ�J���7�����f�2>��Ed�](�@y��]�����S����e�ZPp[H�D�H�_L��tR�i ��;�[(�Ѕ��Y�E������� ���R���Tj�[_uJ����Nhhm� ރ__����SO���'��Y�5��ѕ�������3��h[�3HÃ^�C���7�9�S,�'�����a(�+p�<2�9���؋�i�=m<���/tTn��+G+#2S9P��]�c ��GtҀO���&�ދ�ȆkQuy��0�:�!)0��� �v76ɓ�)q� ���?#".��۵9�7<�P�w�8δ$��Ľ��{�EVٍ��Jm�7�֤��(Ct���B�U�&��5TP��� Ǘ�o�v�#�d�`Z�A��8������Ȍ
�52����i��S��$/��;��8�HwDGF����V`M+�r�-���#�^-�2��Mh��i��!q?� XnM۰f_��[��T�cP���D����jp�6������?����q�8�IF�ؗ���OI2ATz�e��C��6��
.cP�z��<��-q�y]QuU�*�� l{K��Q�=���=��ĳ���/�Nr:��J���U�f��!�Hؗ�8z�e[��#aF۾0���!F�p��o�3�B��ӽ�v=���vp7�%�F0���_��U0m��؇/�����I/�T%l�#���S2����<����w`+���%��Nj0^5�$$�:�d��1.��82(訝�e�Wb���F[] �e�?���`vh�#�]R��P�]�w���yE���V���IB 6��XJ|��t�
�\��5��6������v�N� �o(��L�^���+3<n�+�O��G�Ȫ,�ݝHY�)�����K�o�s{�d�(�a�P,�`-J�GĀr;��'j��vw^/������Z����"q3������*�x%>ڔ/��b|������D�"W����?:��
�J8ٌ>���P��F�Az��l��d�Cn��nt�5Y��IP5m���B��7����!�A��򧍣�����Uk	�1^���c5�K3ͼؘ�a����e�sW� L�J����'bBYE��T���}�
EJd�lD�h�7�H�H*��]@/n�&�~���� L?Vz�	~=�g�@��v�B��X)�&f��UѥG�r�5��2&)��#jA>�17�����[.��.,B�(��}�`6��2�ʑ�smop�,��+��h}WQ*f��$���ڑj
��:V���d�RI,�(�K�ҊQ���-�J���|gCbmf�ys�!H�_^z�6S�����K���>g����q�j�}C	s$b���XJȔ�{)ԉ���֋lv�q�ig���W � wVYğ]wg���T����l��֋��Յg+��V8,4w�l��\��/�XA �Sh�V�EM�+?�� �#O�)����|ux�x��^5�1�@�v�d�)�� B�~��YN���c��E�T#!���<�]�X�''���x��X���*�x�\W������E�r3 �e���j�ys�"�c����ɰ�6�����7]�R�)�4��e2�������rۂ�*N�~N1۫��-�����UU,a�����P�]@k:�N;����+.*0$x���"ؤ) gG�<�fHP�m�h��;����k+��`]rОMఴa�����(�:#�>�����mr`� 3���HF� �u�H�y9��}��(�Zn�#sZ����
ڦ�z��h����X�%s��
�H�l���' g+�g���o�� �<i>c��ƹ_P?I��QV�gd�G�7�T\z��Hm]�T���@�W���n�U��;Zku�ב`Pj�N�l�͔���O�@�d���d��5����mr���l�sQ�z~HW��wͩ�����S�0��ӝ�g܄5�˗�Q�j#k��������[��#���8y��B3��Ep���r��6f�Ƅl��`�լ:x��Ie��}���E�,o�]-����O���8֑6�\>���x_��?�v�������XV�"%�?_��y� O4�Pe��uYh�[6p`�Н*�3꼭R-��h��2�U\6���n������p��8��4��3$Q"����n��*!���PjS2cta��kI�˹P�I���t�~��ڼsܛ���X5�}�;m�[oA�h;F<���E���{N�Ll�k$mz{��m^c������W���ΰ���4��5 ���1����!Q<�w]����I>�6�����zI4�H��
����<�d���N����)�(k�o�+�7-�����K;���@������$��Sf(' nJ����NG(H��r�;�F=1�`T
�**������#L������B�4�Y*�S��ĺ����^��F���v���}�wfc� ��^2��=� G�Y��w4шQ�߻�g[O���!���E!�:X^sVH��t'ۛ�3~r�n�e�2�(`����/�O��Xj�o�����h�c�/�t#��y]}9d-��%�&�*��Y
��dS��UF��"M�5�^se����V�&~G���n�)�)�S��T�x1�ҥě�PO��m/EK��8q���r���.���v����#z�<AtP�I�ܚ�H��u�� ���9��xMR2�͵�&kR�!�N�Ǧk12�� ���8�R<� m��f�p�����z�DWCn���