��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ���!�T0O�'b�O��μR��MJ���q<�[�ń��,��ݷ�8�=�Щ�u�iuж^Uu�~n�w�� �biD��4�y�G�z<�%�9jT���m;\��P�?��;�������t���Pݩ6鞐]A�S0Z��M�i���'}�*ʴ�K��8���ʱ�L��P���g�D6����Ehsc|�G��2g`Hڄd����#�)��ݓ�Q�����.Y�W�Ĝ~A��C`�K��έ0�Qm��<jhf�C�����G���D|_�����C�S�%r�~.��HDNiI)�D�>�͇~G���Y3'�(~ Z�����w��ǌ���8f��m`k_!c����b�*�� [���_x� ���u���#�G@�Ҁ�Y�Y�(
GwK��	��,4�;>W�Mn��V�Ĉ1z`�����u�������5dͮ:�0�������5�+��p�U��D����'�ƻFb}MRҧ&��!�N�zɃ�͞>p�u&���a�n4�o�l;Q;0������[��PE�����4�N�1��PoP~:����{�΍�¨ٕ����+�Q�r�L����m���j�SȜz�!�����7��Rr�[����,����z���J�uc*TG�L�6�B��=�ͽL)����l
�X�p�Q�S��X�p�AŎ�n6�/�1���Yڸ��yѪ1�nVƝ��'D�� o���z�����|[ښP͟r�96�R�G1{Ly�pt;�n[Ձ�V�s��J�z�e9�����>'N^�O���!w��.�N{P�%q���6��@�[-�h1���	ya�`��	l�ܷHYv���#��9p�����dY����﫚07�^����Ì�/w|�aZ_ i�W�?I�4)�r6��'=�܇����_���Nb��x����S��9��u*�v��o�����J/�徠d�1yn�CpO>�Z���E䖯_v����v���u��m����hʟ�M\��������q��AӰ���������h�q���gBN U�I���"�xB��L�$V��5��P�9c�$��.5�������	
 K=zI �=ɕe⧟!�~O�B�qA2��C���+����r�-S�0�+�}K� D�Ro����Cn��ă٥��Z�vJ�ȓ��^N3�%�}��������Ĳ�J�7��87�8��%��z�x��W��4?zH�C�p�I���'}ՉO)7�Tl.��-�90}�U;C���ꬹ���W�-�.hD�B���^�>S~m]\[>�3�8�
�t9A���#nT���) (n�R֯�Nv+�Еp&j�y�������fc��U]>.�T�oUj�ϓ##jTR��>j
��@\9��m
�/�}~�Z;�C���u�LǳXc���aiǟ|pjx�������D�Ѻ��qâX�\<����b��(�B�m�UM�Q�&���_b��O���J��&`N�"g`QL�r�G�|-l{֪Z2uu����5�7<���N�Ѯ��̯/1{�]�֋g��r'p*�8Dg[d�	�z����I�1��r.<�CN����D9ѰI�˳IDR����#<��7e*���̉�9������ϴ^|ڑ��� ���do��%��h$1���l��	}@�����Z����]u	��8��c�n=����tE|48"dݻR�*��)��چ`�m���=���(,�k˙e5%��%��7��=�~�ʇ&�������Bp���D\;,��t1�{Ar�/�_����(��E@��F_
`j��9f[!����y����{n7�o��6!)��|M��>�
X���S��)s�)�j������L�F9sT�_�F���/��Zu|d��jE�1T�dRl��dv����f�l�x�D\_LqE@%�.E�sT�=�L�����"~�n�DS] -q*]O8��T� R�m�eD��]M5��ؘ�$�w�F����yf7x�����޻��|�L���գ9��I.Q��h�N�+�5YU�N�!ݍ�$6q҈���G���j�)�tޖ�� �ӂ�4�N���\s�;JА�&SG,�?	�F�1�G#����XR[���{��oq�6�6W��C��Ewլ8y!�"V�P78�#��j �����6�;C�������B%M� �:�3`�V-�W���u�N��c��ٛ+ؘ"�ȕEs�*�r�ƊS��J#�
3��A(.٩����7�w����m�]���i3_iAo[97Q�w�����T��k�S�V4�?D���i8�v��ƴ��\�_O��o�4���{
-�?6GOq�j�!D�`z�)��q��7̎�Ə�׾_��Q0����N:Ȅ�n��`j��L�;��4�m�"H0��\�n������ l�+I�m��vC�[
Ew�S�ZuF�]�`�'r'����3[(���h(��
˥�����+��u�3KWt�j��pV�����gp�]��=�g��i���`��}��G����uB��C2�La&�~��>[J�1�o��G�ZS����7ߴ/ֿ>�sR�͸HJ�D� X/���"q���R�3y毲�Q���eb�P�B�mR{���,�EG%2K�/��b����:%%*cDɺ��H����W�y��b:,��g<�O�S���P�LE��\��Z�g��	?��V�g]�P�[�r7%�!�^�4����GD��2������)�t�`����a��;��U�;ѱ�~��՝r˛��_�h�������cf[18͹[.V���ʓ[/:���#�`d�^T�9�[�5�q��ѩ�!��}�%�j�ȁ7:��rE0�)�uD�=i�殘�x���h��D3����
�%�x�V����3���Y�5'p�b$-�� �=6�m2нNa�g����n��(�c�=!SJ 1���(S�������O:,��x���%��LM�_����P)���~�2vnKZ3�
9ء@M��|,��8�S�d�n�ک��w-	���(�1�#�?I7���a 0����[�B4+g��M$E��J]!�PG���@�"�N&��pS�������>`}��I�{\ּ��-���;ɋ�߽��גL�gK�,�w�]�T�	�}�P]�F�%(u��=ح��V[$��y��`PT���)rZ�S�?vMJT�̀�M07
e����I�k�Ƣ��*,���[W�
ϗ�i�u��C��k�A��w���H�	%�U�炶Į��L�5R�������A��#�.�/��"mq$�q�G~��������0$���!��t���E1�+L!c��D��q�ea32�v��FdX2"�BJR���=ȘӢ���V�U�ޚ�v҆A*� Lg���]��+�/ԋ]e�\�߅���tP�PQ^�U̸���Pq�K��D�����������s�"òA�H�e J�)8.�t������bg��Lk�zh��%?�X�qۙ�ra�3[nR`�y�W��~D�u���e�r����2��W?�|>+=�D�D2�L0{�*�i8w%^������h{���K=`���H������@
ul��L͕&s`?�	�7�-(ҿ~�r�o���2[=u��D2*�7G����6��y<���f�T3��*�ə�a_��>-�i���	ND�DP(Z����>h���
����Q�����ZF��e>{Կ�K��7�9���j)�Z�K@�� `��ԩI��z�;��P�5#�h�������z��j���w��f�^D�;o��zp�ԜXq3�C���z��8W�i�W��`F[]�����������bp;�;��V[qLfj��c)7���Pg��U�m��|w@��K$F��
a�����7D�P�&�B�E�F�-�}ǵq��a��N2TA�P�@���2�E����s�I!2M���v���疺�J�hΒ$.R��a�	��spf�]~z�u\�ҕ�s1�!�Vp�C� I���f;}�v���w߼���Y���2��}������cVhg�_S�f�D�=�ϿB�;o�g����M-��f,�)pp(��O-,!���#� ��p�o~⸿Z����}hX��Y�R֌w�֞n�O.7�� }DjQ؍�D�2�y�]�kD�;��f��'��JS��%����h���F��ph���F���K�ڡ�vp��������Z�:Jޒx6]�T����=O+�1͉d��f���5s�Zb|%G��7[�">%�;���BT۵�`W]e���T�Lv��kBC��E����a.����E�L���T�E�Q��w.>��΀g�I��x�-��#>]�~�ե��wޢ.�)_��ʼ�#��x���~.�h��4��8Jy�ç�������F���,�~� �*@|�ݬ�ǩ>p��4l��DZv�k%L��fm���6w ]ܿ�5-���M�й�I�<�X���G9h����Mm �N��"q�Y �����ELP��yu_nC���XC'Z̂F�2�ѷ^�i�DZf� X�=��FQ61-���!Y���3({�vt$�,�%U��V�1� �xf�jL����Lz���uF"�&6nW��b)�Ԩ	0q���DvLOi�M�a�%C�<���f=F(�-;>:|S5�������5�~e��k���b��qʇCm�C4��A���e@B2c$��!9��3�@�3�S硷�}��S�2j7FA
�^}�Ȩ�k>�~��ݙ䩅�k"�y�/�a1x�Io�pn�8���Ml0���S�bu�"�QIX�z0OAz�}��9����3:�ޱ������� F1�;�.�}C��#O������ۮ�^�3���a1�$a�#ݰH�=��^u�{�Q#�U��X���C�}z�
�t/�i,&���G��h��q���C6�0���[<5��	�T��H`�R�R���o��7�D%ҷ�	g.�:Lt�s�WD0��lv� rޖ����qE�H �aNk��rhR^7i��'�C�ܙ0��tyO��K1�Ε�5+v�_� ��v�CD����ηO3����'}Ǒ�����Pq��lK��J(�C����K�w%p%�b�$1��ll��o�^\��.�9e�Ua���7N=ډ�@��Fp����^��
�(�����������s[��d�Lkչƿ��b*����D����/�MG~%r�P�>%�8��L��MmUc
�����?,�	���S�M!Z�L�'�&����n�Mw���f$1�|�J�+�����ﻝN���|I����Э�X���&Yp`V7���Xg�"��pv���V����u�M��A��GHJ5y�ߔI�"+z$H�XN�9�H)����C�1��lh:ۛ3��iZ8�ʧ�B_I��3Q�����VaY��o����f��*n��4���ǭ�W'�x����xM/���M�j�O;$�C�_��;��/�}Bg���kB5���>��K�K�
cl�fˢ˱�j���3u �to�JQޡ�vA���E�r"�?j��l�ܹ�S�ꏧ$֨�+n1���N�d�iI�.�`��.������F�zֆ 9e�� k�0A��N :�u5_�h������Ĩ�|f���q�U��v֫��2�ߖMv�h����jU)MVQ����D�����^��$�8P�"�b�5Q��1�Q�}���n~˸�vhڕ����H��&å��
�2�l��5@�v�6.���#�E�
^�(f��N���ρز*��ca���m���\������I��~�0��Y3%Lޝ��;z�X����_����8`��3�h;��ruS�,�u����H,��J,Z c�Օ���콠e����4p򗱜7� ԁ8J�E��5U��ϯ`n���R��������9�lU=xP�j��a��\�T����Dw�O_gvʖ�W׊A�t�t��mX��˪�8��E�&̪t�v�g��Y���
�S<ҭ��
�m���������i&�
p��`�q�d���e��G��GߒD�=6��g6,s,�Yw��u����!e�Lijb�26W�	M�t��������GF���(�-��ݖ靑�s����bޥ�
*�j�L��T��>Ԡ���.u־�(G\Km��O͊*N�w�Ȳ �?}1t���j�̢��ژF0���������������_�M�n�D�ԙ�$��f�)����;���ܡ�R��[o���Ѫ@�q��`��wr��d��y��'��r=���}��(d�m�W�6֌��O�[h�L7OV �/�Cp��DO��O�u�0���x�y텹/��yꨲ+^5t�F�Y�۴��ܻ�s��̫-Q�j�\��t4����b�쯄�S�u3�qF	�#��[�����i�PP}���89�__-��UQE7�5��%/9��x	-@�����i���M���`��SǏWq5���POL����O*,��M�[�e�R�r��i�`�x�u�ZHh܀$���A��Qx�����FPE��H��=u[}`�����Y�D�Su�.���r�o��D�N�ri��v#�7��3ZbIn�/?i���?��5V�_R��.�7	��K(�B�n��0N:G� �6�	�BЈ %x\��(�C�z(��4t9)�A}衵P��y�MF\@�c͈S�$��Z����=�IS�������E��۩��R��`5H�Yd�y3tS��E�� �G��:��h��yV ,4Od�K��/�����GŬH����nm�wA��q8ZD���)���s3����¶�Z����zI�8\gh]���>�[��Yq�+_��HnC�E��3�j�A���3�������j]<��Ѣ<�H؋.�i�Ք��"h�j��EO��D�3�ʃz�����i&�z���࣐���Z,G�z֪x��jk��_��Y�!��W4�`f/z�O���LY�2%bN�{i�eJ� �
�)�xQ,���-�5�;`gwn����"#P�Q�叟O�a�;�I'��4&�1M�~�O�:][��*A_)��Kb���-u����y$C(E��l������V�����ڴ�ޝ����K-'�~u�(D���-?Yh�-7/d��Gz��~���h�3��A_�Ķ�B������xġ�Өs��":���k Le`��UCf�����՘���`���g@éƟ:�s����+Y�&'��t7�ER%8��+�u�*f51����M��ћe�~	��)*
��C����Аn�X�I~�j�����ؒuT������<�0\y�f�?�k�i�/���:�i�\�/#OH��5��������+��a��B��ў��j`����wo�ghIs��!_�MI�/ƹ�E�?���H<%���Ɨz�/��ϩ��3T���{����`m|��"u�݇X��+�$ A@w���禍7�hK(����R��t�i"?�k{�D�k�S��F|�����ˁ`����MW���S�w�̩�f��8Ν;.��W��{���ɕ�^ǹ�[^ېi1�;�Y|$����M��ArI����K�̈�O�<��{�u����צ��L�y|� ,��q@J�������t� �Ͽ�W�5�EK�Zx#؃k˚��ܐ�3ſ�#E[S{#<�2��r5���i�#އ�2�ͷ��DE�Q�ەx���2� ������=ziGι�o��5�
>=����d�K;���`�H�Ǒ�*�QBI&�c5��Gu����A�E`7���	hRv���#|�G�ݶ1�����`�a8�|"<3�;ά�����}�qh�B��on9���_��
�%�H����f����O�-���>��^�8���+�8*��eB)�����Q�����m�C��S_��!�E�i�ey������|�N�kg����K��؃W$b�IB��P����'a�)��%��^'��rs�����bs���7��:��ۦ���|4�÷b;)5���&�K3;zGWLѯLX�� ���`��59����h#�jӵ	�JE�������ȦX�ot���d�̃��ŉ_?Wא������֨q��Kӯ���}^����;�ݘ��8�����o9���D'+6��*��]f]��o�u���]�*�Ϧ�;��/�p4���U=A#Ӣ�m~^�`oz�X�+�vZ��UB�#G�-o��&����x�U���I���E+�4�愒B�k��-�,t}���ng��Q�6�JV�C���"t�mO�[�Sr����0������`*��f'��s�f���hx``f��{J�{4�謹�&�g�n�$l�iR%B�ӯ��CJY��f�D5����n;�P�$	�����ZG7V6�ch2���~��u�Kxh��-6�mޤӞ��W��\)C~[�Z�"�HK��Қa/߽�8`]u�	��.�'C2E8[�H�� ����s� �=�p�B[��T�!��4? �#�t=�����r3��O�&«�������2��&a�Ժ�|��Ւ���d|�xc�ڙu��*��D��)~�WD����@�\�#!�S���s�+�>*�K8�R��Bb`�)�!�/�!�ַ6j�-�[*�VL�n�$�Sh����s��vO���0�{��~�Ʌ�Z�/����a��/T�4l*:����խ]6����n�#p3�,dª�Պ���R���ODVW>^
������f>ٻ� R@�D��Ú��ძ��g�m�9��B47���