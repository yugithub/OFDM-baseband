��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�'�+2�H��;KU������hM��>KW�ʊ2�e����|ѧ�^�c}e���bc4R$]�����(�s)��$j�]y�(�y�����G�R�O5@4d��_�N6�lD�{�mdH?v�x\���\N�`x"�ע�)��o�\V����"��i�h�E$\Յj�%�ğ�qE�������G�Yzl_�$.�r7	�9�
��m��,����b��4��I��5gL���H�}�B\n~U W�ҟ�1�i�����&�����2�l�r����uR�l��_nrY�s}z'�C�|v�	��z;+����N4%����b�w�}C$�.�ԟjKf���*��T�K����I*�0v�}�po�N���e�k4Q�PX�D��4��~K?��x{U�=���1$�(B����~/=a��� W��R�����=���a��*3iԹ_)��+�������m\v,�+!���/?���DwB���5�2z�W���659�<Ĥ�AE�0ɭ[Y��O���d�z-K�AT!NT�ѕX�W^֓�kY�e)P<\~%
s�\���͔��x��T�`"ۂ��ms�cq�6����]D�>��L�o�t}���D>�5/\cgoe����@{fEK���%_#�nK�JI<-�%d�d� y��c�k���mq��_�x�%f&�9Y����/�Q�DQ�M/kڹ=5�r�ⵓ�q	��m�C��CȡP��9��.~����7���"�Q1>�>"�#����s��	o��2�>��?�9К#��!�k=��n�]��Գ�$����1��������It+4je9f�������y���u��v�)�0&o7���7�z�1y<��5]7��pc�а�z�J�&��#Z6ͷ@��������G'�M��c��"/p<����Y.�,�I󪹋��
[��@<>⠲���
T� ��	�n�-�b�94��`_�H!dknd���K�_���5kZ�����(�O���@�~B���%� �Fum����w��;���6��R��<!"hwB�W3��x��&�f�ܯK��K�{-g|&B��j�g���0��T�7�x��W	�~����f�Q�ky��X�(Ч���Oϩ�8p�:�����9�
"�G�|�I�rE�~v���aDP~�k�4G����*<�q:Cd*���)8~Z��Wf�ʪ�rK33X��$h��p�r*o��\��W�VE�7ў��M��8M5���kG�?�����Dg҇�G�Bt�j�����+�i�A|4ar�7� ��7�p1B�Ɩh+�iv��\v��>�]x2�����P�T� ���K8,q����`x���K*l��N/k��.��r�}κ��4W��jQ���,?`�Gq�T5Z@F��*M F���3��>z��\�*(���ي�����Kk�r���":��X��l��-�>�3�<Lۿ o�-�1�E@�z8ƀ�'
��[r��7M�t�Ȓa�	���2]ŭLZ���fߜ�Sv�"�.]j�w$��	Gn�EǝS#o<QJ��RR�F]NH�p��S��Xa5-��Cf�f�\D��O�aٖ�|p�|��q�U�����ِ�${	lGH���&�X�j;�Kf=?��L�˒��	O�b� �J`�N$�xm WDS�k��t���۹�-��=]A�SW�:���KQ���q��߮�,wZq+�C��w�-n6]'����������&�G=�9�b���X�p��|��*�+��(Z��v��ѯ7?�D�F��J@��sRr�݅L�����g�����eIɲ?�j[�m�(+��+�,�8ֻ�1�7`�fk;�*���%�[��"MŧZ�|���j�-r!/oDF����'�'A�v[$$�>��f��C�G�q1���'�AH�@�/�З_I#a�6�����F�����&�G���쓟:�|x���M)�wҏH�F�,���"��5���y�/<��Yv�*ѿ	��e�5��]4��U�O�ދ��C��J^{5���v�d�H�o���4���X��ɹ��]�h�7 �{��&'�-�y��;��Qv��bf���/R%���Y**�m�qx���.�k�
}E$��3{��w�@Ψ2hˮ��<Ġ�T��	H_->��%!_�50�ٟ&����ێ8Q
�n@8]��F�����_�e��X�mQ�����J���z���4sѸ�i)��Q�ry�z-�ˏ���{)tt�]te���uwl$��%���_dZ= ��;�C颬�]�^��똬j.�F����YKl�V��.Hq�}��"m�~�iхCp�H1K�aq��zXK8�P	�'�Y���f�G�p�pI~����Z=����j��2�Ӟ�ԑw�s�� >H�O�4�)�}?Q�^~��� %�H+�����B�>���&���a�_�3&��� ,_4XN��{�����	�oD�{��Ase��N�M.1Yrt�D���͆�q�<YzNYS/�~4��?��0�e���n���~rg67����)��^ϼ�E6"T��g��o�E=�zW�Ȓ� ��R=���YQJ{^y�G����/����wlj ��oˡ���5h|����k`]���-%⃅�����<��r��g(�Ak��(2��?K���_�����@�³Ĺ��������TH���ë���0�.��M�r�)���g�!%�q���Y�9؝�6����2Hʁ���}��v�.�]d V��v!��c0�{#�\Ѯ��;��$�I�G\�i�_Y�E��c ���A���(�_�3~z�)
8ӿ�z���9/�r���7<��x��ѧ��}kU���DN�[����ȫ[J@M!�{g���u:�ku�̆��2���{���	%��-�9�s�^錐��S	sY[R�~��!�'�z�/����$M�d��"qu���!$��&��H=���|�˓���@{���'��c�î������
�-wH����i<-��'�do�vݪ,�<���T��j&��XB�ǽ��$&y����ڷ,@��XO	L<_�^ x��O�ub!�Y���p��L����"�&�~I�&��k�HmьA��EUƘg��+�W�bnU(�c���O�3X�D|���L�ߓ�ߕEQj�W4����E�³����V�i�*��8�Ac�E7(q�zAtwi	�;@NN�'r}��i�U'�W�{�߅G/un�G@�R69ak�
c��nDC�R�]I��)�Pc��)�B	�L����N��"ծ��� ֽ�����`3j���z��������S��V\-�
�i����b�$�D�@�gē�Blb�o�K˼�oLNtt����Ēӗ?�sMfE����%W�mJ���;NL�6��h����PY�/��j��#���'�_��J.����4Me�@�m� ,��w:��P�e���M^�,�,�x�!<�/��1K5��sVß���ɇfH�y�7��wQ`>��!K7	�z q?��k#����*�%~���ĩ��D�Mr�Ӎk>�#�� �K�3&��� kR?.I����̠L�im�������l�p��?�|�ת�-e���rc|�Z+b���ф���-�j�k�[�Hw$����qA7VZ}P�C�0\�t���}�׊j5�,u������i%���N�{Pyi�����D?�[_gߖ��
�9b��ا�G�o�"��Z�z!]�	�vI~�2~���:V�J}��d���S���t&��c�HȄ��Ç�n�:\��ݡr�`�5A=�o��Q�����kޝ�Q���LY���D�����m[���0ʼ�͖r6�(I�6��mk= T� �XǠ��a�1�v�B�����[�7�<K��d��k��i��F�M�>��J��t�����|r�:�Є�5ac���:�r��}�q�w�~��r�-Q+����k�V�����y$~�+L0�C:��b�Jl�k>*��re���C�f+�%��>P�[�1����|�V]����1��<�_�I ��)E8f�[�{ǋ��^l�j���El��1����2����>"��ߨ����LC��,tk�aҳ~�f�I?����3���0��d��R���R����.
-4{�� ԃ�S�Eao�/X��1�.���IJ���^���K6������e��|�I�M�"��1�����Y��O�9�����GQ�Dq��	�|����i��̀m֧$�ѧ".}s�SF��F�7�!u�;G���������|,��W"t�4�M3XG��t��^�Y���bg������о���5�(�5���=�O��17�͈!����5TG��_���i�o�I���<�:;�����о��\�&���Zݸx}�i�Z��u'L4#�^�l]s�*� g�`��X�D�@>��`D��4��msw	p+R���^��QūA�c�)��*E
���S_�Τ��<��?��G�ޙ:���Aũ���T�4�/���2^�V�q�I�L����.:6��Bc ���i��z�(�~vx��������ȯ� g�G?�2m��.|2�6칿���Nd�֢myV���Y��D6;a�/�wu�m5��zxS���b��*��>[a����1�H|�SuLG[[�f!5�e�F(�גM��ы���$�
$!�ݐI�6����V����iR/�!?TL�~���x��"�+��K�����ցΰ������-�H�Տ]b��dȳ�*�j� 3�����SlvK�g�:� ��<[���u�w�����riPb��7��ةx��X�k��?-L���MG߹r��S��&����ntt��� ΍�a� �Kݧ��<��KHݍ�~���@�z��eF���3��`_j�S�4�E�F��3��Z�6G��N?�Q&�ܯ@�s�Ӡ�.ɁZY?)��c��u��(���oG��8"l����d����L�B?��Մ|�NyL$��0]p�]AJ:��f��Z�r�"Ğ��{����}�*j3�cN�s�	�"*��l��4��w(��`�R��a=ڨ���~��u\J�8�	�î����B� �'�K8L>� ���K�X�����{G�X*P�Ā*�M�͂ݐ�Dߤ�}1�{ԇ�x�ڄ��������W��E�Y;�o[�X)���X4.u���A�=���g�\#��xR'P�``0	O#[s�	q��ȚH�]ͽ%��dRf�fŪ�Gd;x+�$/<\�i��Cl���,��g�n��5Kh����Pl*$��~�/�f�1}�Ǝ�:�%
�r�O`'��J�@�����߁S�[�3���ՃU����@���3���գ�h��|�$���`��-۩r��ƂgPo�t�ඃ�ԗ����fAPJK�0:��u�^څө�Cm�!��R�,�k�JVI�.�����{X�@�-<���/ӝ%3kB1V���Q&�R\�_�z��.��@���%�6Ūq]��<p�sp��w�:�@����tx����7�U����D�L�]T�x5&o���|/�l�]�k������d��.
2i.oP����M�ߜg\$(t��=�2zPN�݁V0*5�%Z�+]ł�Q�.1|�������3�x���2uj�R���9X�3��٘S�=�.[s���K�Nu���P�tImX�ID�)��cO��&/���3�"t!3Ko|G@P��?`#�����}�Yag�Xa��2{�Or����&�ּ���n���� y-*J+����'��f�L
��4���T��j�&S��[���Y�q�0n�*s�M�&�t����_�шS�rK����<,~k�NH�ҋ����G�Eإ(�'��'���?�7���R��/{נ�aCl�ֿj�i�:�����;�J���4�ͪ
�$���PD �BS���7��Q�Ny��<i1Z2��p_��|��(�H@��Y�<r�~�+�я��C��R��J�N#�;-[����(�� �����xv�]U�ݣ��	�N+n�#� �<�uq	L���
Q~�K<oJ�DCJTN=��lz<_N�J�_5tcO׬�\�O�T���K�\�.�j��[!� z��`�j!��M������r "mt3���Ku[��%'�d�Vtq�̜g���#ȳCoEq9�}ұ��lHJ�:g���^�����
7�\zF����7,Sڣ\RH�}��ppU�	�����ځ�%t�d���΍�a��x�>J���fW���Ç%q��z�Q���Q�Z�т���I�
qj��*���g��" �)����/��.Q�7j�J6Mt w�S��6�M哸���.��(����o
q�E?0�_�غʌ��3��j���Y#2��_����%0�����Ę�G��`�~ʟf������wx'�Пn�O�����ѻ�3���$�(l�ҙ�FI��
��Ta8~Jz��-��&�����?�,嗤Jh���ܭ�� ����(��}�i���o�Uz'���7�����"6uʝ ����^_�9�f�X��z!N�R�#"��G��|����v/Xcr���RR�k�=� �io�=�L,�P�ع	\R��.UhF5J�P;PE���_9��C�T5J��t��w�%����:X�"�༸P�����a *���E��gXƄ,VI�	1{��,]�#�H�/��"��-�&���4�TQYų�k��߭�1�gQ佱}M���mh���w v�g9�L��ng��� ������ *Ѳ��>��ǹ�e���{��
�Q�#���1� �"���RX9����u�w��J�����"MF�߯$&tXF�6��Cp|O������s��,eu��i��H�ε8܀	��=�][78�Ӳ���4�%�Lk�-5�.���@pb��Qj' �:����5%��ֺ&/4e�ǉʙW�!�����.:��Bu�A���#i#��`��&t�w�v��G�jT�
�6��7����6Ҽ���3Pt�}��\���V�0�Լ?0_Hv��2MXM��FȐ܄�q�g;
�*A��p�� �Z��7j&h�w�@���� �2�� �r�pĘN�9ms ]Ȩ�e�}�ʹ���N
=`
��_'�����D��d&�P��ְ�sQ	���h�:��1�.rP�o���,ꑜ������¨���Xi��ޯ��|A�:Ϋ���� �����;X��~XAE�0H�&yޫT��+,�K1��,��-V��=c����lJ3LDQPڡ�����3�ؙ�c'=��4��,n(��� "��O�0M;}��~T���L�`�����6�5�L�]��1���^�n�5į
�&A�&��|2ӷɢZ��$g-Lh�ա�<Wk:5�@[$�D�3E~v�qsT0l�X���+�}F�i.�v��;ws�zX�1���	32��\:�������<��c�+�%!�AR����~�NXX��+$FctD	�8�<�6��S5��XWj(ȓ	�c���6`¶�����܂5J�X'c�V�VM%�ł�$w��E��N�%+�A=�R�`��$�ݐ�۬�T��������W=C�Y��@��o�ћ*���$��;�x�"�yJ�*R���}�s����X�����pTF�����2��,��gJ@����m�x��J
�N�_��۱�Vx�
��\C�K(�1aHz)A�����\R�����,��p ?�5寚؁3�ᒎ|�����`��(��\�*��kI�S������ydl/8��Z ½����{��-���hn��=C�Fy��wyok�y�\����#��b�\g[��=��xCIF�O2��{^�D���e�%��m $�� }f���e´�X��E��	����$n�AXh>#���ŋ������B�8;цd�~���p��& 3PP��qǅ��{�t)��E��1auUl��Zi���bQ�h�!S:�be~_@�B�EwxsWg�-�uh��t��l	IKUY�Sd���7�*��)��l7�qhk#8�6׷�����s��@�܍B2`��{����* UJ�p�]w�y�W�{�hD��sK�������ܴ��1�"��qYU!*VS�5���LG���p0��Bk��9r3W���c�#w�uiƱ�h��F8����(�b*�)���;.���Gѣj�$���mh&�_;�.�f�&��ͥ���}voIS7�6'�xv��WS�h�
F9�иH���M�w��Z���\׈��	{k���*��6�t;qD�6�Ʀޣ͈$�[)l���M�i�,t�y�^�ZyT5��E�sh�ͶB��7�:�?���7x�_lG9�i�I��j�?R��:q��
Fh�6�n��^���u�OI&>hO�D<E_��FDVa�0/N}��FFc%Qpu���^n���c�a�-_�L��N�O #ؔ�OI�8�r���s�1x`�eJ���ޕ�/۠�d����My:��a���8�)��8
�*����p�hq�vx+��o�2�:A�5�94D�=�H��J��g�����;�v�*�/�a_K��������ם�?�I��������=�Bv�e�"�bg�8�9"(���&�c4���[�������/9n����If!<�~���t�墶�� ٖ+U+}.e�CZ@�p�<���ng�sT`Ɲ�I�̎�r�>5��D	����:�j�"�4����DXK�)}*�G��vm`��;�r�!�9A4�ꛆa�x��w�3>[��"���6���j*�BzJm�VJ�AV2�=m2ʠߕ�w
�����W�G0Y!cbC**�6W�6����j�q9{x\���ubW@P3\b�J6q�5<S�a�9�$G,z�XWK��)Y)��_u8����7�6}ۿ��1z�\�f����
���1�ޑ��@��v1)q��a)�G%�̀����w�����p��?�-����J��?���#K{�g����0Z_�m�H#BðJ�Hxġ�ib�2	�~k���p�#ȁ�q�A4���7���G���}8�=��������"m�db5����5�~�9/,⥑��HI���;�3 �����~7`v��<����:���t��[�(V`�4.���$2��N��$�/�u'�
X�-��^�)ܑ-��`c�9�~�í@i��љ�4�2l
\�d�����9��\TVt���-���-s�z�����5����}s����j��t�����$�Ƀl��9r���I�-��uEz������9�0��9�L�V3ֆ��^�}U�<\� x`��y`����.H`���N �qskP~�i�q�Rr����.4_����a�CJ��K����2�N�<|]<��w#�(��g�x#^�ł���U�ܟ.�����uiۿ�XS�h�^��i�U5�{�����|�l��7���������\%���n�7x+ԬU��-J8���>��4;�Lь���"��Zk,�������ឝ��#����W�7>�� a[�[ ��l��!ʺV�U5p/����3��t��f�q
�k��bQ�Đ�t�P.V ?��Y�i��U>}�W� UyʀJ�	��JK=z�q��Ğg&��B���|c(���"��n����{@Q�����6�	����z;X��ތ,q�R@}�)��4�񒅽Mz-������xh���q������	3]�dH5 ������2D�D7���e0?�V!��~�^!���9+�j[ ��᥷�V�6<46^(�a�7q�Y��{ �=L�4�� ��qs���M�3F�1.A#�>���א�yx��grV�����fi��j��	�Z���)o,��z���8e$�6��H���Y��([�7i����� �N��f�xQ6�7������Sk�k�TG��<��%K;�6GL��i���综�r�c��U��O&71���L�{M�<���Mwx7p���p������c��jj�滪��\�u��U(m��a�|�+~�����騂�6ora[���q5�!��)��[]W	�}����II��J�}m�@W�.ݦ��:�h8A v|��d�$�����u�hI��	����x�k�2�E�$.��2�Y�R�Lȅr�-���5\�X;�+<v�Ù}E\r����(w�!��� d� �۪`�6��}�-�~�&l+H|0��� �f%1#�ƽi��d�������[
1����=!8�ְ������>�I��"�~S!�R8O�܂]XQ�V�h�J�Ί�E	m`c��Ê�`�w��c*��w��mAV�w�y��q�]>��2!�`L�	T	�~�K�0}��A8fe�/�OW8+���ښ��UnO4�Tr<(�|�A8��h�t=�z�����JԠ�׺��X{����0�gU��R�%�y�VĝJ�t6�;�>mPg��L��_r�Y��U4����ޏ���QrT�,eߪ[��,�\|��<h	�D�������kB�;t���^��~�3iPM���)ZI�鎝�"�P�iQ,��.�:mf�j�fk��K.���Znp)z��f^y��Hm�(�p)g]8�Z_��VB���4bP�J�H�_/V��J��,�G�]8Ù3��Q��-��A�Q8c0w����b�(�5�Y�tE���If�ii"1����.����Gr�W@��ۺ��WҐ��s�� �?5E�	)b�8@�h��%B�������	�O.����,��BRo�4��=��BO֏�3�C�]h�0&��r �l�~[�l�"\��ӎI#�_$�1X����*�֡�Zqn:$��?I��h����v��S$
T*/�q;�K������h;Z��8.ԁ ����,��뾹�e܁��1�1�ږ����i2��S�����!G�$���3�f�<� ?0�ަ�������B�`��􉾒�C�L�"�q�,�P�P��M,x8���&��W�
�dy������j'Ix{lE�]�O@�Nb�O��qc���Z'0��o$��^$y��9l�/�<��tu�Я_��ʗOQ�F�<�-"��Y���W�{c���ߏ�[o!�.4Ê�Q���%ұ{C[��A�?�$��d2���z�!4��$���.v	�i[�;��-Ź~�KÆ�ZXX�䩀�+|GSZF�1�W@Pܢ7�2��n��>I]���M�棃��.�D|-W����ج��I[�"��k���C{���$��]�0i#�ٰ�L}�X��-7�'���D�V�B��+1і���?��ʝp���4R�q3E0�;r�m� ���i����2^��c�������ޑe�|�Wh���0�i>��-Rs������k�gC#��[4htF`�HI[���d�u��ǨiU���X6��kw���r��\�������*��{l���Y�z��.��kݼ|#�b�O�����Q�LD�V�f`/��>ԏԡ�[���B�(x�2^QZ1T�%��G�#�M"}�9�ފ�GQ8I��a%�2�(b$�Ny`�G�?(I��-��ZV����lƝAjX)�Q�Tt��d=t+��z�裶��	�Q\`�~��coSeX�Y83���+<gF6e���3I1<�	�p���J�$po�F�&,�(�"-�ui%$���� ����G-lN;�}�Y�FM��3=�W*��=*�D��~k��Ql�x �u:��t����?�����C����6W,�0��C�K4��"7�ү��?At�7!���="K�?J%{�$kt4Q�t��}�|'ɜ͢�L>���� %�Nn%B70 @���+�q��H/|�xp�C(�<Gi�����o���߂�| ��������͝T���-�?_��P��&���oh������ˌ�+�N��/�],�d`{�P%�o9�rnφ�9F������c��}@D��`��`@�IUS���j�C#��p|�_x䜟h�"	H�梥������w`��H��A܄Ʒ%�~ ��"S(;Cx^[�$ꩤ�&���{�����q��V���$9���ㆺ���3�<ng9�`�M��w���bV�^-z��\Fή���Sy�Z�����>9�f�s�#��l�1Q�aghAp~s�;�=ѿ�K�/�a�9=��y�p�a��icAQ�8�	:iFqn'>~�.ƭ:PQ��C3��D��i�ܟǱC$H��i�����YF��]�n��׼o<y�3<�y�*���3�s~1��~إQG������;�H���>]hOV߫�u����{,�!�
4yȋp8YMS ��dX�Fd�Qϟ�de��"�#�r^��	�k+HU.�U��}���8�+ �!g�V*�.�֑HR"�2��F�wLjNSJ��� 譤ud.\�e�[������2�\l#`�����x��>���'Qt���Q�����b��m����A��tb���.h��X�$d�O�(mf�U�9A���pDQ�7��x��O,C0�z�����\��&�� �ٽ�q��4ϯ�$��R����-Q�,|Ƚ������ce������`.~T�opQ���9ک�` ��M�d|��t��1H���!�m���i�9�2���6IL5x����Y#~m�^�)r�ol�~й�YS�.K����#�>e�'	�{&p�ŤO˥�������Y|��C��0����YӣN'kb�T!��K��n���b�[�e�.�Hq}aA���@gHB=�s��46��+7�JqƂ,��S1��u����y�����>����9�i���н��l��D>1����{��x��b~�bH�TD��k�e?�S��N]��VUMc����U��	cj�ґ��]��B��F�:"ð̉���$ 

�`
ٕ́��ն��\���t�������CzQ+�ER�г�mG)j|G�w�g��7Ӑ��4w�o��QtC���"
�����_:��ʃ�*�����)%�o�����}�G%رS�_�E��9e���5(3�c7au¼�]�5�e���(����1���G��	j\��1���65F�P�ȅz]�Ыj��ST�7��8�icu?�)�gaж�Gj-sݵ�\�/��Ăd�ضy�
�6�(��;�1����J�A���r��S�O'��B �A(+X|�*�9�o�0�,s���,P^˵'$�9�ڡ�u�͊�zD�<�&�D�pp�-45یu����;�ocB���	k��as�x+��o�ie~�y�|�x����9����x����I��}�.��t�W�xr�=7����O?}���Z�4���c�p�-HvO����	�˽� �g��,'�1�lϣ�c#�"Zd<���/�x��*A�s�N�'?q��
(mvCbw��a��z�j|h4Q��Mb�tQػ����:����eX�DN?��� <��qyR6&졒f	5>��0�$�N�_"b�����:e�=&N:�Q�I���W�t٫W�ΛU�-ii�����vz�{\kƚa����pGz�=7��5'^n�J4�z�+��l��h��
������G��*!���ñh�3<�Z�'��S�����2��GhW]݌���{��� ����(NS�cPh�<�
T �.t�*9��m]��q� 26�ڗ��%j�\�|�;އ�^�1'��[�t��aœ���07��:d�n�!{�M{@�X� g�JT�^%\��c7�+Xk޿8���V(�Sxη��f���K�;M�KLG=J���h�&g��./��u�F���c7�ϳA�\���u���:z��h�?�;�@��5�!n�!'�Y�f��x~u��kd�[��e�ی����)W.gz���|�J���~\���/�3�2ȕD8W�j�5-jv!����L�;��Z�q��`��u��b~�g	r]���Y߹?� S	HɘŴe��$�P����$��_�Y�s��`>����֘C*�ƾ��Ú'�ۆ�E��+�pd�&;����4?
����B�<a&�U!�6-���q%���̀7���裵���RbK>����?�f/�1�L֔�}��0�l����`�?���@��dT�����"x�y�� @�s��R�Fg�zv�~�3&��;Jk$�8�k �F=T�@�x#.�Ҷ�o���w��
�e�D@Nj�w� �}]��P_�����Ű�f��x�,LJ�X��@��Q����ަ2S�@�똖�Y�_��m5v�QsLk	Z+]L��-��WAu�
�b��{;�[��/
�M7SӃA�a�{[2Ɓ�	�X��2@ĲT��W�'3�~�ַ�:��|'��I�6}��[�C��$����f��!��!}�.8p�U&�lp{v�W�z �Ժ�Z�Φ����f�zy���~�;�?ۧw�
�:�{�3��*�(�G��C`�?�������-5�f�6l%2���J�s�+�+2�qq���'r�o 7��ࡱ��*"��HC�E?�i���ε�ש�o���n=��J\�B�7�W���h�3��M�J��*��/Y������������}�RU�������r'��P~ʵ��l�>��v�ň%$���Q+ϫ]޷�0?@�F0��q�nΨ�K�_�1ʓ�3���������;}V�������)�cUH�C�՛��y
 ���:T�P�<��cҚ֚ރw��2��N���U�(���m��u�j�����͛���FS�N���!y˩�o�� ��n�����"�O2�I;�,oq�[v�ʷE^e����}t��?��-DΏm���'�\��-���)����iONn0�_N\�,]l/睲���N������}�<,k6�d���X�xP�l8(���Wc�);���)M�Y �G���� ��R-��	��0�%����c�s�*�Sx4�/ٜ�5'V�g��b><I��~c"G�[K�8���m`�	մ߯�?��ܖ�|U՝l��o�jz�J�p���T���5b>�U���Df�4K�I�@O�~�B�~8��t-�i���-�C�} 1���ϫlZ�%y���kDY��8�0+�qTF}JJ��aGId��n�D�cQ+c2�C`�B�/V��_0@�u.5(�NEƖj��  7f�y�C&���<���
@�V@�H��e��O�qJ�t}ṱ̌�	�^�}꣦z�X���M��E���\��uV�n����]�K��3�%�BB��8S��>
��4$nπjB�<�Y��v�M�����!^/��ރ��;l���	n��ճ��Kwb8�A	9{ ��jX���I K՞�5�qA3��s^����oүW�V��>��������w��y+��+ޝ=����a
"��l�X�)�OI�������d�����9i��Kw�%1�5)r��'�����f��N40Dh� �e-��2��6��X��B� ��8p�b�q38�M�O�QF5r�h�Wt��q�a%u��A��a���Wze����9�k�UJQf��?�@&�^�1g�C��QK�19�&�!
5*��j�����j3�YPa�
�/�M��Q�Ƌw����'���{Mة#�Ty#�x������0]?��ܣ��*�3�]p�l���/�A�ؕip�ˈ�*w6vV'�E5�&"�y��Ӈ^��׈���h�����q��5�c3(��Ld|F�Nܳ���jͩI��=�T�2�F�m��7D�qX\d?7o���D��4��!��A�Lp�������K^�����E?n!	�Q��Z�m�pV��ˣׂ���s8�=�f�Xy� ���o�8�=8��`_�?m�e���i�zp%���W=/ZC(�i`���5"ǉ�ӧ��������to���|Yn� ��h	*�{�Q��	e29�q�BQ����a0�ܪ�R���VU�0*��|BKjUk
3�_��c��B�W:��EI��^�q�LnR�Ft��;£D��p���Eq-@WE���Yl�.Ĳ��ٍ<t �膉Q�%��iT����Ӄ���hP[�S�S���V�S�F���;k�����=����X�"2�Z������	�2: �%pՕzX�D�ʉc��K����;��~m'y0�1� @pZξ�ywU���vÝ·��S�Y����Z'���^=g��P�0N���Ņ��FEs�+�[��Ku�BI���I���	`ܥ��}Ȋ���h>��i�������^sX߻jjx�s��yP�5�P^�_b_�ٳ'tX��w��e�#JPܡoo ���ӱx� �^�z�'S��m�i�W��'҉�	LX(s�����C�y u�[��b!m�.��w{�|��C��+#���U��@�5/C�>�����'CS����Q���B24	kz��F0]J疢O�0$���E���Ph�<�+�j,Zcn�XB٩�L�{	�Җ!�)�����[� ���,H�Qu������.	r�@��l0�wҎV<���!{�
��R�YYhu�;G��*�E�Y�4�L�ӦM��"U;�Ta׀�m:z1yǃ�9�@�x�o�I�*jA�1�F�=Y�"�c�g,�������R������Ǔ!�=�Tѥ�.��Tx��Re�~�i5P3�򗼫g�9M>�֗m��ή:�aԽX���@/Cڂ(��񓱖�;��xd����Z|X|��)-����)aq�����Y|3�v���)#��vL�''��YE�\@���~�^+u��]�nj��Dg��x@�B�0Ih�S+�5KF�f�2���_Ǒ���n,��W�mM��V�����(?�sU���|&�
��LB�J��uR��\��t�C+[��� �SC=��b�:�yQ :�J���B�=�\�g�k�)֡~��t;�,�и�J^���w`�Ak��}�Qr֝�'��='`~�w��S�`X��ﳭ�I�M�8�!U�s���M�u, ��`�WX���{�W��P�6�Op��ُ)����}�^���D��D�rP��&s$�J��
�85N	���I0�"P�0�[�`v3��?0�o3������5%Ҿ���7&�:��Ug�� ��I��{��M=G&�����q�zDL`�>Y��}<�DBh��]�V׭�*S�R��[�i����i# CH�v�_$n�-��R��z���ޭ�l�nN��a��`����,@�l�}�[.�D*u�W��c�<Q�\�2�b-�'Ɍ�9����S�D�DQ�,��̛�q�lIʒ�8�k�]�����\b�u�.��-���J�	���;�Y����$���ں�mM6�%����l��9�U�@����L8y���g<�z��^۟�/��H�;W��+A��,͋q����`Q���K6G#D�\ )�C�x��B�x&7�ۙ��~��e�!������~����(�WP���6���i1��8��@Nq����P^�l*�O�ctWGLR�:T�l夞��jc���89���b@���zA}�~�(��w{��.M�d3�[����!��8���Ƿl�$&�/��W��%cA�F��	��˽�.�#�_�Ƶ�<9�ޒ�{����p�ꢧ7���-cA�ly B���t�Z �I�V��a����3�����8�&�������qn��M��_���̃�v��FvU&p^��R3���_AZ��X��ZMI~��#Q��p�������KD�L�L�2�Q�I��H���'�;�p_q�v�Q�DG�X���ՓW�x�9�Gy>�������_˻y7����C>L9|�U����=j+"�b����T��-m�;%Q%���Zp���m�`>$7���߃���T���)�獋���}�\���DzC`�|P#�,D3?}$��{��9����~k�sJ�O¾��b���Þ�?�$@S�1��5�,�:���^kdw�P�|q���b2��K��v+��eR�r��Ɩ~�st'9�[g�+,0�M���ȥͿv&I��C` wG��~�� j[���w��>KlG��|!$e�b%L�� �7���i*�$W�x���`D��5)&����]�^��y"Q���i��w'�{>(o��`��0���ӊq<��D�Ҥ�P�-;�z�$����OkM-22��bi��*es��j���KO|�.@�=ɯ�/�A�,V{Gp�:m<����`Pg�c�a1��z�4�hs�i��>J�h�6��#�5�2����!"�x#p���;J�\�����)�H��&�>�Ոb�c�S�&�AD�BO63�I^�m#��~{J8-ф~@�N��֜z����j�æ��rs��#k"���*���V��/ ;ߺ��|-T�"9 ���F�A|�{�vI��K�U<��N�SNzԙf����ёf���IJ��L����]�r�%�a��U��� 8�0�Յ�3U?EX�������+�	M��U�������L�ܽq�7�k�
���
h%YTH������77,q!��M�yV{ �K���e����*+Hi���T̡�#"9%�|v$��/�'�	+���'<�)��>��{�V�'�O�0��j�U��zjU��Ϟߪ#5;W-�T��G7Z;���f&v�嫕������l�[:Ի��X���o����3�Հ��>n�_�~�\���)��������.A��j���BDV�vM!�_	�?py#�l��^������=���8#���ĩ�b;C�2�9�5��q9	ڔT{�9Xh��f��S��n��s޳tjP.aډB��w	*W��;{�?�0Q��]�P�I?f2�yT}��Uq��������+^`hA!�C���!$���i A�0/�o�5�{������2�����H�ϴ�T���\k�u�[2`�MmO�2��ӵ!��G\�l'���;�`�|s4�����=?0O5'�_q@�vC����,-����=��x���o'ء�E�	����9WZ�$l��p>L����!��/q�r�v��X2�$e�]��x
YS �:}�8��އ�[#����*������5OOMB���FԄ*[� V�|)d��r� �,ІC��U�A11��ϋ׊O�u��e��sZ�0iΌ���m����D=)�΂Ӳ7e�����H�ɠ�sb��s{k���3��X�N��GJg:���L*q�ޑ�7��ڇ��Ap���9{��V��`��vd�q�Q*��:�Ɂ��� ���vV�V�)�����Y��<��?�$`5���p�MGci�v�������®�����M�͍^��-/.RHB÷�{��O�&��,����=+��Y�[�}��X7~�GG�3f�Ϩ٠�!F- ?H��J��E(A����9�]"B����N:�Jf(��×��4z�C��_�Z�bp�D�,�~87�(���P�o�<��M�X��b�m�����1�T-dCpUéP��F{k���\��4�-O8U�E��%&�����Q�FmW����g�Hf���k��[�z�������?C�1���%>a�?Du��%���Өr�1j�9��0���࿼k�hI>��],�x��б�b"��?o�2�v<��y?G?�3<�:��l���Ǐ���<򚣲��[.A�ѯ�N��ŉUT��Veέ����|NP�ԓh6�h|!-]�Όz�tb�|���u�ч�aN����Ȕ����X�ԫ ]��&>1�����w���"upx�et"i#�XCG����A�:YT�X0��%ǡ5�[8S'a�C��5�f�Uvz����e���]8sn�f�=R�R~���9���w5:���o&�A>}OTnFi�E^�ʶX�i*�Bc�u	<�X�<��lQ��z@���-�5��3w)�/7_T����/�)bs~���)�(� jiq���x�ș��Ij�S��I����"K����������\��q0xl�b)��!�.H�:�}�6.�����?}�N�M��=�A�8�52r����f�E�5�P��|=i�R�@��i{�V�}�궔l>��9W{kj�hp<ɖ>������e l���ro[�K���vD���uꡡ�r�x����`�dM�6�ĩ"�!�p=mA���Va� �\��{�Y�*�M��^�9���W�DC �5�<�����J֓��e�՗7��m���Џ1'K�MX��F�Ґ���kD������1j��S�H�q����!��7v{�Q~���k��#���Q��q.sڔ�)0�5�S�&�Ww{����½<��Q0���sZ|ȁ���#e_�Y�'�}����pء�B��ZBN��z���	hx��L����3^�I�앹Q�J=��P^[6���,6���"�&�5���\V�É'��o�Z&T��2^�gw�����-_N)̓w�E���f�*e'���_�>K��j��v���c�V�H~���'�p��زH)n5J;����r�TK!0�B؊U��}&�.@��cj�n��V[W�N��z/��ҘJz�����E�D�m$Y��/�{�\T��%ڋ)�����,LF�kV�Bf�������<	¶�׳^,�+�_=��GQ=�$S�w�����;�$�Q�l���c��qO\Hh�y2 ����s������e�<\�@�3�8�ez�a���\�.�a�Y�@�T#r��b܇Xr�D,4jג��gA��/�Ĉpn˹��X�k{G�����=�鶐"Ep*9�^(�ʢ`��G�>W�}Ɉ#�X�߭F�Ӛ���+���	�z1��I;)�^v���3�1��M�,��%�v/��/�}${qc%ٹk�N�zˀ�{P�6}��|���S_,p4���^��K�fSaK�t5i^.k����S��Ya�6w*J�(Hڎovt;����j� B5y9��s6M!j_2
�_O��>Q�1mo@c�;h���m,�)!ϢOpywC����7����$���~-��jpm'��4bf���%%�	���� ��JJUb�ޞ.Q|d\���~�硲8kL��2%�� ��߰"PS�B&��n�M?�
9���	���w�!�1�����#§��*C��3��c_�J'n<Ȯk�Z�5u��x���u������^p �������5��՝��X�Oh��+_Ļ���{lYIj�͆�~v� Cm4l<�g�Q��T
|�����鵓y��1�\��4���!an(�B��4�!74��i��Jl\Xk��$,�8����Y��9����F����]�"<�Ѹ�o�_�V���R�m�^g�N۫�HA�Of�N��v�u���^���̳��L�i�sg���ƭ%�_P`�|C����KU"h�Y�;�P�����|&&�o��n���w�mv�9Y
@�w��&)?�5��w��{/�h�����0=u��dc�[	�EBUW��h�dLh�.�B<@mO����R�j�u�	��u5!m�ޞ�
��-�/aU�C ӆ���k��^���֢�)#}R�K?YB�EQm������^h����r������XG&T)��-<U�e�e�]��!!��kα\K����ϴ�g�����)`'c�̟(0����q=�������O�<��K$:L�(f���܃ձB�|��Y�fHI�������G��.�=�����f��'�.�����2IENʴ��$��9����۽ם����^����?�d��Vk��d�f� ��t仌,��ˣ��k��X�5م�>ɌH�'���_jԳO���i�I �sG�9��V�j��s����R�������<�<������Y�������賙�~���$�Sn�쏩�X8�!@�d
�>�C������+�4���������nmm�����Q��_iOJ�ɔK^��x����UKB�Ή�	����҄��<�Lj�ժ�� hAc`����vh��ySf��l��(�B�:h��J���I? �-]�ȁA��qR-�� rCj6CWU�;V�Ǚ �<�'����8��Y��W=X��"u��CV�<xO�Bs	p.s[!6qk��m| ����
,�w�=d�%�<�Ո6n%�Mu���YaS�F���r�{���q�kb���}���Q�޶�8o��o���>�"�;���^�5��o�Ob�F��di�2���g,�LM�gI�����[P��Y�hde��X�>� ��D�ܥ�'����ݗ)��{�3��fYB����~
�V�9cRp����5b�v�c<�D�m��zJ��<u>B����q#���/�Of�a7Ѣݞ((�{�x�y��<}�D�M��J�� '�-�k�s84
��t�%{�/x�
�Ҁh��5r!��!�O���=7Iƍ�cG�xJa�:_�����o��'�.Ơ]�'�C�k�{G;,�a}����^e�+UQ��<3X���@p$
�T=���,C����ᄒJ����K]]搛0WS!H��/�usLWږ��A%�F����گ����qGk�D��T>�eV(�c��4�����AX(N4���d�X�p�9�7�
��vLh��2z?��А�X��VnL=�Z��w�~2R������e&1'�D�i�6�\bӳN�;Fy�s��^�������`F�1����`,��
#z�ˈ�^���a�4+������$���i������@�:"Q%���Ɋ�C۠��8�T?0>l3;*1V���,�4|�}����5���6��Ē��(��,��P��V�I6ζ��}H�f�j�C�TTX^w<��[ 1���ST��=����c�<ڎo3r���iT�Î�N-�9��$�D�)�����K9KQb\ac�a)���`��/�K7{Q��/���Oɬ�]"�����p|�%g¯9����
�G��j�*��s8LAp��<��e��k�!ĥ)����H��<��	��3����="5�7t6gq�w�|ܭ�YA��,dҙ��q��Dŭ����RX��-藿Б���x�������1�q��85U�N���S[U�ϔ�<�gȿ����+�5���B�>�V���/�!��4�@�w�+·�VwprW�ۀ,J�T�~��`�'p4���������Ůt���upJ�Fz�}�p��ԍ��8�lw��K�4�B[��}/4=`J�iߐ�a�Kk�S�-G��WV�3�&�=�G��2�vn)�`��%�����b�Ĺ��$�sp��j\�q�0����� @�E��<��6ᖫ���$Q�\b(���*�J�wʾ倮��vbH#�/���O�OE⟙1-EZ�id6���J�:FL�@�l2��8���tu��i'Q�j��}̋n�N��<�����hN7T���`����Lx��/���I@s�?�	;U�4��=�p���
��o�<�������|:z�>��j���d�N�/��d�]S��И��E�KsH5J!	�U� �epwP.�y����l�$����r9���]�ޓ*�"@o:.��YEꛇ�"�K�Y��jQD.�4	�c�xgu]'��s����|�B�}h�	��g}$�2�A� ���P��~g��|���3�ݛ-ej�7����i�Ly]���.��c�E����V�2� �����>�yym|��2R�r��KH-r�"m�ܙH"i��t,�����dR��,'��I�}QCXvn�ҋxا�􅝖���Y���3�ö�?��vAºk�j����
�U	�><�n��
b��+"d}�U�:��.�=�<��3�3_e���S���r)�&sE[L�h>F�_(��9W�ٶ�v$`LZ6x�S00zy�eC�f|L��9-�H��z~Ie臠��L +G2�;j��}،�	ق��:`/�V�ɳU4}������1�\x�n/ɛ�������?�������~)�؏F���a+���/��給p��M���Q~�( 	�����!UE�$��#��N�Ua���-;��Vxv��d�GS!B�xȨ�b�����a�`!'L�y�PWю���e�MKvj���u1n^4����ڋ�7� �)�̜�s�g��1Ok/��F(�SLtx1�dz�V�|E	���Q������>��*���)���ڭ��v<�9����^Af%u�z̀dB�Bw��<Yh��cL��8)�0�!Qݥ�>>3&j�T��Xȶ��칽�c$`��@�	�KN0�
$��D~o�8�ۖ�_�i45�E���9���z�M����]��-:Hٙ/y�.^GV?�ܡ��l��w ���K��ԛb7���G~���9&�	:�<%�/I!WΜ:���^��*6Є[ƥ�E�����B�|+�'�T�*ҁ�Cf(��P���W��W�!s}A'"�*"����p�5�}qe��aC��} =a������{���>�K1j]��I�S�����?�6G�j�cZ�)�2�EK'=HE7%t!���φ�:�7Z�_�����Yq9@m�;Ȉ1�]gaf�dA���w��)�0����DG_N]��_�� �[�d����+����K��Q[Ɣ�ߖ|��f�o�]xcѳ��{3S�����8���ʸp܆y#G��yx�4 �GS��Uq7��U�D�%�Ӽ��c*�(������;�f�޿�uAs[�`���^f6�W��2�����`D	K�8u�����'���9�p�9���X��m����Om���{��e�]���g(,��#1��Zc)jT�	�b�PהK.b7[_�Y>^��+Q�1��8U��a�,<���s��!�����٥ϸ{��v-r�j����R�Z�3��z�~���0l�ϼx��x�y6��4X�>X����JZ�t�J���J��'���K��������#6/��8�v+Vw�Q�]N4�kp$�O[*w@��"O]��^�G
��!�B��5Y�'5���z�{/����IE�h'���<=7y8��.ʦ@�4��6;�N��/,
X�?�<�1�z��<��Z�K<L�!���ٸ�Re��m%�k����_���3�V�q{�v`��W����5b���>�����>F�ض�8��F�yed�{��g����Eo�W vkk�dyt~�N��|c��p��J�.�����R�����\>wm���C�zؑ��ɐB�o��ٱg5>n[�wd��OsM u￉�m�^.l5\=��i�B
���܊6^U�IN�э��/�d�P<I�d��#�~�r�IvIb��=��Τ;�V�^�~���_8�3�y��f,>��*�'�L�kZ���G0�^��B-|'e	{�x׸d�C�6c��yZSdv9pg��}�n}�����
縈��݁����nca9'"���nN�z�W���tM�'{���|Y��u/����r�P���oT��U�@W'n�}?�����r��H@���-�� �fIc�@Rz�j�rIu�V̩"�C�C���S�i(���_���̽9rJ���$:�b����d�1;�VM\�l<K��FKuI����G�R���pgP���Z	J��밹$iQt���"��v����c$��{*�k��zzI�� �ՑD���Q+�������l��A+F�q��Z4���>6HFj�%���vC�z������Pq��QYjfԶ�B��k���	� |�2�ۏ��A�OG�B���}�V�jO6UF���9�@&�}�����|3Z|Oz�ȼ�?�M�@�e�"N����A4�4F`�c�6��!�a�t����pc���^Bp��K5Vq�"hA��:׿�с߰�R�]�����B�Y�?��Ν"��Urc�@��iy��\e�s����$�)J���Df?��7�ZY"���,�Ը��d[���� ��FٴLY̠��Pk�C�����I	�z�뉋��<xX���'̱ ����L	�K�5��oTz��ׇ�����ۙ�!�6$���.��p��	i!���z�aV��juf�{�3��ʊ2Z\�\��_ �s6G�}/޽Ý;��7�Dн�'�"�C�>��R�叩�~��ø�c�8��+bp��3i�c$*"TeQ ����ʬ���B��1������P�� ��a������~��<��{s�u�%s>���ѷ���i��g�G�н��S|���٧��F�I�J�	o,|/�3��f1��҃^+����wo �G
���[{���ݾ�
ŧc5�' �T�H��\�fE3̪���j�:�Cd��uDF|�?�I���z��¢R�6?���l5�����>7Ijh%T���m%�9O�N�C��E�[��X�b��餕zx��o;���%�PK<[Ý^Î����NZ7�W�ٺ�&�3~���]�E�2;�\�X��P}\1J�U�J݂��M�mL� X���V:��;ȭ/ｗ�ur��1$��Ď'�u�ܓ���SC�Ltٟ6S"�bT��L�j�M�3�PWD�$U��G�!���&�kx�wIj]���0�+7Vx����]#��*߆�����+u��-5��u�5oп��hz�Y��ޗE�d�p��!Ȩ��ܸBj��R*5��A�$CR����Ţ��F����,�~�dԹSu4���Q� ^��z�o8H����������.U,��6s�oK:a�W7�8 �N�rY Дr�h�p�������� � �$~����_N.��J�y�ڠ�:�dpK��3ڞ�[���E��ݩ�({�w��\au�Q%hd�=:��K3�z��Q�׸GqƳ���f+~�r���7q�h�T?����s��*���H�{�*ȝ^Ƶ�M#)*�w������J���n:&��0)���'<�5��e�P
E�������:������Ƕ:ז�K���m�l/�ȋ��9"	�h�sP�Ƴ`{x����W���@�ْ�O�$�")�� �W�3V��;w�=�Te����/v3BW�цPNa�I2���]�F�BJ��H��k�����x��M:mm�ۧ�X�3�r������Wa	��&��3w��Y�̊dYѠ��H������Y,Z�N�TE�&(���T,�~�I7e���$&=a�ə:+�uJ�l����'`�Lk����5�,�`>O:��eI���m���/���)�N+�t����;H���t�4N�=�C�Q�f��8�kĹ=3�)��Mp�Wèw�8����*���K�j!�6*/o��;]�B����v��J�՝��o$wm�H{mBgΚ�x��4�y_l���3��;��f�ϰ��,I���W1UK]�xENK�!�b�A��,* ,7�1��V�(�<�Vss�֡X��RGZ{���ES�a���~�_�� G;��~�i��4\
hs�5��*�i���m��H�oݮ�.�H@8�b$D�w`�D����g��rOi��ev��N;	��E1H�����S�w��(cLtuE$�ɌԿ-� e5(�ƙ+�7��<,3��}Fw��*���?�ˆ�"�g�hX4x�����Ϧ�ao�