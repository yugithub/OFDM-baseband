��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ �V^���qQ����jH�I�
�!�Kq�y//�`��~t��
�|4-�N�ԏ�:M:]���UއE���#J��;��Gt"��Z����/i�K{�d�n�=�Y�7`IpJV�,��.�ϣ?��ׇ����f�P��&/�Fkn��v'@A=`X�D%-:sI�nd��I�K5
���ҷ�֜D�=��?3�C���ڲ6XO�H3�%YD�k�<�'��F�����`���OML�������:�Ǧ� ��3�5�l��w�""�{a[@�*b�Mo�s$[�'�P5��#�
�v`�?�=A֧��]�{S@0�3���F�}��0�]�R��'^�s�h��"��I�%<�*N{.F�~BO^�^X\��D:��"�\ٖ7�"{��0۝M~�Q� u�Pc"�o��T�;e��Cd�@���
S���/5\L�8w�R�el�5p�z }v6*
/�!�8>�v��N�gr@�4�����g��O�yl~H+h�^s�3�׀
��N�E���)�{����m�S���A�g2,�H�+�n�h`F��q���N�-Ԃ����Ϙ��mԊ���H%��gL,�]�Q\ڲ�u�ȋ�N4m����!�{�T2��7��c��͚�UB�8,Jw�[I�tĈy�Z�7��RJ.��gfA�R�� IQS�4 +p#�ݸ���Al?��0��r��,��� ����=Fs37cy��yu��d�!�D�
��`^� O�-b!fApUH�o7x.��͔��`1�H��3�&�n(�b0��蘼R���N3:���X�WfY��HT����e�8&?NH���($�Gh�ߒE��4Z�V.�%��K�Ha��N_��Sޔ\�bHu?ij�����q<0�X4��U�Do�!��Ju�rR�`��}�E���H�^�bF�FݤKWG��'�ǌd7��
&�Y�K�s���	rE�������mOȒR,_��0@�����%B⟃j�x������X�Y>c���@T�_"/W��1k�PB\u�;�kX����I=�0����h�˖�$w��qv�C�Y�=h^
��"=Ik�&:>�_���,l�aj��L��X��#���ӕDr`�F�h����i'a0t(k���'�'�HNd������2���:��'8CN����fL���9Ru�$�ܯT�O8}ɐ,H���R�R�-Bb�uaD��_�"�N�ń���d�c��｟�=#�����Ĭ��شGd`h���ܜ( ��^�**2^�O�L*m�S�� 5s�;5UG�W�&��R��)O,�<���1
�:L�xc��IŒ!U���d�+�q�k��,�m�p�!�]� �������!�Z=�������M:!#j��P:��AT�zdQ��nZ���M
� ��h�W��� i@vQ�χ3_����c���[ܼF��<5�^J�X�~������^��%L̩I1�Y��)�q���ɝA�:�!�i��O[�壾?���A�7��Ԥ�M�Mw�%a%�/E�	`{�����=�,Iч|�U��C����p*�wx�[�k�h��)X5=r5��߰�i1�B��_���7-��2�1?�9ca���r�1�}�dF�>I?"��� e�eͶI��D���l&:7��Ȧv���~�����-��������8�Gfb�����R{�`�����S��������D!����Є�$@�XZ��g�'���N��
(d#���먼N!��10,F}/���Ņ2�5�t�K_g��� �b'�?J ��ƪ5�r���t(�5����mK��J�k3b��1n
Tw�� `�*�|ݞ̏fi�7���f8��I-�Wo�����WD��Ɋ3�l*�����g�c�pU[�8w�U3(��Q��Z�Z������ף���Zܗi* ��У��!�a0ET�4jh_��������hO�����S�{�jjG���SS����:$���OaD ��#�ݭ���s�4t�������w�'/IKL�Z�}lSN���Hܬ@	yJȭ؂�Uh1�JW�]d2��FVs ϊ�4,5��M�?L�d�*��@¢��&�N�ɮ���5ū��D�g��!7������T$�d�i�71�a[.,�>Y��ڇ��?CǔI9\3Cl)ݘ����ќ��;�]����U�PAȆ�"�-�_|��OÕZv�� w������(��)�_����e%wnI{�l��{�)	ir���CM����PA�i��X]D|W�Ƥ��wdD�k�)��֭6.�V���n��(��u�Nmj���r/��m0�.#V��u6��{�E!qA>l���C��&c�����v��FY�ӻ�˾�h!���D�	�-�����CP+�h�K���M0�"�yCC��ޓX>��\��<yL��s�R��8 �&:�ꋘ��=�Y}{�_Z��{�#O�����^�/y5ֻM3�n��?�.�e����.�W����Q�E�����7t��
�<�������U�{c��1J�M���{�5�0O��K�&��#�A�[9��3zr���3��+!4[�k����o�c3f�wZ��E�&������!K��IB�tN�WpњBh.�!�`���p矢��0¡
��=��c|�-�-6s�z�����_�׫�}+��dN���J~Z�HMJĝ��C�Eb,O�ʯ�\!C]��7���HE�)�v������̆g���8�Ŝ�g��*��N)/&5hÜ��Mm�B��0rY��$ʚݥ[�&x�l�$L����	�T?��p��rV�1�h��%X��6�6 2X��T��zC�n�Of��]�51=��)2K�_rre�4!q��d�F�I��Һ!`�v\M�|>����C2Eo4h�a�!�ɐ䈂y�KE	��\�Js8��jj��|�٨�E�l,Cї��e�T��$ME)���p�V��Ԫ�̚QC�,�������%vʔ4������hv	w'�EE������tm����@e��V�Rʧ�^ٝA�N��������j�,[;$�U8	��$���_fu������;O���6� ������=�|�~�D�3�%p0��E��Xb��t-���,$4��N8�����3�������{�5�`�_���������Fv\�*���Zջ�a�dH�1���!������G%�de#�{T��7��^i�k�q�˜G�m�}R�E�U�ӫ%x��&�9��x
�l�k���4��;���c�V�\��닣c�}7����"<���Ȱ��,�\/1𖺙�ͺ��?��DC�kK����}Ci�����l�&����Tν:��2x3�	�:�����������MgSp��\ȁ#*D�sĺ�����פ�7��1��1�X��=��F�"�U��H�����}7����E�%��E���TnQ	�h�}��#�$ݯlJ�[)Ra��}{�t��a6j���y�-*bh�+ʴF@�zDg�~*�E�Rd�Ht�5�Z���>ˁ�m$�������HG�e�S>ʎSo\=�>=�<=�xl�{��ñ|w�Okf�%:��$���Ks���4p�3�J�)�؉���y��O�C�̎��ӌ�f����U��}��BP?�`��ڕӘ�����坃*�|�,,[i)-5�nv�v	<[���PP���i��S��� ��?N����YD�fj�x�u�qV}��yC/˿�F��-D��W�«�R�鲴h��pW���n6̙���X�9���5�r�\���op��4�]n���
g�jY��`�O"z�S��2�L�Ŭ%�U���1m7,^�/��t���>��p��3���Њ�>�}�a1��'�-5�p���k�sJ�U�|�TI×;P���f�i�[x��#���4�� �`��_�qp���Z[��|�u%�_},�*]<*%�J��a=�ي�eI2�"�x3Х��'��N�ߡ��Q��
@�a��Ѝ��e���	�k��|�H��t,Ax>΃;b��`����U��$�6ѷ<��l�;Ϩk�A55�#��;;M;��b���9�߸me<�1'��:M%NJ�wlj<���F��Y�s6�Q� �u8�o��l�YS{M�"m_���7D�E�1)��D����{�Bi��,��s�B�}:�� rR8ܭ�Q��죗p,�G	��y;�+����kbE���˙k�pe���#�l"�U�M+r���jN��"w��I-�G���\�&��w��F\`�P�$c}�:�x;�B�\�9�r(�A��<0�#~�E�"~S��A?ϖ��և��a��7�S �a��&��s&��y'9=}(����]��[�;Z8�貝�H]	^m�a`�e��2F7������Sԕ'���$��u��2�����X���E�v[�#��<i���9��]�#8\��Y���Wv~��:���NVB����R/��*��1��c�bg�ӟ�O������/�Np>���e��tD�\� ��c�f�Z�?�
$�<j} u��bz�������Ɠ����$!;�ƀ9&�9�g2�E����pLh|$5�:���6]���g'�3��7�d"Ujfk�L�:0ڿ��&�x~���Z˂��ie����
�W��oF:J�,�6{ͤ^�m�^!bְc(�PNݰ�l�C�λ	��k���`�4rn�x�`_�͑{�1�Z�D[�f�B�(f�8�['c���w᰾vB�^�)Y�y
x 0�,Yv��2�	�&LKIE��{J���VPz:��W�@�K<�8
���ގ��4��3y�+���0�V-`�850�h�@�@��C�R�?�y�0*���3����sib���Vn䨽V]������S��$���F��Ъ,J��k_}t躻6�j�GC
a��% "�c�ԣ���N�srv��ub@�]Ub��kB�kh|_�&H��W�kƼ��G��'4L�(�ZG6�CRP\[^��?��	WЖfs�΂���_�5��\����/d����<U�y�ۗM< �#�~h��U-����; ��,��t�'�Ơ�٪�-�Zq6�D���n�֦ؕT���F���d�d�F����f��Ia�^��ƜfS'6�Ӗ��_���G�2�Pd�Ƕwm��zSަe�M��HQ���y�y����YK��t��4�銡��is!Ѡ�۵�A�ԕ��j?J�I�kk�����̟NGDZ�ho��|�F'j�%WK��6��"QJkT9����h���/����I{7�~��l�I9������Ǵ������5�m���������/�`�&9&o�w��a��]<b��%w�;�9����̢��*�;Y�TʨF����(��廳��$ۤc+�Z
����?�*êߴd\���C�l���K��H՗R�sA���������F�M[ю���C�;`S ���H	�}�s>��15���5u���QMG��wbe��� u��|�܃p��őe��}�������\Y��[�)�>�X�C�n0zN�t�m�u��:*F�L�{TĎ�5`Y�άh"{}��j���.:�-�+�M ���X�Bϗ��zE�d�I�
!�$]��$�oJ�B���3�Z+P���:h���]�L����F1����sz����H8��C�T�E��)cKΗ������[���'�������1=e%�u�[�iX9ذН�D<����B�i�+6�F]0iÞi0��͎��bCm�B#)O�Vu���	>)���a�F)}��V���$�������>��:�#DT��-�?�k��䴐��w�[~Q~i��8�0������*��.Kb:�ǂ�dvuo�e�����=4�i��$�0�UN{e_����\rs��ؗq�x�v/�-����%�@73�����@I�mf�����&���t������L��;�`f���8W�w�ЕN��~;S�z�UU�W��y��6h��?���O�#A7�^��Yʤ�2�OFʑ!�!v���`8AKN)�l�������v�ptSx:�f��ߎ��%�u��K(?�:�� S����=-�JL+gI�u��pR���H�v:���L�~X��ϒ#�I��&D~n���1)DxF�f��G��z�A�^`=��
EI��QY�NtV|��6`�.=�G�8�iV=4�� xU��
��O��V#�l�BI�?M��c29U$�\蒅�P���*rYn#�e�?�u̖���q> ?m�׆m�)���e���Sa��O�5�/b��Q
{a�	�MhO�T9�K�T穀��a��Ĝ`����
�B$$b�G�g����^��_�����-3q����Tz38�~]�EjǷ��g��.]�b��������À�,������W	�HRI��O��p��[5}Q��,,j�K:�|j�¤?Vn�Z#5n��&i����IZ
�؈A�/���PR�j(�����ҽy�s����/ީ>���MCb+y���sgpN"�Rts�slʹv�bׯ��za���b�{�7Z��:��	H2q���ԥ�Ԗb0�"�?��q�]/v%h��u�)�X~h�'�=XEn��L��>������r-����(f���#Z�R�!�e}FQ�N�v����?�
�<a����WV�^S�]kF6RAa�\P�u���q �آ.�W�ǋD�[A��[�z:�nxYŦڊ�miL�a��v�Ä�E�����K�]��������/6;�M�7X�L5j��(�CB��EM��f��n��l�Wp9�`����Js�,��b�p��e_[�z
Q��]��LRKA5�Qɂ�V"�{�J]�SN§&�e9���G�3!��e�W�Z3��o�u6�
�R���͌��[�s����v�ľӴ<��Y���~�B�v�Mv\k-t��}���}.�=���L���#f�����Z���辶���"k�^U�v����S��Z{�ֽI2��jrwƠa��#�Pz	0� s�󳨼���ۀ�yS8̄~��W$�ԕw����A�͔Q�g�h��� ɋ��=��xT��a��C#O��*��x�Ҫh�����_�����I*�K(W�A>9�����K�[� ��|�<�j��J�'���6��T�򷄅���	q�npiY[�a��G)O3{ؔ9�`綥�ARɽmp��C�:���m �>����x��!�e�~�}y<[F7�]���m�z���`��'v~���m��S��e�̩`�s����DS";���rb�=��/�DM:��hޅ�z-�o�Y�,>���n�?a��=��kk��h��|��G�(��~�O]&j�������E�ڠ<Y+����0O
>�=x���/��w��>�GM�Bjt*e0���L`����K�,���
B��+���_��;���il�p&3�c�K�"��ZT��	P�ks#���C�I�c呧B�sz�*�R���!�ߖ��[tU(<2��������5k�W4�
	O5�]���%�[�|#>�ώ*���#i���ļ�q+�e�0?��r�:��3Q=�[��r��xѹf�T�2����(>T����gC�����f�ޅ���G}HlQ�'�j!|S��Lɥ��W�P�&M���j,x{lsM`�3s�e���?ӧ4�}U�ZJ��Ʀ0S�:Y�H����Kn���`C���