��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ��t-�Y�n�.>�!ɸH�*�o��h�PG�J?!i|�Ws�����gG�s6��&(�e��U�ހn�p8D�~���Z�#�q����ē��1���˛5^�ɢ��w��f�hW�l��^����ĜT���*VkէL木���G+s2OܶN�f�v��m�eǴz~4N}8@"�����G�:p��+l��ä́�m�n���UV��7�Hh$�]����5XN�\G�����Q�s:��	�|c�� 7�b@x��[�,�3�PN���{S�9{�h��ӥ�����3�%Xn�;t��E9lt�z֟-d��:�Fch�IW6�-]���Z?'4g��n"���s*=n��mf�Z|�a��'��s'6q9:�������G$]��z���V�	����6��n�}?�O9.˻��4��	�v\� ���L��fo�zO��r�'Y�=&��{�{G��8���}��K���tP�:��9Ɓi���%%�{G@�y|�g�(����*�5�]x��ROi�
A��o$����(�yO����� �>�}AKpl�Zz
��������N�Y�X�����G�ʄ)���X���ݏӢ��$�o�p�uL��:F��׽X�(��d������9Tv�4�݃0 "?|�6��X��8�&l?P�1Gـ��1���Mh�L�Lb�N�@}_Y�8Ju���ᥔW	��!�g�D���0o�����rID�.>���͗gP%e\^����w��Ģ7��V�j��o�A<jaci~���=��Zˁ�|��@Z
`;w������2��Y�5R���'e��l��h��rmb鿫��c�r���z��Õ2�
>ѮTo0w��;�W��7�i������F��2�"7�7��y�|i��}a`bь�1$A3Z��f:�Cm�u0�)b����Uu 3�T@`���u�x���&�UT�븢�Os��	D����}y3���CB������5�-�����!���Uz�*���f��f�A�%|	�� ��.����+[�5��7ܲ&J���7>O�wsV�|� �*�a�C7��q8�P�^PR�Yy���!�����{��" X��i@��x;�{�s~�%�m�em0�Iw�X+�~1N=G�ۈtL\Y�i{-Wiģ��cV�R_Ła
n����
�E�YB�y�u��a=��j~q�L���z�#�������O�7�b�!���>���D��l��s�^EJ�������p���bF>��J�O�~��n�=�X���i&^־�%���'|��迯k�ylPQ�N���k����4(ӳ���</�f�|�C��t��ڍ�C�v�D0�HQ���W�>��ҧjw[��+]����^̤�Mz�}cU�����@�|���'���	�)���X3JF�A�Aj��ZW���ߎ�*�m��3�>�[d�"�ܿ�4�v�&����tǆ���X�1D"�<D��>@�j�>Ep��l�JU��K˚Yx��&��	���~�X	��:;��ٮ�Ѹ�|������ݡ*˶Ab,�IOFl��a������¼��n���V�� P�k��k1�d�IKͮ��/E'}��>������k�쌧���%贼������+e7L��G�G���-qD�[Hv6'�^"�j/����
rlpf:y�u������[mX
��{�0e�s�$��C�oeU8�1Y*�����"n�A�F�S]�Cn��`�z���D-Ӣ ���I�E�.�Z��[�h��l`��ː|��)��h�+�xhˎ\1Nؘ"��^)�#[�����͖h"-B�oe�W|��M��l��!��}W˪YZ��W�^��eP&��_��c
�A��rR��/����<� �7')h��\�I�}R�h'2��1�"�il�3}�j��+��S��k���%8�k6=O��4P/�jK�L ��.5��	�A�¡�4R]�1;�i���}{�/+�0���n�4��A�SA�W�efC^��I�k@��w�z��(�4����_��~�RN���N���*�T (R�By�6���譂�=?	>��^?�ʪS�O585�VtvBcd�1�P�%eS ܚ/��A%o�9�z6���7���!y��4٬a3�?:~�ˬa��2I��I��9�?7����P#�(C�b�<i_�F2ht��K��3�ѕ?c�-�4����]�vc�u�o�Ⱦ��rF�� �Ǵ����V��MJa�^S�R�,���;�}���e�
;�������n��u�+R�;��Lϋ�v \>���t����R�
5��!R�5���r"�p�/�9< 2X��1K;pWK!� 1p��3�.},�ٴ��r`Q�i
5-g/���'��'�����|ٕ6��'��_�j������n��ER��I��摲�}
�����K��H��G*N�/!��6��6
��WN����`+&� q=�h�0"���};1�o���i���(���[Z LG�b����N��f����݉2�M�G���wȔ���܁�&���<W�~t
�r���JM�LJg�}lA"�,��딢p�~e	p�C���]-��C$͒x�>QE�!g����?y�qN8��R	v�h�5�Q��� �nt5O�2P���N�Q��[]}��%"ZF�#~���ZlĊ����OU�Akם�������5���=տS�'K6���h-B����;(-��)J��%-f�5H���ߒ��v�oä�:R����� �;��&M�z�!f���q�3�_�g�5��Z�[e3�L���9��=V-��d�Ua�n�e���ȵ7����@x����4�G��@�6�O��hib|��/nڻ�{~s�)/r�+m���A��m�$ԟ��85bwEp�}�h���_��%#��l�*�P��y�3����(ֻ;��q�
��>MN'0��{Us�l�X�f_~���D��Z���FJ~��K #R����;�K��l��ڄ��ƚP7��AH��U��rĲ�nq.!�ʶ��Ս�h6�|2���9�P��?�|�5?
۶}o��p������l��~ɹY�1y9e���`�26bL�,L
�Rٜ̭�@f������B�������l���V�<xsR�!
	R{?M#&�+���8"`��K��7� �~����H�|��R6���ϖ��������NZ�!���f�ލ�/\ɰk4#�,ɘ$�{*MX���m����a,XG	wz�<��{���!��Tͻ��y������м>Z(��kO�f��u�_;X�ĉ�s��f��zj;v=�>Nm��pc������ �4�i��̉�_��5�rʊ�dpO�*�?%�iP���lWƁȎ�Q�X�;�@��e��7���Z�x�N��\��qű�y�X��a3�E)�S��5��'������0����D(��D�	�:��}��ib�y��8��+~׉��u�b4��2�����Qn%)�'~���
D	�6�ZM��ʋ_��N���
X�=O#��K(�DÍ��<a�����}O�Uӆ�|���2���-g��z>+��¡�Ol]N��( �땮��,����5c���#q�?m���.T�ΐ��%S�m���ַ��xJ�KgQ��C/h�IX���@Z�g����lPPOO4��eX���ٱ���K�����d�e���Y(*_}�M���zŝ�|K�'�W�bqT`��{����N����A���ċ�N�\+���Ŕ�Oԭ?T�U>�B|/�����;���\I����y����7�6$%�x�w�T#�!�^��Q�Ǩ5�t��A�P�Rl�� ���-`Y5��W
3���b�����@WU�s��O��]͔4��<
�+JN]��D�����N�L��A�Ѻ kc�2��*˧�Д�ǖ���.�.�~�`�������pkH��aW֫���Z6�}� w��ؤe�8�{��}��3:���LZm��
M�ֵ6:�G/�� �޸�߱�����R�s�g��$l9u�y�
4�M$�A�,F�ϟiF,d�RT�dC�.z'�0}�S�D����&��a�fC�����{�2�j�Րfה��x�v�YM�K%�l(���ʢ�$3|�n�����灹e|��ْ���<�!4����a�)V��K�)�ks��U)�SME��F��3���̳��a?PˢVzᴶnL�Fw�&qdd*��o��� �]Qs�)��R��O���Ap)��'ʀ�v'%�\l����8�S�����Z�B/���SW��7���Gkg8hK�m����U�9{o�3��y�љ?�H��kt�k��Y����iD5��_hb=�X�R�j�Du��K��a=5��o�X�����߸� �� Tr
��ֹ	ӊ�g�����a&\���EӚ}����%�yO8�
��l���W��Ɯ��lb����݁r�<���! ���ڲ����A�дT1���?�#N5;�S]�h���f�?�=5�KϞ��m�&xn��#����Q	zY�r<$�����Y�6�q�:��^,����b@q��[���Y�ɰ}"q�"����6m�`�^�k�WA-��+P�EI[�SE��cY߬֌U/�K�_�A�*a%_��i�i�Q��UœX?l��F�O����R�N N���y	�(,EPSY�TH*��A���$���d�w�s_qB��u�����n0���mU�������kJ�nj�-̿��Hp�~A]y����ȞߑX�1׸�l�9���D{�<vRגL'&.*����}�����I7Gq�X0�C�(�1�� �Uz�����\n�\N���ˋq��&װH��l���?%f�($�$���_,�m�\T>I��d)b+#|(��D���w�Ip����D0����WY��'Ԡ�C��'~Ƿ�n׬�H#�"��G���iI�vg�S4@�����j��5�HS 7�z�:4 ���2ofa9fV,�{du8����F-(0�/0�%y6:]\�p���0����*�c����~�2S��p���Qi$̐7��X؞�A���[t�v���Q/��6�­YW�k�V[��$�`+2���.�ہܜ�aW�V��a�%��4�M�!<T~��� wU�u��Y�b,���k?�7���eL[Ek3;�s������,����W��~�V�oz����7�3qm��`�9�Ej>Ι4���!����Dv@A/���]^��qr�+[�`�1}�\��l�c�g��q���f���`�Oi�S�������A��;�tQ~�^�9=qO,��t&�"�Z���F�md�Em�v���G�wI�F@�ٸ'A�� �}�_s�\�9���^G=����o^E>�X�BƇW �HG/E��j�qP���&AE�9p\�Z��@�����V�郈���a7A��d�K��9����f]�qP@�#-�Qy�u4Z�0n&'<m���;4�b\�O��K�' ���c��n�'�$��G��2py��a��f�| Ս㭋B�����(��{�51��b�?�K�o�����Yf�ɠj�~r3��k���nƒ���f���+���)�@��j��3��p�rX��7��%l��I/P-R���RRw�Mo뫦Ax��:��������Ԛ>a�tQ�̥�j�Ř����H����{�cE*�y�������H@���b��+��	��d�R?�/���CS�����J�qbC�4G���OF�{l�`���Fid鸂i_mD�(��_�r��,�K�*��������}���l�Z�C���`m���O4Q<�4C�Lk��8�_����E;ُ��ty�M�"���C�����X���Z�Q$�~�4"�6W>Rq��=��n�n��U����{I�TJ�6��<���d��B�|^�L����N�@J,By�s�Z*�NuK���#�?&]vnʉ�7�2'��^Iʿ�}�ʲ��/�h �̀�v�p� ��aB��-N�3�}0n^��լɣ���Z؋�pC7��P8N��n��#.zÌ/��xP?��1~��W�v�ga7�c�N�J���������s"������x��ZFu�k���rR�N�,�m�|����~� |gf���|���SZ]4Ct�̋�	 �-GS,�%��g��U��D�:eZ=
Ó�f 7Fݷ�E�%��_��a��*.��ң��橭�hO����0�[J�jה����lN�!������.���R�,O�����+�7�*�j�I���_�m�Ս��`7�r��s�T�`'cA���@n�)�ad"��;��Θ>ӿ���x2~�R.�����O�cX܋�X���[VK��/%��j4p(���<��H�>b��w&�G���$�+�EZ������F�ɒ���p_�T��/M�EJL�����ɷ�~�����,-w�f�R�+�K���v�NKۅ?7z0C#��6������b�Ǻ|q�/�V¤C��D��Ǹ����r��T���"���X��Ђ��h�pV�U%�9_�0���>���%���W\>ܚ_gO#�ܝ=��}��-ڏ>I�O#�c7����f*�oe��j8��R*����c�!ivJ���������X��O-���c�.O�¶ǅ����/�/�`-v[[��޶K�wa���Ca;����q�s�f���"�����h+���~I�7M�lᷦ3�y���
j�_&:Aa�t^z#e�!Kc�z81�������6��V�D�����&�MvS�9����G��q����S0���4� ˂� Hd��Ҥ���m�@t,yi#����VH|�$���V�~c���� 7�՚�)d��}v{U����YN���e�&�1�0�4���J��.Z��l�N��+�����IW*T{,�}����X��������P@�>�Z���=�D�`���EMab406�S���/��3$o̽03�>rfʓ���}Y�dcBMB��{f�ʁ�T�����y�����4�g�/];�Q��F*�P�������'���6{��N�p����\�~�H�EP;^�y��U���U���ou��)	|n�V�$�]z��_9��D�Pi�$u�̷�@�%�<a�?ǻ\��M���{��^��jK��L6}���UQD1�nV1V�JUVL7n��ƇK�NR@��l�<M�u�@F�-�N�%� ��9j�tR8r*X�U8��/c��Fd�D��Hq�3�4kRB'�AOc�Y���q�9�J:(��b2�=U?�?;}5�j�_�5qVn�g��������W�C�8h��e�@?�Lvqo�a,ی�9��؛2`^-�&�%@�~�7��ӹ�y�99�<�j��V��E���I�F.'��CB��d`��J=��(���թ��<���Q�S���!*NDLW ��lG7�&"Bw�F����|`�Ϯ7@ُy;.߆������"����-�m����b���`�)��:G�\剫����eQ�m^��hř�qo?��8�6���>=��DUqֻ$j��OZ�6��4��"5��rOxڣ�w��F/�����J����BE��!z/�cd�l�1�Lތ�� ��8�Y�(VV���w�)�wU\��QѾ*��ӁG�M�DB���X�F��*� �i��o�Q�m��A��,X@E��d��i�eW��$%�af�j���t��I�˨0��*���s�5X�bI���x����>w4?�[�2�q`�ٺ�:Ρj�)O�YHi{�D�`���
XY�Z����'	b;o֗� �
��2�M��E���Pr�>�sDa6�9�grM/����b�`�V�[�f��3�!�p�38k�b�:�k2cяC��1+��,�K�����E(]o�_m�O������$KX�vRq��#�Ԙ�-s�9?޸�ӷ�/�-����^������G�J���t��e)e���Z�v��e���-��	,�ba#����Ua#�h���w5��t$���QXVS强i�c-�<0:� �-�t\s�}���>3��YtB��NP�����UZ:��V1������;  ���R#�Ỵ�[����=�|��ʉ���X��[��6�c�oLi����DF��v-~1����P�XO�Ʌ���6���/�"Y�u��9�/�J�ۻ�I�\�Aw*e��⚮�j]�X��դ���)B����<)B_��8lf�����-b����Ƈ�B\���K���mFW3�螱꣹�j��ҲeCm��p��AU��b=�B	��^�K�-"��+�8^uN���E�Ķے8ǃ���m|��:_C��Uܵ��x~]\�\LO݀�<`��������$�_J������ �|"����U���^OKHj�/rv�����������1|����jG�{�D۱�.�	*�	{ĵ����Ղ��s��]�a�T(ir���f���L~�<0*}MA��bD���;m�斢���U�:�8q��%i(w���Ei1�[��0��RHDX�dsEy;���R�#���8G*�`�>��U�&w�����q�$	 ���?����V�J�9;tJ�S�;�$W��4��̮dH�Y�c|�t���$'$M�EJ��L���~)������}�3A^�#[�v�D�*��m��A�X�4$�;�/��??�F���X9��aʟ�(�o�=#"���������&�W.���F��d����ǘw��N��5+��##�C��T-%�eZ2cg�����w/�Gē�D���p*aN�r?���is������+¯�W�h�,���I��-s�C>��2����E�]��J���tdU.�/!����䆐��6�u������0�a�-�C���������L�����Uf��u�o�VRS5�O*1��) �;*�f3����f��,����0�>�`��&�u����D�4�u'^x����fwJՍA`G��_OQ�fR� �G��`�(�Yg���-'u�p�����m��mE��u-��͓] U�3(
v��]��F�\�u F$&)jC�W��)S
�����Rb�ō1wb���"����d���^.汷�˕~�������p����F���#i(G���'$9��b���6?���W�ZN&����`F���, ��M�sM��3�_4:zցN�Bc��*�J�m��md���>�09$]�w'!
#}8S�g?�Ojd#.��Z���o�ĉ�l+g�?4��L[����dw��R�&�'��Sst-x.05��~�:�P�{]��<ߧ����k(~w��2m��նPN<�YȘ��&�+�O��^8���5S1G	Z��)�wR$@x)M�6f�e�Cʼ(�&������WM$�a�J�ۄ�s���E;:�(ɳn�W?Eٳ���+H����2��3)#���(B���1�eOp��gT�*'�ǲ�dѴ�%�NS@�3xk��o0�7��iT�����5��+f�鐎�d�i[�i1��I!=Hx���A6��_t�}�h�ΨQ�����^��R^���9�=�@�/�D�vL�)]�;it���ȫ�yt*س�Ц��F`�Ll����0^ ~���&������.sZ΁�ȿ�D������P��t�_4$t�lv��������Rv1�HK�T�i�pb|�W���f��D�X��7Φ̩3B	7�@�C�*(�-���2��b��4 �B�
��[�&�i�K�@C|�r�Aӌ�rf-� ��|ٞ[ҍ���k~����?8�!�z#^�+��q��o�ݹu�GG�3X� �Z�dco�*�,+�fs�6.���.��#�j�uR��*�Wٞ�/t$h�y<4G)�I���+��H��t�>�V��-<�r��cK��Q%"&���#�i�oB�I�K�}&S����-�;t٨�S��S�&.���JiY���@�0����j�-��K�LkV���J��*�4P����1���`\q\���Lr>�!	���Ε�	_��+��Q� {�+�ҶrS��8�a_n�F���+VFH��|�e��q�����K+i����	��m8����:B��W)�Sx6��"�2�)��C���Nr�t~�c�,���%�I��l^����	u՗�,�pZ#�U�����]𳺅=@3��)h|�C)1�-P&%V_�E��-�Ƞ��bE�{	�k��L�! �6V�Cu��3������wxcPb��z�Y���8�Ī�3Yl�<!�$h�%^�3�L������Yܼ�.��%���Ni��?����X�~2\�q"	�yq���J���8X�?]ȫ/�҆��8@���$>�nh���R,[Oe�����auI�%!&m��e 4�?Vދ��aj-���m_{��̨�Q�u�N��Q�HL��S�))���w�!�}n�m՚�����4�y	����(�y��a�P���t��M��m��{u�9�-���j���FeaI��$���& ��&���!��&�Y��͹� �@~!����C��ӎF4գ�|ֶׄ72P�T#k3�m�P�z��d��+�"��Ey�}ӱ��6�0ݙ~�#��c~#7~Rr6�'�����-W��ލ.��ӫ�T�N^�珛�A��p�"��J/ᵣ�
N��� mMX���E���d�<�<jF���fs�׿�Aa���uj�*X�`�i\�K)�=}��76�����q+�@q��$)�yw����+x��]o��:;+��j^f���U��S�pJsoQ������l=uj�i��ix��`��`�L�E+�-��e����]�Sx�pwM�$V$`mXW�&˜A��h���� �W�1���kŞj���ꕨ:c�.��u�H�����V��Z��������T΁!���Opı�#���O��ۭ��;F�.?��<� C���ZQ������{�3_��>B�}$��	����2��Ҫ���jv�5� ��ڼ��5��\�K���s��F�ʽ^�DoN0y�d-&����i�&��� ��5ר	J�3UK/"����-&=�F�k խ���Hz��^#�Ҵ�?�/���fFt	Y?�f��&>��(�-;yG�C�1b߯p�T�Am��K�5�H��ɚr�x�ꌊ[�USw�M��༃L<�]���>
�ۑw���+~�݌#R*,���H�~�z/UP��]b%A���:�2�M�Y�~}�~�R�� p#�j�c�s~r,������&�w�8*����L�q������k�bYbj��]�IG&~l�����:y�#�O�����c�g���5u)IbЧ��b���삁�P���vν�X�Ί)�:~���Tu��qo>�����P	�Ɋ��wuպ� ��:��!}yN��\�_�����l�v�*�h~L���tq�H�PH:qe4Bk�E�e�T�$&���2~��g[-
R�z�&g2� ��C�S�����j[W�)hNXŻy���k��@�k�a~�]x����d�d`���[�
�Vs{G���S
���&4.`����崇|z.'�y�FC[�/�ŋ�˩g�v
\�,㜢��Vl�R�
1`΁�e�u�mՂ=�7O���a ���F����ȸCSyzue�3�^�̲���$���G��շ�E�x.�1�l���~��K4����{P�/l��0�r�^*d#irʢKr���-�J��Vʘ���#,�����]�[�dH/- )do���¼2��ش֎2מ>���/rGId�U#�!� �v��a�ۖ�.��
I��r^�0a��.s��a	|����@�jZ�0�V-�����w/`D�9
�WP�r���0���QPW���4������}�h��l|gtW��۶oV82L���#{
�$��(��$��'�B� 8m��x��j�7@��~���WQ���Q��~7��]��
����5��3%��,YHO�bm�3��\�ORkM3�ŋL�/'�]W/H��๤H�jb!�d?�]�稰���0�p3�<Ef���l�H�^�b'L���X�)Q� af���x��ۚ�h��ؐ
@��tqQ^]��5x�b�Û�i���`��S����G��u_��T���Q|�U]bT��L�%�z�e�k�j_��e��V�-mQiXM�vؐ��L�?�6گ��f�i$�KYo��N0��&vi�'���OG�,n�vx�%�pR�`�+��l���"��i��
r�IHs
�����f(fdWM�u��+߽��ٺ�_�>�.'O��3s���!]!	�*��	];Qٗ�~��3�K��j���4�8��(�
��=\�}���73~i&�f���n<���ɉ��&
�\� ��n����Yُ��>4_��;,My<=+��*����4v���\�TM��Ǐ+� ]�N%�PTK�? m���VгP�刵x����V�x%�^7���[b�+�������s�,���*��E�
y�pt�[ et�2BoA�O��S��)!5�jۢJM�|�R���\*.�VoE����׺�--��r�<�2o4+#��2�ն0=�Ʊф�+�/F\��b֝�����V{���!��q=