��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ���yY/���ԗ�8��@D��v"8��	`T��*�3�&,�_��h@ !�8,h���P֗��L,5��ٞ6D�(�ob��S �A*�F���"�Ϟ&O�^P<�!�|M�jO�S��v��a���Dsv����/�C)��B�~J:&����?|����k��U7�ot$Ъ�@�)@�$m�~R�ջ%&� �@���޶��om	G2�]BFW�}x���=�`n�/ڃ���q�`�{x��9>��bx�
�Q݂���:T�~�<@�.�2�>'�Ώ���ι����BӺ�i�
�nd�� �:��
>�0W�b&��[��w`65�]N!{��*	(5|���1E�ԇ�9�c+���+��FI�F�!<��M��C�o]����OZ/W[B�"T���_�VP��zc���� d��^�06��Q�t��Ob�gV(�njZ���UGd�ճ��t^\4d�mrp[8N�33�B!d��0m?VC���Z�X
��������_���`����s�*�ݾM�))g7������z����6���t�*���w#�.T�B�\���BJ�����i���p���lE}8� �00�f�].~c�a�g�K��;��ԁ����o#����.�\RM�Y;S!��D���ګ�"/S�C;���M��n�fS4��S��.�o<�~��S�,AP�o���ʆ2�e�8hR���g�G�/��w��l��&��M���n�����[:R��HQ�%8^�����k�T���w�Q6+m��� r�~!�oN���j�.b�QC��!څ�U��W��x��.|#e=��^<�CGNmDc��Dy	�+�%�=�)�(��e�&��1�y��P���F׾E܆XxGE�);(q]"�C������d���SE��6)��J)����'7��9
���W#}�5�-U���`W>
��G�frPe�E�X��ȹ�����cn��mY����p��rP�Rtg��1��,��j��Z�x���@c������0������;7�P#�ЦDT5��wTO���"�?����(i�eh�S�t��yB�V���_޺�C��N�f&�I+��ij,�s���Gb��M�+%DАv�����D�fZ���ڕNL��o����v����B�-Wޱ�x�B ������<8F�K �"9�H5q�o����l$���.�1&[OZ���	Hiׁ>���1A>��U���')��w-f�ݏ�;TF�����"&h��Z��܂-<�)�ozۘj����������?��S��g�]�c7{��ѽ�����j�{���5�^�D2&��2��0�bbg�c�>�'��(�4F]�N㺽(t\�c����Ċ�ݝ鰊�9!�H!6��@k��A߸:]+{[��fk�)���j�I,�s�o�j�j�;�d��4Ϣ%��D�vs �N����b���ť<�L��ֽf�
D�x�X�9�s�Ӭ��E��d0�x5`mC[�᝞�tY�F.G`�w�=Z�� �vڲ��8C\�i��R �j���eɡ}��� j�q&E�����M�������`��@�e+���aN���Ѥఄ%J(f��yM�����wi��M�ѹ�	�{#�.oa}η�D���z�	��m��7�l�����(F�`�-��{���+,u�5��ni㚏�w�q6K!�,��+�d�����i�"�ٯ�z�t�7�H��{�kJ�.����
�3��>�������Y�Ƚb�1�[��uܢ�8]
O�o��+J���M�yx�00f�a�
n�;���W�7dsF�p��sjT���-��p�p��2ۊ�5Y�Y���R�p �d�no�h�-&C��Rzt��\܋��QCw�taW�%-r��c����J#/V�S��M��}�D�f1U�����\��t� �0�=^�K1���!��;T�Ă��d����v�A��L5��c�~%�~C�h� ��ŠI�R7Fϥ*��L�-�(��;�Xڃ���c��~�~l�+�)M���eHB�=C#�~�+l�.�T����ݟCj���b{ �*j�8�$Nf8��R�TJW�ʏ�)V���n�b�3S�$]NїZuRI�.h+�˖լ,J(�����ʎ`ߖ{�p�w��}��
�=n7ᩬ�.���Ə��޲*�O��9��O��M�i:��	���f���9�@g���S���i�D�h#���'մ��:|�R��������d�L ]�H�[��nt:"�ˎ�6�U!J�~�|��x��F �bSLTv���L�D�9�+OB(�������Ͼ�i˥-p�ίs.?�R��1�j�BȚ�{2��)*�n+OV�J��M�lV8Ӿ>�ަ�ۀ���F&%��T���~CXպ�Bk\<���x�r�E<v�621��ʐEՊ�;�@��;D��Km �cu��p�Ǚ�j�L�U�H}��E~�q��+.3ô~�>? �o�<�Q��h��Q�GM9��5�����5nf�ɒ��yDl@���T5�O�*��嫡[l�%mÒTn�a���bvʛeq�:���I`���.�Ϩ��5%m]1����'^����َ��Q�i�޷�唟!�!�)�Ԥ��!58P|��G��aSJ�)- ��4)5�� �arܗ������l�MU��Ayh��?����$�h�%��̔��~�9�YlZ���c�Դ�	�������kˌW�*�������~�b�1V��gv���E*�i�*��o�[�u�r9��>�$�[Z'�"􎱻y%��Ѓ�9L�*��Bǌ�}F��՟�aZ��lAP�J�d$eY(n{�Gi���f }Մ8%1?C�X0MA�D�|���>6U�� o�yP����Qɐ6�D�K=ћ�Omם�LӘ�Sە�NG-d�х�����M��yl���+��e�r��@[��g��A�0�SAŴҫR��
�PsQv�4� c��%Cne>�c�-�����ȋV��k�c'O]�1�4�n����aȪ��P��7��d	�ת��R��Նݴ�o�l�>0���^�����	����U�`8�ʘ�m�NbUu�+�g�5kh��D�ïB���'�����>��%�=H��0ޭ�����ǃ����Ąr䢖H��\�Ri�35���
v=���Z�qe�=�C�^��'B���;:6ŃbCk��H���U��pԨ��S)w_����	����� \֬y>6ٜ���W�h'>�ig-�y���v޽����\)��J	�̐k�Qh0vw���*�� ���u���7(<'o���U!MA.F� 䎡?��d|�r��2�<W�ЮQy�6h*��y7�w9�∊M:k'�ʖ�
�l��D�il}�˹/i�V�d̢�]�RL�s�Ȋ��3�LQ<x6��6�F�g���pm7.�:�!�ܞ=t�͆=-����V2���1yH������_�4-r�2�Ϊ%�Zi�~n��Sٟ7UD���.��� 	�(�&�Ei�䕕V=����H��?�)�ҙ�r$�����8q)��f3�t��CK��뎶�f��-5�#�C��>=%C�.(v��=2���1��_�	�)�+g�+5Dc2L��<�o �ؠfN(�\,�*�.�vQvV\Ϫ�6a�c��Ȉ�m/�V���{�/���M�cn_��!;���������h���F։�A�-r��!c�ؙ͉���>u�3�ze���~�����m@\�L�H��EX��7y�`�����9�q�fU`�.{OMqZH�C#��FKp�fX{'d(R��
I�����c�R�j��)F��R �����-��
����KvS���ȇ�~]�K9�ɓ�F�SFU���G�����E;��YI�_{Fk�n�Xt�
O���憭.em�/@��E�:������=�I�l�����8Tz^:>i}�S�8 �n��J�L}(F�;���i�9j�� �E�[�1#h�@ʍ�aRμ.oEG�t8��e�:m��Y��x9tǅ���+��8%��*T&���G�<'�~]|M�04fX�XH:�*R�aeS���)/��U�P.�KQƛ���`T�����[�N1�
R_*����1�%���@�Τp&1/��,����d��5/v-�P�B4���/���6l�H�k�T�Ż&��R���<#�<�V������:��?�o�UВ�F8���cG�V!�O"aC���RyEk��)]�(��S>EG~�F�R�l��'�J�h�8���^{���E�l�x�&:�� �AǏ�qqJS��5�1�o?��q��`�Sb����4MH�g��ԑ�i_k����$�oG�
��$t���Y�U<Wo��}1S<:��6��<�o:g[�����Ȫ&�_X�OH�P�J�6W��H� �&��]u���u��ȍ��֗d�?0��C��Y=N�_�!t�k���u,.m-r��_9��t�a!�2���"����� �G�˺~,N"]�m@�cC�M���x��i�`l���2f�����*��a���3����V~���lR��$������}j�1��8��|�F�AAE�N-��1Q����~g_�C!�����{���G;C�P�hѾ�&����~�ʰ��WZ�ަ�#���Q����t��z߈[�|��-��g`�B�4�qy!y���I�0�!1N1̳�+�G)��YR�X�MDB(�%7DJ�h�ьZ-o��A�؛޽�ʤw a�-���
}��'ʉ��d�{v�V�9��tCp�p�x2*�d��3T�����|��ۭӱ��U&�9 <��E(Mp�j�_�T|�%��FvMҎ(�8�~Ԓ�����.�Wb��T߅���g�ɤV]3�t/R��?��O����G�&��Ճ0iFZ��׿��5�����5���j��/ֆ�;������G��X8<�ZƗ �X֢�Z�7S�'' {��⛗���˴+ ��T=�YΊ��Ȯ��k.��D�Xe���t� ����Ȏ)��n�\,��Q�q��dv��*���P6�El�Ξ�:'��<eq��]����Ç6�*�<_�Y?��8�C:�xX_Z�V{6?�Z3�@!}c	y��J�ۋeVp˦�(�V�}
vKTU�����.x�9�/�'WD�� :k$���=��0;��Orm���=K֩�������ԖҢ��l�����V�m0��'�$n��Z�L3}m'fP4w��2��a[m�/��3���mѺZ��D��+��E�4�3�|��N����!g�g�/\�����*��0�{���1�3ʭ>qׁw����i��*%�w=�f��ؒBOn�s��Jr���Q�*tq�c*)�C������Ɲ�8�S7 ���S/U\*q�Hh�[�:�ݘ��	*�R=�]*��H�B�¯�]q ��ܗ]�Jxe˛�	�%�k2~�9���ݱ轇&��?��lV&��<e�<B[jI-@LC�)������2Q͊{a�"�	-�/ıɦ!+�5�� (�e]���i?@�Lx�����,��q��I��'er��Y�*��7m�.�Z\qG4P�P02��}Q=#���VLfw�[��
Ǩr_���t�mȡ�/Ey��[�O2�U>�i�De;�.���d-@DAA���)pg��Mfq�)�
�X����1��M6῞Y�٦��|��i�_60�����74{U��&�''�^5����+�8�F���Nj]L�����
���*L;�����p�������k=�(�ERG�&_ۇ-=P�E@�8��,�4��k�+vm1p*����D������'CR��Q:N��*�` ��3B��L�}�\���N�;A���`�;^�o�3A'ar�?����I�)�{�E����Y'I{�9-,Zw�"0m{��O���|�Id$�~G!v9��/�����g�O��rV���t�fi�5�ސ]��+����_`à���M��ӷ�X���^�L%�k9Z3m����cy����)�E���me���2�[��梘PA��%��J1�6��n��SW�rk���ޛ�&��-L�F�G����¥TM�
�Y�8f�,���ȕ���I?v�6u���o�w�ݠJl����H:��3�S���"~���K�y�`�Bu7IҘv:1!ѩG�śZ�mdB�1��|�I����s��J�.�� D5b㲟i$pm�l���0��*���7�Sg��jv�c1tϣ)�vDhV��GK�I�~�2��6����Ui�?�}����J��kL��V����ırjk5u���5��v�%���.T��<�L����uG��c@����©�
����(�\{+mi̸���<OJ
8�L���gac.����W/��
6l�Z�VEs&�ye1��y�dn#�=�؝���y��W��B�iR��[�Z�H�'sx�P�4���_��$���ʇE�tzitbX4���e�\B프��!�w�8_U=�2�C�Ǐȁ3�oI��W��G�G49�\����4��I"_�Dߡ-�5Wd(�� S)�Ψ*f�ZlK@�Р�w�\,�B.�u�O�#���P�*��<j!e f�;@K��8�u���wm�>N;�mrW$�Շ'}�j��F��IY��,_<qD�C����yM�A� `�<�B<"5C��E�a֎t�K��|WW���Rͺ�[1Xs`Z�����9*�$������"ۡ�f��e�{���]~�ϔ�l�9��۶��F�R+m#x.g��Ñv0�>Շ��g GSj@̼�%mc�h�]�pD�mX��Nз��!���%zC�iQ/�� 7}	y��+� 8U���am���2���Lm�[�R���m69,]�2F�4�%%g�8�8!k��g6�|z�ȉ�2p��[�o
.O��=�b烇�����tҕA�b@���A�	eG�r����ՕC=G/��n�	��RL{�hTn�*����!���l0i���$d�z(�aF�G*��:9�GSN(N}ܗ]r8O��1��Cye..��O�}�<1u�4�#��Y�+/�k O�b$�^h� ��o|M��O�E�3�"t70aVJ4�aV�%bc��ț�=�x+����u��C�"JVY5�������̟n������n�8WI��Va��r�YAg�x��A�*u���${�oIR��m)p��s͕#v�s^�{����F��	:�mx��j��a�=���s$�C,���T����"e.���9WXI��ՖYS������`���$�]f;��i��g�F��G���0P�����޽��S�{ƪ�W}:/�海ֺ��ғ��dOID�*x[]��=��)P�i>�Ɋ���|��i�+3L*��Tj�,�s�m�&�+y���}�1�$�χ�Aި�B$qA�d[��b~����>��t�ޭ%�)H��Z��ҳe��Z�y2�g�,����~�-I�T<��� /m��:�w������h&"�h�*���N�����bq�i&�7�SC[|�2B�+E�}m*�IQmײ��ΰ���L������]1C×�����O�l�X�y�Hq!g2�������0� �[�ո����T:�͔�eə��4a�`�ɳ�U���Rb��2{��T
K@.: ��h���ǠLހ�������4N���_R'{l����ս���i=��i�2����
2`L'��¹�5����{�k��V����c�U	'���fx��I;���" 9Q�T��
�����Dڽ����U�'�%*���f��� Flu���g7�
�ټ�;߈�{�u�}[��nw��Z6��D��'M�RV��G4׽�J*U�-ڞb��� 
�C:^B*4q#hV�g�m�uL��������3�n\Ē}�8��!HU3�n��V�rȆ�^џƕ�r�>n��t긷���2�x������L�龿�q34�	i�I6r��u�>9��o/f� Jx��'�1׆[(&��Z�?�/ 2�ge���vv,(���{��T��#�
	�l��(���*�3��) ��~U��Lѷ�E���h`����w$�d�G�񛤈�/+�.}�����_1`#��~dP�7R����.��O�v6�^��Z���a���s�m�3[!�i�\�X����R9U� D`axZ���%���u�(m�TM���}��7�9�,��Vݰ�$���ؔ�����r��Xv[޲1� e���Q�Bm�&��Æ�½��#�Ѽ�уw�80g ,#+���zВ5x:��{w���+�<a3���0N�Ed6��`�*|�M��ݯL=�Cx`j�yK]�:
J����ZGW^c+� 7h��߂֠�G+UJ��^�De�}��>u\�.���H�jb����D%S�� ov�''�Wp��O��{����9de�b�.�m�M� ^�e��@�%�d@��>H�T�>m/�:�/�v�q��T���B����ܡo�~��\BG�S��:�=�.�[��h�-��UW����p��$�h�`C%
d� �\���\@�_4z�+fgx	�D<z��e< B,]泩�9�w:e3���3�t&�;0�-@�+�ˉ൦��n��H���	�S��j<�5���L�B�|��0T�Kׁ�r9Ib࿟��K��O�������4����xr�M���?}�W�C�r��.�����O���n��C��+������{�Oz6:Ú���wm;�<'����2�&+�v��l�6����������G�V����Ҝ\������qx�2�3���9.U�6b�8�%<X����R������H�L�yǸ���ļ\2�QT��}����W�����l��q��O�����:�k�52�Q��|� �����>���OO�ZZBj�B�#�KtZp�,N��{��S�4�+��{A�H9��Bf�-����F+q[��W��O$:-�\�5i���a��I�Y&�z��
k6��ABA��2+�)S�^"����loS}���NA�@��� �j^y�!���@ش����
:|��Y��z[Ny��vXa���m��?y���Kp9���+�@���9�Y�k}ț�񻾴�t6<2ׯ��4�<��D�7�h%��oBb4\r��,�fў:e'�&c��D�����Ϫ[&y�Έ��䏔��}�� H�B��ؽ`��7b�*g�Vfe(�W%�#��\�E��g���2�U���9�4Q��~m�u��k��#|oQ+�%�(�I�O��ܞu(\�<0U�0�*���w7�)m��P�䵹^���ܓ�v�[-e���3�>N跒BGϨ#�"�l^�Es��m��^Q�8z{C:�����z^ɯT�Ol�(�"��MrG5M���
����IU�����'׹�ڶt�+g�y���	{p7��ܰ�8��F���`������.����-6�[JE	&��Җ���=[2�H.���"G-�	�0�
%Kބ�wT�\��Sc^�\*��f�m>`��"�+�������|��Pj�77��f��8�5��H��<<E�����B�7���:D�KZ���ۦ�I�m��,�׹�6Ymr��ȯ	8j��M�J��`�ҧ�F	�^kN�����kw�A��m��mr��0�������9l§� 1DE��:p����\�(q$��	b󙖿�8<���ϡ��J��'</-�ṡ�0g�=O�闧�\T�
'�*~-$yA	���,���t8�D�IQK @}�B`�;����o��D�}X��ҧ��fJ�\��PZ���E�����tq�w�Z>��%�O�Q��G�q��<���fABB�bѿ0̊��~�6	i$6�.�_�+�m�̈́\����3A��=C`ît��R���b�i�C
���������G{�𕋑`siM��t�OF��73ڭ4M�t�V���-��c@^�	��$9M����됭�K������G4t��U��mvB��+z�ի�{�����'7��2_�sdƜ~�{��gg���4��O������Z�J�GF%qک�/�.��k�$Z̀y��U�"�7yuQ�ljG�'��H����b&(�t�O���m8���27�u��7Lܨ{م	�(�a�>�Ńr�Z9�'S?s'�K�~Qn���稌����?Z��g��|�]����":t� 9(�U:����.�`�,�@��0,Ff
��r�R�M���j#r��꿐��?;��]Ok��(�����#|��t��v������J� ��P;�be#�Ӂ�ώ<)��]LW�t�.9.E3	��4�R�I⢍�y�}��?�b�.�@cj4e�Ur��f�t� ��G��&�o3T�ӿ�(tms���!7MI�0����d��rΝȪx'�K�yID����IRye(�u�L����A��ϼ!��ʙ<��-*��
ݱw�"yx���Ơ�� �ϼ��|�FB��q���l.��c9�_�C�����KT���@�; �QKTjO�a.�U��m�-��X
T�:�C8�����.��D�	�q����u�'��II����۟"�F���^YF�֞G�:�I9�vc��]���X�cD����蔸����w��r�̉*��<x�4Ql�wb��*�"��]�f00>q>ѫ�T��JD��2����vD}�D2)��Q����S'����}�tܫ���%F��������1(o������{����m54�[�Jzf���|��g.�~�,%h���r��)ھk&��E�Y��ׅ��,̦�_��m�T�w���VL2Aҗ?@��~k����C����U�*��a�գ�9��?4Se��.��HNu��)�؆j�溃zq�7��*4wXGJ���>��zm.�U���������>���%�y9OM��'v���ΰ\R��`v�uX���egc�:x��i�Auny��ܽگ��(�o�sAt�(dbN�Q|�~�0|�՛p�d��?㣓��Q2������N�&��u�m��$�Q*���^�0�s��);3n> ;��]�GQ����3,3���/x��3m��_�I09�����36��v�:/#W-�6���jZ�|L[��N4)/�����=;~beLj[�J���`9�̭Ŋq����q-�|���!��ة�˔�,��H�n\�9R���h٨th���+BZn��~�^�R��e��O�a�iJ2�%pB��82�{�t.��|xC�0ܢ����z�rF�4�5��uB� �ۇa �9�����.�>�,�BW�S��V(�n�H,}��!8 /RM�aH^��fs���_9P74飜)�������3
G.�a&g��"�5��-f���{�bR��im|͟����܊X��'IwPڢՅ��=7̬<�b�ܫ�v�q��h��ЭؾC&C�aQ�"(8��S�_&^�LN�r�t`^���G�P�Jp�3�u��6#a�"�jOm�ATrΚ-����@�,���=W�y_O��dQ��CLH˛�*�߲�W�YF9�Av��/���F�Q_���Y�%�l�