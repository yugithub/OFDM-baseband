��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛQ���b��E}z&(^��]�E����nC�kaV)[A1�Q��ӗ���U��}�CR��d݌,o��,��?��4TB�)^������b�U�]�
�?BUhL�P?�r��f�ZpGY�����%�ݴ#��T�����𷮖Q�)�wȷ�AֿFhP��<HG
N�_}�H�]N{T�Q.���BC�5Iŧ;GG֖B�Ҭ��'Az6�͵M41l*9I���Z/Շߣy ��I���
Y�����3ot���S�=�/��K�-��qr�J'�U3�}9y�vT��[�o��9��ћ)\̑�/���}��w!�YO�3�j�7I|�|��+n����,�ě�!�����'�h�k\��oI��%H��'�(}��_����~�w'~�nzDc��|�7�c
�:���5�/�8�1lB� e��hG{Nr̭�/�x����i�q	X4�����B>�VK}E��S�HUꐞ�¢��(�c��
��8����c�X���ϣ�pߛ�čtj���K����&
dݞ!�����7�('h�?r`Y�.z�ɩ{��>�=NJc��x����(^V�ٜ�~�	м�����lphOp�&C�C����B��^!��Ue� �e�ɻ0\#��g�_]�9��?�/�,)�J��.�m8��������u'T��a��>�{3��#
|^ci}5��y�Z�S����>�*�4�T��zR���a�ߡ]>h�	��F0���4Z�j�_��e�,,�-�l�L!�f��n�����K��t�ٻ�-��� ��7�.�O�K���P��?��bO��@�Z����odT�!mh&)�2������>��5X8g�?�}b����U��x�G�A�EXs����ǣ�M�y���ia��:i��%�kO��c�혋�-q�A�KM7s��r^'�r�����!w�s#�� �C�K0�+�Dl ���y��Ϗ���WG,:B����=xJO��le~
J,��V(�����?���N��l-�,��(��m�q�6Xl{Vq2Բ�me��b&1��Vx��tjr��0�W��D�s�iÅ���q3]���a�x]�����C'���>Hkd�wZ��f���/����s��ë�T��}xy�G��SicCZ���9�Օc,`�h	�@A"�?{q��1'�yH���g���9Q:�S�? %q<�Y}϶�sj����)��	�z���t�p�ִ����I��Ђ[��]h���a�z�j�c@���5D:y �a�흘���ܾZ��'F���(^S�E�M,&w4{�e���4e�R�H������9�7�>*@-���a|r�l]@�a����zp{�?$����D��b�Zg�j��S��-Sn��1J���)�vSR�B��N�Akސ��#��Q�'��m��W �� �Cӱ���=	=39�¶=��Md�]�2���I�64�ˌ��U\Y����>O�gG��6'��=nwp�9ܼ��w�r�u�5m�jy��1	v�C��*�ȓ���o���tv%�^��3�Ǒύf#��(�7�|vC `{1G�OuE�2��m&l�ޗ,�y4���ڰn����$�\���ܩN0�&wف9
E>1�L Z+g���P�����xi&�O�
�ܾj!�V�S3�QU1=�Ӈ�Hz<�R�9�\����	x���\����cD�����t�<rY�m꺏`�ʎ���e���N��XP,l�z�����L��VJA~��:Dǈ�J8pg������Us?�^|��pcW�3aZwV�5߿z�
���qUtXz��=T���dk�����/����4�顊;���ȇT���_�Y�M�B�Z���fB<��Az��-�i����.b�BK���_�^��b�'6�Z}�YL
���7]я//]ԯ5��pcg�MU���wb���#�V�-(��g��,C55�w�\��;���g�h�rN�z筣=��S��Q�Bt��O��͈���Sc��0�����V��ar��a C��{�2�����A�`��ww���)}m踗#{mtg�k�ñ������G�\?`�5���Y���eD�EǶI�D�g�*T�h�wX4G���<h���z�а髍��}��㑽��2 ^�����e��o�޻Vf۵du���8l>����~
��0�b��ɶx��W�Y��w]�R'�K޷���MNȎ')�H܂ȸ5-����	5��w7J�aaٴK	��î\����~�2�+�G���;V�b:��7��O�}4�?0����<���ȑ*��XomtH�����������m%k`|�Q��{�8L#5��t�ю�oA���Y��o���bl2-35��7[��d���23���ݜ��Pώ 8�ߦ
;G�E�#�R6�v�9���ge>��ʇ�4^�Z����x�Z�zBK�n��+�Z����˔���<p��UI�o�L���RP `B�=�� @��TwR��~O��P~[g�b����YF���Jd�(�T�����X�#Smз���S�����(�Z�hIjŜ��p����iٺ|g��/qM	�ȶ'C�R{N�
�<F����[�lOfg�DM���ti���ۇ�om�7�l~4c�z�����@�V�?�Φ)Вk8��A�1����c[�i��徨Ć��-��bm,!9�;Am�ho���{?a�������W� =�x/-��|�op@ �B1+�ep �L�V]�b:���Ǽ��X���=��zӯ�+�
�?V�t��_�ԭ��	�^hݥ)8�����H���҇�ڤ};�5��c�P����e	�o�czD]�O� ��ă�0��*�f�kne��0T�
��w&\������Jv��5T(��
'�j��D��Sm� �f|O�$o�ĥ��f&��N�7�<[�2��pz���O�o��R�kn�^ K���fe��R����X�eA:H�iT���9�'�7���F{5��+fŨ|��TW��Gn3~ 8�ܨMa+L����QUĪ�=��1<F��W6���t�b�i
�+���/~��^Y�Q��[����d�?l݂�-�#��޹`�]�!6�֮�5.ƣc˶
S��y����l���t�H	��]���w��{;�z�;$�l+?!�E�t��BHL#u�^�y�ӫ�j��л>���l�����-�/r+�;à{ч�A������:�"�w�^�x�[b�KN*�VCF�:��m0��C�w��3Jҙ�T��Cz�ԥ��F~Ӄ�g�G0�.y�2�JGE���~�ɹ��D�q�ߩ���pNȯ�����h/�x�p/C�&/	BŨ�s�84�/xH�(K��+hJ_�pY� Z�Ȉ��\Y�ȫk(0�-śzSr̺���������ڡ.|:T(`|�Blc���{��ƾ*;��R��ͬ�`|��:ҩ<��)�ͼ���T�����VV��Q���\~��M_�֕��R�6Z(��n��o\h����D�w��::�CgT��R�΍��;.�A���ځXf��^��M?qk���t�V�k-q*HLH!n��Ebe�r�b��m�սyVa1�T�;���6h2�r�vU�����dm,ºj�Q���#4n��5�"��O�B-����}r�����n���4?&��X��(����|'n����󙇰 &fC<���0j���������|�`�W���?��\xA��z̧'���������i��:b�v��g}zZay���<߀\
���X�.�gGф����{D�i��~l&<�8"�!��B/Ȋ�[����6��Tc�V�n\��'��N>l���D/�-� ����3��ٝ�B�H��M�Lck`�G`��x���a�w&h�az�-��яx�)
����CV�,)�&���8!�����_�-B�vm�=��-�u�\��=m>��h-I4����3���/p�Y��4ҽ��2�$0\�_E/�#������ƭ9UV_���Q�.&�K����z���hLQD�ʦ3B(A5U=�����>���T����j�,E�u��Ae�(�5�B���� �yO�|�Mq�B��Qo����m���7�@>�ʠ���'V��6�*6�Z+N���䍜iE�y�	����ndqw�k�w��Ԧ�7��o�S��
?Z4��Dt�}���9��c��E��Q�����+�A�A�7�YE~[����d�~��ea(�Ȑ���k�IZ�e$2��lT6�i����4�_������@y�ȹ[�E�e��w�����RT?1/��?Ǫm�&]�jJ�pI��2dS/�ή7ZKʿ�׍^�_\�E32J��.��� �FQ�;�����&n�<�e�M:;��ֳѺ[�t�E]�ܜ��@��23���a|��G�����9	�z��yљPz���uo7�����Fxwr��n��=[�0���"P�����w�]?j����j�
����~l���RaO�>Z��-Έ\f�F���a��i9�����w�F�~��V	�(O�B�>l�{�@g�XK�	|M@�HS��R����~8�C� �ڠ=ړf�[�,�~ã*��`ú��Nlg���*��x�B�U�P%��Wr�K2]/�;�{'1-��۱� D�)v�w� ,#I ��������1�co�ҧ#� )��
i,��b���e���~�j_Ma�A��d�g�КH�G�c�2�d��Oܳ�0R��E�%�q]Vd�w6�BC��A.Ǝ�m=��:!�ΐ��ip�P}�k�z�Q�&sn~��4������A�&s�����Y[;i��P��[�� �R��g8�sU���W���L�a>�
�D1d�r^�����{�62J�.�i��u�.��S)���7]�Ɲ��ۿLQ�J@vn���+�����Q��!*�t��ػ�"�x6�Y6ņ]�\q]T�^�gi36�r��9,_ߚ�Ys�D�>*�S1gi�;M=N?AY"-�?7�ʣ�K�<�2��Z=�V�g��i0�`vu��I�Oo������qH�����,�����? �\rh�l�M�$�s|h>����Q#�?%sO0;Z�ع*�a`�G�(��.�S\.��I�/��5�P���N���p����ь2�t��G��Co&�X>v��ʰ�]ۡ�2���sz5��6M��z�����9�=K�[-�}�3���LZi%�/f1��b���G�Z�>��g��Y�a�J�� ]��*��f��EftT�;SH�|�h��}��t(�x)ǆ��r��X濷��<-����R,q�e�����X�
�{l��w�Η2I@U[��=��G(��v�n W������~�<I6�&�{�62&"I`fQ�"��A[ws�����rk�f����z����yAG9r
߀"�O�G� ��w*'`�k¦pe��n���D,�����nRp�T ^�Rދ��+�8d�����:�6�ˁ5F>���@5٬`]�YM��$��W��+�H�����ő��! G��jCV���=	�>�i(�����:>A��s}����l���%ZV�+Q��;��L���Z��=g'h�Nkn ���%4�122����J����ufꨶyM���N="���ڪ�n?hxl���[�y�a놊��:�I/� �D9�J�'���C�x�EI	�6���iZ���/�xUǾ�D���GhD�� 3���x!p�2&4�R�ܹ٫���=��Ŵ)ڤ�j����㳧qW%,x	s��&'��m�����@=l���XΙ�@��C3x�w).9�Z(��q$3�NA �6G��wN/�
a��i�S��B[tU��۲��/ڣ{n���W��]�E���=�7���+/ܲ����4.Q{rJ
a�hr��$+��T�m��>��p�����RroWȳ�����^�9��C����!+���!�ԯ�T����ݔϨ�\G�x����