��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛlb~�mʇG��CY0�p��u�������-?�17�A��07.R��P�37Jl$�a�̞�)��x��G��P
]H{�_�U���}������,4~i��z�˧��A&��1'�<�ϓW�>wY(~|�6S��ޖ�.�̡�oq	ݻ�*U���\��'kI�>了[�.g�'��gۼ����I�|��8��?�������<{�ږpC��{R�[N|O�E����(��%��l���VSҡ�b��I��L���wp:��8�V��t�H�$��@�mB����T۬����X�`\��@vG��+�q�_��Y��Z�6V`s,W�C��^�%:�_���PDTYɷ��kvq,��aIٳ9
��M�����v.����wF���ȋ�;zr����:M�#�c_����ҁ���IH�j�pٳt6���11>�vp�a��<���p�������&�\���"Օ�RMo�y�h�($l1��F
�?�01�{��9$��Y�Z����蒟��#���X�e��aY^'�/[&A��Γ������+�bӶ�s�?}��}ח��}�m��:�&u���Fp�tQ����6Vl��x����+&�f� ��My7޾ju�h�x�O%I��nfr��Sc%N-p��J�}��0���y���B<��3?�f��F���)�n[�آ����~3�mU��mpB��5HјT�޾�z8��-�E�a��m��~��� ���arI�Ũ�H�����M��-�!���d�V�`���RjR�3u�>�j���A���C�1��]MY7"Y���3^)��j cx�%c�B�_1�BI��Ր6˞�Ǒ�%9J�u5X8�X�0)əKn
{E�Ζ�|@��UDp�U��=��[������,����Ȋ��1��G��t��ݸ^�,wjR���|��7�Jύ,���&ƫ��è�%	2ҽҀGc��:^�l�a�cd$�.E�2�^��V?)����C47��I�o�W�E!�50Ӛ��~�_H�t���=�1cbPn�w_"��\�9�j��f�l�AZɀ<Hwܦ?Ź��`c���)�X�,<?Xɛ�S�F ��Ub@�b�XC)�H�!?e���B��hv��6q�gw��V��B��R���=m����r�X�q�fi�C�j�*}����+R(g1ǃ$wXp㾝�йB]w�8���]oc�J��%Ąt��յ4SjJໟI<�z�O;AAl�s�l��f9n�ȇ�?H�o�����,S�kO3��&&�O�R��Q�Z��6,%�nH���3�<���`���~m�	:�4�I�#���Q�#'c'Lj���+6$Ng��;� &풇�VV��=
[+�$brd�Y7�`n��+�;!��ٱ�4�_�v��c��HAb���&�"��8a��Uߵ M��OF�x�]�&`��*˕��^vh�S5�t�Ѐ�Y�*�Y�q���{%M��9�L��l�1��&������ ���U#$yd�N�
+���0�$J�g�d���v������7��Q��
cז��2��(%[dY�%��&�R+��M�=@�����CS�At��� ��L��l�u(�p�y/_�&`^�����h~�-x�Sm��Z�������4��G�c̫��L�'\�ps��b9�Cʷ7�2_C;�OT�Œ"a
';n��2F�xk�p��D��0k���QsҌ|l�� e��	���`�i��M>b���F�\��kר�mm��[���곹�##i�������d2�MG��)�Zj�::�D1�e#{ �������*�.���U1��W��adS�Zܸ)/e�X���S���BC���Sg_�c��b�e��e���0-(G݈��qN�� �����(��v��BX��S��K�˵DR���2jIE��D�iu*]Q����Ѩ�t��6@
���vP���)S�tF�ؒ�¥$�iT��٧��[����
\��\/�T��-���,n+ڣ4ΉȗO�Fsq+������s�D.c�ma]�y�ӃC/�� ��<��kV�^��'r! �>��4 -���[�I�@��{�3[�ƈָ�7 ���GN�%��a>������\�����L�B[L��j�9{�a�"�&\����E!�x!C:�Ւ�;(�J	�X��5Q߬NU��D\���P��%��v���1�ǽ[���P%gOgZ�}���v!��6��fi�)t�ʞe�.��V��4�e�~��j�����}�|����A�?�A�l�
���^>�Y�"أeg�Ω�+4��F*�^6��fd��v�����`I�k�S�Ȋ�We�%��	�E8�_;�e���	� �N ��W�l�^6��0�f)��W��6�ʺ>3���ȅ�6g���~�i��I�pD�

҂�"��{#Z�N᝝W�jI�9W	L_e�Z6Lsy�EM�u��Ա:x���B�����.5�!�͏U���U�Ʈ]Z�=�s���!�����h�+:g���W�W���C+I�Q|�,��c 9��*�w*|4軤�6x- �|:���=o���ގ�'�,тݬ��V�.�4y+x�j�
8[�,֗�^
��H�#�5b0X:�'��$�o�#���N���`]5*�A'����&mQ�����Y"��x�_?n2��fʊ�����0�y�/4�_l�4��˹ź�X�w���F�z5�����MX��?��jM�p0��`N��H  c�-�`8}Z�t�	���g�d���I���g��^�p6&�����]�tG���(���V �Ġ3J�2D�����>IQ5�m:P���g���k��୛��
 ��sF����Jl�z
�ϕ�yݦ�o�Z?�jb����*��k����P	�׬}��R�X	�t���A�W{ö�1�L��B������y��y�/�B������RB�gJo�nv�� �ж� �?M%=�L&\�UY�K�^�W�".���mܼ�.�C�n&y��ojI�X/�:���e>�t�Q��~ Cm;���e�5�Ϙ�D���R��t2��4� ��e�C�k���B-���T엵����2z�������L��>��]Yd����e�<$�{f�*p>���,pX�{�u��L�pG�!Υ�OT�?"% A�px0�p'�'���2tme����"g^$�
�#E����{@�5�YCY,��ư4N�g�0G��8=C�
�R��9��'ά]�l��I�R�?n���MMA+��/�ADǢ�o����T;�&Zg�V)�>̥�C#�Ӣ t�V�%X����y�$2i��^�m3)d�b<M{��d���8�H~Ev�JV�=)f/�95���N_;�������[�&�8��c)����[k��8����T��<*(�b�	��NLM<OkN��
]�"HRPd���-�Gh��<�d[���[0R���i'�%�2ɠ��Sح�N��=��H5�$$b��>�Qa�gpd�3�ݠ�v�XM+��<$
a��ZbW�Z8�;<�4��=>�so��|��5DM��>Y-�~0�ۻ��1��=
�4lW�G�� �2b�����^����D�r��e���_��&�f"ۥ���%<�S�,��+BrG�o�̏<A(8�Re_��(� �.�������f?}(ϴ	9I��s�y���n{�A}+��lb���i�f����%�?E(��ķ�>����ع^��5C�@B���c��k���� ���M�~�MH�4�>תQ�ҫ���;!�z��V&֖�G��-�ܢٝp9����́D�CQM�m��J_-aGn~���F�*Tە�An&��_-�K0��RZ?ZP��t.l7��,r���c�/��ԣ���G��APQ�@���4S[����ǌ�2��4#�ݤ�Ţ��Ƃl	j��a �i �9�x��C�.��O�(��jX<S�o� �g�.A���G�gB��`��ʶǼ�Y�A����z�5)S�
+�@�5�����tt>�b*�����b�@�s�O{�f��H;�b����w�R�V�p����=-=��v������p����#���xAp�&�:���$	!�9R�����iY�����r/�� γ%�
x<�_a�	Z�^�,��?�p%@TwK��C�~g�Q!	}Ow +��Q��䐓P�ct����3��ѡg06m������֏%g9P�Ku�h�Vd�;�Lt�Z������z&U&��VU/ZW�[�o��ot�}0^ȡ�F�c��l�̶��2�|���XFB�m��{��{�w�1��{=E���!E��`OZ`A�ժYƐ���t�����mM�j�voN��[[��L���@k�8���C�ꗮvc���u��3���`�B� %-5&(�+�7?.�;�x8kJ�]�2����2�?����d��Ё� �������)�7��,�1
wz��v�~��ж���>�V�%���i����m�<���{.�ϊ�C��N3}�r�'=�X=k|��U����l���zū/��H:���Q��ɧS[��.����fv��'��_va�:#�ċ5*S���/[D3�y�#X#B�����T]��'H��,�|O��^T����ɯsuq�a6+��c~D;�C���o}���*+	����Dq�Pl	:ہ�R2���]\ٳ�E���3<�UW�<��j�`�bw��[�9�T��4�����,���we����
�!+\H7��p��~�f��5��{Y���(rg��}��#(�t�V-��Z�8�C�CM�)
���S]�Q�-��	8M9�969�3�){�h���Wŉ��H�ܮ��åPYhwe����;����#ė�f}��Y%�rB�3��5C���ʅ�n��c! κ�j��8b" 2�V}���a%�-��!4*�թ�,���Q^ F��gF�fF������2k9q���X�\���G��f��a�ַ���Vq8<��թ��]W�然1Hm�����YkS�s>0*����:�H�ou���	���ڰ�v��o�S�F�h]0�mkJ���]�Q~�ρY�p�p��u�erU	��<�I��#��x�DV�X�E��D�'&�<Ѩ4�v�%�)�+�=�s�ԎJ�H(��حL���&Y�]��[�E7�$2	Ƅ�/U�Ӥgy��޶ƻ��V��� H��o���j��'&�ꝲ>N�:1�Q7_�|lP�3��? �#�/+��O�%����stۀ\JD>;p]�H��A2ye�m��1J��_���O�m@�-A0�U�Y�9ff=|\ԬM="͛��͹�*�wBr�=2~�*hh�D$�K�ś��IS��a��y$AD��ҡ=�O���*89�z���5X�?�s�o�Q슥W4���4><X�i	��Ɗ6.H�)�/t�����n8�\�"%�����d}[��=�� X͘Lz�l�N=�(m�0�D]{e����X6�i�|P͢��	(��!

�~��Ж��G���|␚��q��#Q��L(�����ƶ.B�w��������W��12|��@S�Ϙ��=5�o�j��q~�2����1#�>[�����θ!�$W!��I���X[�M#�_Ţ�`W�vK.W$e�'��@S�7�M�].������ >D^����_yh�]��r���i���ݷ�MIG7���^�j�.�[�`P�:��C���/��7�X$!���Ǎ��mD����G�v<�Tw��b��XtG
��Sڨ���H+�[��A�ρ�����Sz*'UmI�N>�6���9����:���a�ʉ��](�9���hds�$��� ��1�n��r�Y��:Ke��Ϊ�K�q�p�d���|�Y�n J��-�q����p��xQz=PB�g(&5��ɕ]H���
\#2}�=7�K������l��{!��A�uQ&���fUq��
Ht܏����̣�:�ٍ��~��%��Z�u��`�]x��:�Ν	���tJ�,Ip��i�	g�����~�W?��O��#�)�T'��x(�����ӣY�������*|#�	��+� �1���f��Qv��lq�%��& s �t��҂凖T�� .W>,H�\a�!F���Sx67�hĕ�G3 ��3]�����`�����5�
(D����rH3�P2�{���p�+��kjy*]sh��Q�*ݢU�����)+W�3���d�juB�XK^+���K�޷f	hJ�Ǻ'> <�UBV�!v6z�s�4A稅,�6�S�Q�g��@q��V:�-����:��v���Ǩ[ުL�U�%�bS�>خ<��/~jv^ڭ�6�I�eJ��d�Y�0��9c�xT�dQD�CY����2b7�΁>>�U��R{�rvܷ�8f�3����#$Tn�*쥰��Q~�y����1.�7�����-�x���	��1���w�q�rɉ`���>I	�Dّ��&I1�LᬀJT��j���aUo�>��Kʝ�q����9�W�� ��I.������w��su"D��N�C��i;��]���%��s�J� 1��Ω-Ti�R�����J�t�����`jƟ�wG���#��������r!nc���l9�L��������]��['�V���e���\�U	���Ҥ�x�V�Eq4w�/�tb�t>��pQ���ޏO��f:IVZ�* ��M6������Ss��P:M��.h��T��C����, �� '~6
����!a�TD�q|��[Λ �*ڢ�h�w7�F��:�	o$�F���t�Ox���y�a_�-��y���e;O{��6	0���fn�k!��'�/��t�	V�l3�z:�{Ԯ"V���`5b��av���7S%U:����*�{���0�u,�	��LCC���z>�k�:(B[�Tl�Qs�d�F�Oȵ���DO'.7���)S��"�P��P� ��*Ǻ�RDO���9w��9'-Д�Cx�EK�,�����x�uy�U���Qt��^�
�Y\�%f7�(6?]��J�!�Y�`���nٗgc���Y�i�5Cƃeh���M�	W�8���@LcfdED%�BE��b���j
������nzg*u��+�����GPŝg��e�4-�78���`��;���/�.�����S��[�a��ÿ�jF�h7� 
w���n[g��*���*�A��}v��u�$� ��N0SAw�fΌߵ���0'������Oe��LH�aBq2`��.4�N����������	����K,��!r��텫d�OYe(<��a�h:C�����g����(*3&%�3�������`|o�u���QNR�����;<�`n/�H������[N����k+2G_�[r����x����v�b�G�,���7��-�M�M�x|? P2ɒb�-Am��uaU�I��{&����I[��D�5��Kŭd��SU~E�gB?Ȥ�!���)0P��3��ռQ��Γj�bIX�%�Zj� ��f"���O���h<Y�4O~�Ǡ�90["�]&�7<֨y�R^NR���}!2�1��d�48�r�Lz9�}n�ꈻ3c?�_�bb�����1�!��Pm���ɠ4L�K�.�r���.��> ˳t�1�3����v���F٢v���+��-E�@8�ɝ)TJ��*�Q�(	���|�Y�*"����w�J��y�]��ڶ�,%,%�@9�(8�� �J:�Ky!��{j0���*��W#��(A�Ҋ*�6ݘPThd���|���ܛ�Ɠ^�*C2|�v�؀�u�}�vp��?�U# S��kO�ε�C�F��Ik��l�KRO�0��Y����2�e��� ��8_�+ԣ�3L6�̱x�Il�Cp�_�`:"�?�ziϵ1[�-f.���*pf&4���2��X��<Ui�5�?@�g�$�9Ă��V�ۯ��$Y��4_�yT�j[��Z�RM����n�N��$�LQ��y��dr��������[�C!-�&V���e��Oka52G�K�mB",X�7��%�R0\��I.�3:]�*�nD�	BT�T�����Ӂ��-��=����h��#�_�kgP��"[��@&"�1�n�1i�梡b31&}.3} ��z�>vƽ�0n�9n?�� R#Ԝ�D7����T��L6�;�C7u�W��d���{i^�C-�(lb�ǹg!fV��� ����>	'R����̬���Y��Qzb��2;_����2��9Qp2�t��s|*P�( l����v�iZQz6ř��V`��a�urAv��d�g���Ge�/{v���������������I��0W�3�[��6-��~�{��#ߌH��K�h}�=aJ�'�9LJ�y"D��M˦u��9�ו��Q�-���R��}a�z9�Ǽif����Ua+ē�r��}G��w��tp�D��s�θ���dF�N���җghl]*^�K���d7��ֳ%��|l�%�4͘I5�r%�gO#��@z�K��y�]
dC��nP��,(��1m�fb�#�I>��z���oP�H�� 8~���*Y�j�Oֿ7���jY��w��{�}gj8��-�B�0j��+����o5iFO���1T+Da��~ۀ�`�>8�ݍ��Q�oV�5��4��ä2v��]b��mw���\֟�"U��@+,��iЙ�ˢ���<)�hʅ��}Ή d�W�1zr[x%���������D�:�3�����_ٱd��u漐'y�1��l�����w7&  m�Y���&���/�.�SlL�[3�?���R��9�$����D���	_���L�I���o��s����K$�s���EtW���U%/@C�O�Zz4�| �]�HU2�:t�tap�υ	ġ����S�j믋WRF�O�����4?�d	ɴ��)q���uY��!w̴��F�jsMs�͸�W�b�K+~(WVqe*���#�b�ct1C�R�AqѪ���f2з`��.	�V�Z��l&���N�gO����>Đ�>�X�5@��A�6��N��C���(�D#��i�9¿1w������$�kMI��h�bWX݃�^�����w�d{��
6%�������{ 3�_%��()Xt�!���Y��p���D&���)��5�{�E��#�Hֈ�u�o��D,mk��*�\���Ɲ�.I�&	���@�"�Q��&�r�Wz��CT�����s83�OU��.����g��-���K�w+��}|sJz�p��#��R��gr,)�8ɇ�*�A�l]?��!�g޼w��'ê_��'g���	n�Ც֐ ��5��F Ur&`Z�*d���o]��G�9P�����8�CG)K�K��%��~L�۫�jf�Jv\��	G�01���8<8[iʊ�ۖY��̇$���KƗ�E�Ͷ5W'G_���M��ޖ����0'L�j�`���4[UP�ݔ�����ʌ���05I����a�_L���h[��ws=q�����*�;"��C��ye����uS�w�[���}:���kE7	5������B�
0�-��V�$o�Jr�zI�o ]WN[B��b�&��ä�۰��t��s�S:+ͮU�����H�"tq�"�Z�z:�<s�d�B�_1��=��s��@�x���b�+<ݥ�	3Q�dG>�|���t�����1�(��8��q�$����}gL�r��a��$tIg���T����J:Ѩɟ��-zchϟ+�eb6����tYd`z�0��)�`����[�g=�/6G@c�ˤw�r�)��Ɣ��������v8Yͭ!�bI�0�Q)<I���S���2Q҅Vy� �|��gIB������ѿ� ��`�p�!�"s�}���e�k�&.�z���$� *�!�k��8����Z��s��J�r��P)�A���Is��ٷTν��2ji�͑.
\#�(�I�����%ʁ��fbrZ�1mz7��/rRX��;�HQq?1���_�k\�W�C~��,��<�n�>�l���*"�ff������W6��_�gT�WF_r�Y�q���^^x+� �}Gｚ��C<x���#lwYuh��ꁡBm���@cK�%o��$�	[lm�[l����~E\�Sw4ҋD�Ϟ@�s�[RuH���n��Gd\}��ngn8��� ���4&5g���q�7�a,�ҫ�SY��U�Acl�G$���z3z���Y�7A z����+ɛa�q̀T�Р&,PQn���]�d�0",_����d�/B�+*�"Zp���P,4f�d������k*5YwT^��̡���_��U�y����K��yK|���A��Q��A�b���K�o����0�>��w|~�!��r���LV��;�J؞�T�="j�R	�M�|�'���B� C���>��Duw�[R�����9�&3,a��Twh��5/�j�:1�8���`�b�g��}��19��߅]���7�4K�I��F���F�����t��R�$m�'3��{�`v\\���r�^B �?m����� �k�ӎydϡO)���u�_�@����T�K	P��y�V '�@���ĕZ^���0��.��-��3=�����y�c����ӿE{���
��R��4#@�dd��ye<25��5X��jJkT$�+D\"d�bj�>���יa��iԘe4ڂC�FE��U�+�q�5M�n,Ɣ������[���l�"���p�+�$�B��������VD�4�A��������:�K��˶`98/J(b+����.�Ɣ�:K]��"�M���n��YvK�&���<KqZX�A9�c#d
3�*�ؼN;T3��ܳ��ş�V��X�R֎`��:#��(��D�I�?�=��^^	��T���~	��H�
�������*spMv�w>�}�N?q�4�ϋ�L�A�ϼ3�gy�˶��cv!/:�vZ����]�9$�h���m$pr�D�Y�%�x}�	$��o�]�+���'Z�F���[��#�-��Z
�YEʚ�j��3����]8g�P7?��F/&��<DjY��]	�"Xx���늪�K)�;�N�Qk�����Zf�r=f��e�,�vGж�#=1v>�#~�M����l��4=��}--����_
n����AX�d�vc��T���rȊL��8��A�c�d��N]�&ˍ�UU3�U���iu{�gʫ�P�I�9�*��!�'	z��Uї��QT��.FOX��ص�6z�e}9�Q�5�����}�p8=�;�/��-�3�Q�;�f5��B.��nַ��{>���'Qc�3�e�V
#�!>T��LN�4]0�&;+w��H��JY����_MݟxX���|t�'���ئ�=�竀��Z-/�8�y��F����łJ��jHt<V�;4H�g��: �&�F仒�-pR95�gK��ް��^ސ'����Ih-�\��B��H��\����V�PT��s*P��{=lF�V�;z�	^
w��x��P4X؆�0F��%��^�Yxc")����T5����'��s�I��:6d61��Hn����Q���=���н��<���&KI�V&y�!M-�"�����A��U�^m�k�"�&珯9�+d�
/��2j�&��*+�#KU26��*����w�<�iw��Ia�5t�z~ǔw�d�]\uJV�ZnF�ꭷ�=��Z\I����)$��z�&[�M�����u<�6t�?�'��z�w���wݯ�1��w��������@7ه�Vsxd�ʉ���Xe�r?�
���p	C������`lp�OSS/:�+�Z0|��� /�A-���^s��g�T�6��J�̰ �h~r1ca�ӛF�Me���N�`O�m ������e$I���p_�<�2Ͽy�T�4����|���	Uh�&����!cArb��/>�@��&|��ȓ*-��܀h�3ƨMJ��MP����М�_�,ۏc�/�ing��P���W�U�N��fZ����򑔉��虻Zut���;{[ʔ{�:l�%���+�ܲ���a�Y^�{�<ΏƇ��]����t�-��8���2��L�)���i��Ze��@��z~�����4��ob|��FseH#Ҁ�adS&��ddݜ�6�q,gЋ�K��!כ�=eC�P���0:�X�t�a/@��
>���=d(�#�=n�Rd%
�~�}��S9�����)x1)�lw[�~[
P�M(IH��M`ǰ[�W��*����* m�f�?�;#�vZ��1��������A2Q���7����R2�$=��.����!w�^8h
�AB.��D� z��&�7������	���vkUL�?����8����z���=�-v�HrI`Y��4z{�@@��wm r@0Vx��D0Ew2:�h�x�W�ND�*���@F܇�0�q#%(O�1=*�� ��ʛ�:�z`�=Lb��{����si�����㙳�,�U/���WG�������O��v}������K��Tx��d��ɴ�W�G�;�3*����WΣ���*BLW�����_1�q��p��9w(��0ڞZ��W���հ1�
Dt�[�8���<0dR���!e�\�~O[�� t�M_��M��|RTY�=0o����?Kj�s�\dS����Ǔ�B5��3�S�z�x=0�H5� �>���QYlmU�ɰu����G�׻7]�X�`��������2C)���x�lnN/�4�:�(4c���Ch�}���uH�_At;ONZES����	� ��S*��M"�������3=�}`��[�m�r�Xۧ��Btu1�;������{��z9�~���&k����l�L��&��:Z����@&s�!���~S��`���8ke��E�
߬�	A_�a�s�V�����)�Q�������9s�l%���J!^\���V��Eȓ���4�n6����byF[u��xk=.w�#�@��vs�lk�M�Z�\R��`���9�c��Θ`Ir�Y��8��ؾ�.ӹ漋�m�JwC�7�&�U���DC�ɾ���O��K�%�Ct�#V��v���DA�z|�֗�I�x>�[�t�Z�����i��0��D��0n�9�<��f��	|��<����4�$f,�^v!�W"]��d�if$���ׂ��y�]�+S�����Y�A�콝�,�u�6q0.�'��`�В�����Z/���ʹs�%���U߅_Y� ��G`�yc$�~����Y�����|Bi����%L�����b�-��W��|5 ټα>`IZ8�\E�1�ʯNY%1�W(�>��/ЉY���Ad�wDN�N7�r�v�}/�2a���G���"�P�]s�O��L���鲝+0:�zE�v�*7>�E}���������ora�fϡ�g�;���_��f/]� Oa#�����W����a
0jY	�,�Z�����a�DSդY�A��x��5������,j�g�?&Eru&����$��aC_Ѱ��5Mpi��aw�+��oLG�{|U���R�ݵh�G=�ND]�����$=�?س;�C�9��ƓM|J�3���3_�#��eY�
~lu��x�㴒˨40��'՛�Y9jc	�F�а/��l��5rTT�6G���FX�Q�a/�nzL�#+I��R�����j��-k�~S�����\��^/K|V f�^ v!����/���z�������	���`�FS7�D�4^�a�.x|�C�:��g���r��s\��5u��uA&i�KI�n�2���
���u����F�)��;k�����^����P)h̪���ύ���G�(�9�Q�Q]�7>A�F�P��[|��[�jG^<�n����u�58^e�I�â�J9����.���0ǟ���F5��pɡyO�$u'�$}��r[�1�S��$�Q�z ���Ŏp�Q
C�r�D���h3ԑ��k�߫��j���)C�0�n1�Gw)����)3j�K�>SeB�Z|8�m�h�m��?����&6�N�u��b������(�H۫s[Sן�HJ�ՍF)�u�g[|h�M�^�����+�Y��$7��t�Ap2>x�^��I)J����PT��g�>�yt���P��N�i�6	�������ՄO�.�m!�W�1<����T�z���qߝ?���52���}�T(N�'e?��N{�$�?��q���U�ꨥ��W����X,�M���}Lh ���/@VI�P�B���a�Ư�e��(E�{o�h��@Mщ��!���O0tc��IQu�'����tT�eb�\�#)@��3�y�.���=�E:�4�B�h�F3l�ē����+�;��rB]y�9�4�u��(�s�X7@9��@@�bQ�l���/5u׻y��x���+��2L���d's+�WO7�1ֿ}w�2�.���-]�7o�Ṛ��R&�c6VK�^M�4 ��p���/)�z���5�r�:PCMԛ/�������O���������,��̼$e�@�=�?]A���C\�jx� �n�������h�������-`V��>�A7.�M�L�Lņ>HX����E�L]*\oŔm�jK��/q��'�Bt��[�ܶ���GbX!�A8��:ZE�J�ɱK�+M���q�ں�	;��<��ܺZ��$�/�BY�Ex'�nr��{�O�� �
���[�0�PT	�d��~�-v󫙈�IF�����&<1�Ұo.���],*���C\MQ3�k�|C9��f'jپ�����)��� H\ rعv�o�t��&`�Ӷ����e���T���jw8�K�F�Ժ0C���kS;$	"0Z�������Zmw�}�A�#�uy�,9����^ڧov�S�	�Z���Ju�0��R~5���K���"��iF��}`}�.e/P
`�����
�c��S��C�(�>d��*���nO����5 ���XP��vM��Y`�Mͣ  8Kߝ;�� ��j���q=R�d�f��{H�֐��X|m�:�����C+'��I��U��~Y��fS�F]�߬��Y���hc8���ciQ�L��J��sb^{>l�X��N�	n!f��"��U�"E�ɷC��K�b립�H�x˖S񫩪�,)�F��R���mrf��E�s�ް�i�P�6$1h#�6N�`&�j��A/9G`�� �=�	�������q�Hz��x]���KX��ՉU�Qg+(B���B
P ���u�d�e��Q_�iO>ݎ�@�Y١F�(Zﾏ��Rw���k@^ӭ�ځ�G=L8��
(A��jʓ���yՅp���%��K���4|��$�wh�pжk5���/�Mx�|�"������:ˤ+��@FP*C@%�L���U�����V ���p�(
Q��~�p�u��t�yG�^cb �a�����I�0˝����-���/�6x��cz��L@��������Y�)X�)���g���jΗ�: ʹ�
����=C��?�P�.�O��I����G���"���������i�p֠�_��w%��Tfhr��eYay�fd����ZГ[��ۀ�(1�e�I)�=�h�҉ ]ǵ`���x�/��8B��������st�g��՘1^��q��6�B"��_ϣ ��P�؆�޸��Ce���:ы�I-9�?���_���S�_໹�L ̭ɇ�\�342�R�9I�9ǡ�D�x�_;nhs�H�+�¥���6�Ua��(�(��u�������1��<9��+PZ?�%�_���a�&Z���\N��J� ���\aB�r%��*Q���9� ��ȕ&iA�ʸ�����-i��?9@��_���?�l�,3�C��\cFϮ'�n~5���HFT��J�*��a�Ͳ��(=S��[aª\�@m2�3W@�y�_�#�7b!��>�V��0u��e
�����|�Lv��(��I-�b.�L���e�%B�V�n	��'�T��`�^t���w����iX�\�7r3�ڼ:�7��������ELh0	�|� �x���;-|��Vߨ�%F������6y���a�zM�� 6�=����@
�?���a�me�]���I�9ӫׁ�|h鈹
H^R�P;�� OA����&�4� ?\ub��J0�id�#�q �ص�R$��;�������+ߥ�4�j����%|��"6��&ῆo�ϯqG�up���-����q�=9��!kJ�}I����w� ��DX6?p��b����\�(/$3��_����O/]g�������]�������R<q��D%.��7:�;��!`l7�`�^"��ܾ<�H�8���ʽ*9��fJ^���23��3����G�q�,I������wA���K:{Q���9gr���:x�5��4dc���/��3��~q�x�Fݴ��$HI���$��T����jKr"}q��L�4{(� �@q"�Nz"$��E�~~y��MK)�����Ԧ
������Mv�lb�(�|�+ [���i@>�����z�9�Rv��]�Y�AYi9t��:�d����8�!/E�wc�+�`E��W l�_���;+�t�#�t�~�zz�!b�RP�����,^�|�_����@�߼��F��2����7AhV%ud|iP�Mhcd/������ �>���ۥ�+՘�܃X��V���o�W�5�_���FDԉ�kHH��`�������Pʣ��Ŗ���� ��fj�3��	x&���\a�
��8��g˥��D�K���6_�LtA
07�UiM�Rsz�#�y֡�����/Tık,��#li��g�L��wM_'�G�:�����@��״���� '_ґ�ۡ�1ɾ/ݖ}µ�d�ކ��)�3r�z���:�;�8����SG@� 90�i�*����S�2M�8h��h�J�����.|�?}cѢ����|f98Ӝ8�v����T��<m��b��J����,�+l<���o�����G��?��&/��<����I)V�cp��`̎��c3'�<�(4����B`��7f�������Pu�l�ɚe>P5kIK,�/�-$vK�Y%�i�j����]+�v�N ���jN\?�gr7fūp%t��ͷ�,���2q�ͩD���
,��}����ϙ�� ��UB���,c�u�?�����nKI��[22;�5�e�í�/���6��tC�ǉ{��R(��!D�0����:|[�Z]�0MI�M���>�%M�����{�1��_��e�g��R�RvGUB�P��Nq�į�/��ՏVo7b�Qܨ��\��h\0��g���R+�E��]=�fc!e(�6 |�䆮 _�C?Q�L�&[=��8( �5��EԈD����@��w	�Jjg�ᐧ+-bX�PYp���a^P1����	���gw�Ug�0�N���>�7�GY����7WZ�P287q'��xk���G�Q��h�v��T�S4��>6���ӈ���,n\��G�15'�`�9��gZι �͙�G�Y��Z؍g�B&�[�b�돭c��@#�pU������[#L<\�E�̟CJF�>7�r�WB`}OY�-ɕgT=/��MF�c^ᘽ���\���qu��\ӷӌ/Xm���"���2j��'�|*�BMZ15\Vկ��ƛ�3I�$uw�<��N?���ؔ)�=L9�,�JE��X���O[
B.(�Q���x{l�� {Q`�	S��A)�EF!����Q�VTI��"Es�����vȲ���Z�j�!����m��Y�+Y�w��"��	��Q�6hb���;�fwh�Q{���P�2�NV8d*����<$\]�bX}��U"�E��)M�_ڇ�G��T�b-�<_��ŭ|Z�.ƃ}�u��?�{RčR�����(N�(´�`>��!/��rc;��Aз����}���JLj*�lrCB�gXi^7%�(�:��]z�ֳL$5Ϩ�&u)M��^6�X@��
I��lQ[�zs��g~�2?�T��)P+s�Q�4̬���w�m���
;��
�j��i�~�Ê��^Jؐ�q��x�h��M}	��@n|�Z����cՎ��-x��V�kv	�QZ�xkc��dI�K�,{���?W|�����;9,/��;j�Y9�S��R��њ�X�����M��LȾ�Y�\ݞ@���
�J�52��!`5a{	�̞l0��ޕ�gܓ�m ,���Zy��dj,�n�ͩr}���U��9V�u�Y��O�=�M�7�b�L�eL�A��SR�1'n���=)(P�	��1�R��������/rc�7(��BÀ�44G�`�@�X��v�8S�|�$�`��i�R^f��� _�f
ܺc~u����"]?����6�d�<!l����cr�~�bk���2@�U�	�%Ų,�;ۓ\ ��N��� ���1P&�s���'�ܴ����"s�F�ǡo��b&@�gP>W.�k��j�#+�ja��y�#c4!u��9P*�R����FS͍��Uߑ�>:�w]�٬�~��=���^:/.�����H�A��o���%�2��s���#�>�H 	4R�
�g�%�z�0��A�z�_F�S�r�9�5tH���x������XM
8�%%������0uӘ9�έ���;�o�>*��R��u�um(�Ƶo�}Zȹ� m� +;���ȪIy�iCb����E�r,ޭL������Í��i��x)I���NDhSQF "K��>͋E�^�iT�+�{��%QR^~j7���m,�ֳ���d�i����p���nh����!'�"���]�*���L`ŒF^I1�<(�����tF ���3��%1��刘����B]s�^�u8���N_�p�0F� G-h��Ϧ�a(ss��s�a��n���1�	T,T�̏�YGȄ̼bsS����k�E{��j�lVx�H0U��Utpp ����©�8č6O{�q��KG/1�w�)����E(��c�8��2	�oLfp�Չ�]}
���蝐�í�B��e�o���LB�-p�H�z�{��W�;''�Z +�Ȯ��x�}D�z��S�r<�L����o�}6]s3�]�����G�Ab��1��ϵ闑+]3`���Y�a%:�g}�?P�0�|G&�뾿;¯���q�����{�X�6�4FR�h����AO�~Y��w�W3%C��.�;\z(���Q��O5���8F���8�����o�����;��V���1B[[��3��.���	f�=��s�:C</j�� :n�!�L̕2�%��/Vݑ+�m��A����v��Śc3�٥��]�0׮^�!��$�O���M��Ϝ�N�m+i ��K�7�w <��-��|�]�Y��B�6a�l}a��[�G x��O �ST�ﺪ�݄�=�|����;IݶN0!U�¾�u?a���g�q�mU�o"/1��wU�t�'�B�9C�~���js4�k��g��j���̤D��3�P����[�ȷ�q���<�������Z��2cg����A����+��[S>](�;A�'GPwI�cR��O�s���y�{	)r���h~bɖ ���J",�t=]�Mh�\E�k}e����9�h��R�h�i�
Gz�Hm�j�¤� �Hn��BP45ɶIu�������J�?�h�g��NJ�_�\�_q���ء��:ۮ`���W���X����dE$�.~Yi�y"�+k��B��C��d�=�`�3^�QH�֞��=D��dtA��%��@	խܙ u����"41t�B�nU�pI��r�^������^JN6�Ґ)ā���R6qI56�7�
<�=�f�S���~�r�T��X,�2�n���T��	q��Ԉ��9d1nУa��j9�#�c�D�C�8��&�$f4mnj_3c�.�Ay�QF�gj˅G�;��	���r�N��N�.m/�-t"���k/Ęƅ���5�^)�q(K=��ɓ�V)�#��|^�����Y2.��ChuK?��0�y��BN��ٽ��cF�!e��eR\����itL�X���LL@K�$���¾
%hE~���(�	ߪ~I%����]��U�kaHe���׍[�*֫-�/�b�*=�L�*�'#�O���ڠ3MB�h���*�'`iw��6y l�H�nRwF�h�-x�VX>
�'��*���C��mл	�d��S���'�/>`�q:��V�����p��@�2�ؖ%��v�ӿ�ȡ&9��9/����W�OP�uu�#���l4Y�kkİ����:4����4��:g�L��js�y� �5��yhlH�=�|G�ei��!�;�s�8�ҭö=������wr��#(P,�����`\�$��A��$�,왌e���2DȐ�pm5���.�V%��3Sl�	��vV�3��5H|="� �wEf=K6��)OW�
��E�tc�';������� ^�n����i��5 �'�n��:��s��;ưk����3�=qᝲ��z��r�M�r�qV�&caL��3�l���1�+a:�Ʀ�1r'�+|���֦��������4	�̴�v \���9cN��E�[#_�̢+��I��,ȩ
ڼ��`YOM]R���fN*bUl}�Nǫk��DZب1g޹7�μ}p�o7� ��O��&���Fe9	�����g����)�X=51��|���~���#�䂲];UR"����fta֭���4���,���+\�ϣ���ͼ]��V;�Fe�����-Z}�ې�*s��@<E�i^)�+��;�hv����I�[�Om��Փ ���T���x+Ws$~�+�������4&Ua��ݎIԆ��]��-�OMMk.��{wp30�w���茚Js�2d�3ƨN G����C/�*�RS:*ؚ��e����m�ͯ<�\�o/��af���.	�8�>��ȷe��F��]_���{o�������p}Z�6~a�0C3��R�¦�e!���|x[F����@)�ʖc��da�7���De���A1,Y�{3�����b��`��=�*N��0
�wtBW<��՞`��b��⛫Z�	�=��?�Ҙ��	���>��c~JA>r��J��TG�p y�}b��S\�z-u��Om .g��vAr�����{������K���k�����8�=��~O�?K��R%�NŇ�)�mPM�eO��ٵ<��L@R��Ry���|�) ��t��K%:�!8�F����A��ᤉ�����l�˙!$�����F��(�;:�3`�O*�P��H��~�Q������P�`�M-��{��k���
��d���F�F�]�����5�St��w^�g���e��Kl�Wz��^?Z�:�{�5Z�*���R|��4�ɠ�'��fܶ���+q �*�;��R3*�`ͻ�r�+>g�������o�q"*��{���#5���=�.{T �>:pn��A-�^��`g�^@���A��S`k0 �9]�uz�y�*C�\��ڍ�X�
R�����������f=n��c9�|���&R�D�]7�n���]%lK��*����0�/�<K���Oxϕ�W�fݭ���x�Zw�]�H���� v����?B���H�kcr�y-}�˞'h�Bn����>�]�t��S�IR�.Ɔ�[�}Q�'��D���&��D8�B���-�j�*<s~$М�)�"��ց�2�0���0�"�;*�~���C�`�g�}#�?�Rݾ����4<�<���d��2K)��9��r�/�' ��(��Z��m����-6�jX��ׇ�E=t�O#�\���u*k�ŵ��W��W8y����3���iBv �!�nj��+��BE��:FGrr�;ގ]�
�ӭ���Ƶ�PM$����ۨ���lU�xQ "ꅣ��8lA��i�?��%6�o��4\��OT�H�Q��D�?�}	�t��8J ���x�"��o��h�Y�dH瘭ا�͢�Mƈ�/��y�]b
-�J̢=z	�I��I�+�uh=U8,�cv�&�U�4"j5�����QީK�V��ƾ�"4��{%0�Ƥ�y}�Gd�_<Lҏ}���d�_���+�.ް��ΈS�0�s�[ �U�~�7ʚrm7T+gW�s<�LOn���&e�M/~�'`V�]�6����rp��|�7�EM�.`�By&��Р�B��Xוr�	���܆�!��!�np\zV�k��*�5z�zd��fvh�$�-Y�~V��J-���}"
�����:��o�W�3�*��;=�}P�Xа<��(��Ѵ���g9\�a����J����/Y�B�&�l*a&dPۄ�.uu��P]Јa]��h>�N���O�l��w7D��c�|4`Ks�m&JI��'�f��%��k}������׊�o��c�K8��1�Ö}�E��� }�������ȡ��f,l��vљxɠR9E��}z�L�v#�b���fS:	���.~��E��O6B����׀��{�YGӱ��`��lLI�L��0P�3��M�сf��b�){M��Br�(
�y�+�w��
����B����ѫvа�ec�Y栮���\��o�z�aѯ2�� c�{qǬ�������ϼI#�qV�lI&�:|�M�����ښ���B���P:Ǩ`��`<��"G�W#Γ6
�������{ս+D��͵P��"e}��{��#q��-�Vo� �;3�?�`��u��(��1�,�BG�]�[�{/0M}�ls�I�V'��c��������I��q�?n��3xC���a���hQ���b�d�fa)a������q�ҽ��v��p�/���%�1J�b��ޞ�X�B��iD�^���լ!�tY�~�)M	�{hO	��V����Dc�_3�D��	�a�*�>G���5���O�gϹ�c�5{JCtG �o����wT��0��oU�ѴplYt�>�\��{��,�JR���D��(�n�RI}X�ގ����w���C�	LlF �Y��a����~���Lߡ��7&�;I��&�tP��R�'u�]8	TO@���ՙ��R��sbh��<O��� ���y�97'܅�S���eA�bPX��CKNl��z�D&v�`����N3��D�q�^*�^1���L^�ToP����ab�
��ª��j���Z@���	��.�%�n�ci{�^�}J��UҪM �_:9����2�Q>d�c`���ve�A���y��q�c�v�l�0+��p�i���N�>r�_W7�Q�����Y��"Վ�e�d�y����e�X�X��RW>�}AXO��|�oNAu���d�*���bO�a�o�B��/�@��'Ё���*���&�j��>dk��7aL��^)�W
J�l
�ԃe9����(�>^���Px"#�j�A �C\��tթ�9(I6�?���DF�10+@aë�yX�Vffh���I����p��H�8�ZV��2E3�wAP۾�\.�/��$D�֜�� �0u�m"k6�t��v��z�R�`�)_�_	�Sg@���{�ת���X׽�N~ O����W�����/�K4r�L��������GR�ˏKs�H�	�ɫ��yCؑ���qJ^�&b6	,�0X�I(��'����xL������~�#>���U(��ͷj����`܋N�����J�o����t���X\��}��}K!�$��L���ti����N�֎i.c@!��ґ=o�x��,��d�5t�� �d��\G�L�ȻW��81y�&��,��(s׫�ٷ�JU��k��Hd�:�`�7S0��J�E��?^�-0D�nH��m�W��X-��p�6n$��w��e����!.{���8L�ȝ�Oc�9����G/^_�����P�dG���l>l@��oG$eN�tZ��١x�g����2���|�r�K:D��l\�y˽y	!����a�+�D
�C$�=�i"e]��ة~��#���y�'�=M��1G���^��( v�i�ts�-v%�F2f��$d�F��o�	�Ŗ ���\�D�
����M��$�o��=0��9J�����g�iG����S�A�n9�;�<-,�i]��;Rx��q��D�	o�O��� #|�;I�f~��$�S�L�N�&v�d�=_O�_�m�~Bր��b-`:�:5�Q�a.Ќ�#��T�a&���7�R�ԭ�/�G��id
�\��G����/��S���'����j6emWp�
����Ȥi�[ʀў�����Q[��G[�
>���k��V	��A?ueM�� �n���ք���!�3�>��weOec� 0	j��2�����.���'��9����5����;�`�����/sg6lC�ʩ��);Z#����?�����+��ߍ��N�w9y�IxTPBh]�T�ey��ۑ��禡r�w_�hܺ�� l�ɕ�eZJ������>v �/���W�sm-��i�߀�����iv	C�QI�ڹ��p��K>���>�(����Z�QoF��F�D�oZ���)M��zݖ=o�40Ay2-�4cH�T��vR�44˘� ����~󏳒�d2�������t��3뾲�����y<C��+�+�������l_>b<rÏ#�|pm���ro�]u/�E�0>"qY��Z�����Z�y{)��21��	�{�D������\��*{�K2��֩�"��x^��˸?�^qINk��5]M=���ɘ߱�7�^��R%H���-eյ��Q,d�� bد.�M����:�р����wi#�	��j�2������D�!�n����*F4~9��\m�vw�x
�#��w�8�{;St�ﺗ�ȴ2�����dN�U��N��R ���RA��
)���\V#�7~�D�WF����@L�8I�nc�>��P����g�ۆ����T���}1�GZ���r�%/���L�� �W@e�� ��%�h��� x�ts��%w&�X|܃H��C�a[��Y��o��&Vh֔��]^W6��������)q�&�|G�����Ua���M�1�Dơ$oL�������y�8������HיC������k�n��-p���˧s`$�e�:���i[�w�Ꮶ���x |�%>M��������w���9�R��9VmCG�Ϻ��g~f���{7�:g���é΋�B�@�1��/�v��ɓ(�D�(ъؕ^ �7E��ɹct���KVP+�N�]_��?�y��p`+s��#{4Aȝ>2�˷�����-�v���Sm�R�z�������d�F�v&�uYqg�zY��2�J�0y�Q�M��UF5�7o��9�u��r���餟J}B(�L~�Q$;�'oθ#'�j=�%E��Z���^
�0��)���GJ�,���]"]� ��(���yx@5V��hF��K	�5\��e
Mm��c����]��ԋ\�O�kF�=������|?5�$�"V��EB������bw����J��LL�2E��c���!MOC��E�,K�|V!��u\?+ڕ�B��-b��"kֿ��b%:
���Vu���kN0H��B�VeudM�h�!�M�t?Zs�����E��l�][K�k�H��6
�nCMf��)P�4��`�ojy�!�'i`I�]�[��tv ����3������4R"֨�R3����C�H��v�Ǧ�����toY�8�t���df��`�+��sV5]�� �`TcQ�D�8a������7";���ֲX��v��(C��<� �-4%�z��iQl���	���S�,Y��$�-v��'e)s�a�2�-�8�6\�b�����-?���z����M���
e��O�lI�^ؑ.�I2޻yC�v;���`�e�v�y9c�;_�L�B�ܣ-����w����p�H��9��YBx7���rplk�	���/��?�d�:vs
R�JA�����`�'N�K�n57�~ȟvY ����aoۦnV���%�o������&ݹ��FV�}^v����Xpn|�s����[�a�|NŹ2P��<�u��B�=c�J3h�}� g��5$�,�m��ZO�\˳�BGL�`��u���k�/���?�72���-/���5g�������ո�pbz�Y߁�(0�s<	=��wĽxq��C�c2�u�׵Ď�y�h*QN
dP%�XI{4�~z�2> �~Jt;�:��"�aג�U̶�=֑�u�K$�Ӷ荗�(ԐBB
@�m�ė�;H��Z��yO�I���A݁�l��_�>�f�?x�;�r��X��T����T�_;OS(s}~��׽�0�᪽@M�UV��y	����?�U8��I����m��}!���p�Ox,v���M�D7��}�n]9�d�I�0?}>��V�422��xy�-�xQJ��=\GuT��Ǧ����8�j�o���q�tXu�=6��`œ�_�M�y�9�	@V&�]_���쾣�
��	��C`r�[�7�V�5 S��P�lS�]��>�^{����� ���PJhZ���+?���4��Ϡ�������j�dq-Zs%:Z�	�T��12}u7�t�jrZ=�q)���v�H�oG�#��M9�g��iOe����˕�r+���g} �����c�<$�@�D�mz('wB���J@,��N��6��JV/�V�$��oJ�|߂]ac�y��O!8���m|���A�- T�ϣH~kQZ@�� G�-�;XZ<�vs6�dRɃA*OLcZ�o�N3m<�#E-��p�.�M`�L�K��V4��d!�;W)39t��~5�ǏH�d�0"�N��{DX#v�2�`��<F�v�+��.�F%K�ʩ�x@t�/QWsf��t��kv#�����B�����JO}�3u �7�𱢖��T�ѡN.MV^�dxvBi;
�O��o)tse%Y��f{L��!�����f���C��#�%��M}��Ӷ	��E�e!
J�s��t�k�n*�����X�5��=vG��b�����RF�����M�?�W�m���'�pZ2 ]\"�G����Ɯ���e��q�ۆ�\�����[>4V�@87jR��W Q�0(&O�}a�22��l���%��;��eh��j� 8*�1���2��0��ɼ&����[��'µ/�Q���K�8֑e���4f��#I�o�u�[�ڋ�J��8��c�ۣQ\�%���t@*���Y#9�i	��E�G9���;�%;#�E�A�Y4%i��J0n�@w�����o��E݋�bk��{1��Q$�NiŷE��n�i��a�e1���
q�g
,�N�m����>��r,	>AT���>��Ρ�\_%#'�%�k[rʋ���Z�Em���Uy)�g�(�H7u?a�/�v��~u���(��	����h(���,{;��Q4bU+{���-��E�s� m|�}1�R��k����������OD��^ò�3�Ԙ�:JP����x�)�D.<�'d��N��-Vubg�z���{/Uq�5k޵�]cC�޸n�6P++�H`�ӑ�ZD9���<ٯ����d8��M�53#���lV�]��Z�a�� �K�;,�$�C�V�wBTX`�z'3ڪR����CdC�/�+]���P�Gү���1�+�����3���2!����r��V�ӘE�ȼ�qڄ:�
]Y��jQ��'��U\/��7�O%p�@ ��_���u-�V�Z��E�"Qw����
Dn�
���1BI�}C�N�����VAtN����p�R	���d���������@�P z{u�t���\��M:����S4FE���S���w�yT�lC�E�ŻA)J�1������+�b=Y������(�N�;=���B�ե=�e,�g*��U�Тܹ���+�?cŕ�aɽ�N3\����00�7�F��~ߓ�?�o3�g��%��i)i�ŋ��Q2۽���g����7�I�L�j� OVx��K�d0F���S/�X�r·0/�n�pzz��cRN�zh�W�42����� ��W�`h�Q�%P�˶.V���Ge_L����v��������̭�S��Sb'j�{C���1�2N��6p�=ޤ=b`�E��SUá����)3����C��5]��7R�+��v&S�D�Sǫ= ,�RS�xjQ��}�XV�_�{VK9O�<簁��]���d���t�!4~t�N
���/�Vz}���珮��c"?��e<O8��(eg&���+�CD��l0v�؍v�^5�jAV,����b�XR�A�fCߩ��8m��G����.T1R���i�,�m*�w���	F�$�*�[�p�A��@��zp*� �[��ܥ�5UN��`�n�[s���A����⾮l~��W�	��v���fD-�*�=��l�`�&0����:�R��קZ�p+Z��Ԩ6�>:�� �R"�8QY�s�S��P9�2�iN�|I���ŭ�(d9+K@9�1c{���3�����D�NL S�+��3�I�H�W0݅K��qO�w��{+)?糁��F�Rc���v-Ķs0CБ;�����c�PTb�2:(�Gpdߥ������[���*R�Xg%��X!��k�3,f'ͣ����WWt��aoX��Sێ��
Y����3����NN0�b�h2��\ ��X�2t���@����� ��ׄ���B<�:�[1ڠ�H��tr�] #r�6�85�IDv����"ù����H��~7��Dm�"M��i+��-������#Nd�/Y����'�1o� :s�~%�pst�sJ�T�ʛ�*�ڼ5W���1�o��#1����'P#�Z���]�˕|��d��,]��>���gdG�z�'�݂���>8�N��K���z��`v37_h�����<��� Z���o!JŠ�E: )��?�|*�x8xG���H�}�&G�L۟��-^F��=sd4��q�xXC��5�je`a#��)�Q�Ǝ�7v�-�Q��K�
��.,�d'+ťV$�қz��Ō�����j��>i���|u1
8jqv0ă1���d�v?�WHB��x�`�m�e��=�k"W��Ǫ�A��.ښ}���0T�ܔ[�_���`0���r:��tFP��Mp�e��q���J�������u�Q������ߺɎ�C�I��^��V�<D�-��Zb����\������q�B*�V1��_�/&��$H�1[�[�F�b	�7~J{�a�y.tȫ,��z��Շ���t&4wL��%� �� �Y���ب�tt-��b_�,ALh���i����D��(&X�pi�s#y0 h{q};+#k��J�ƎP�~k���ص =��.�]�R��7��T0 ��gG9��{	�]yBx��`S $?�t����&�Ƶ*(���j`��F� �ɰ޶@
!k�뙱��7i�1g�L�"O�u�۫�b0l�� @��a�)�<�$o;���-9a�A#�(]n�'4F�/8�״�s6X[c�Xb��@6n������ɼ�aRpd��j�4�	Zu�d%z����.48��bT�l�g�7֪��{x����-�q���	��b0a@"����F?/��2������O�f1�F\T��������]�a��fB�a�x@�jx���.4����P$�|���W�*�N�����!�	𕚺s�}���V��Ja?m��͟*�q���o���QW���C��{��-���
j���h�=rV
�m�h��B�k
�@5�9��DЃM��q�?ʭnW�x�Ԧ��\��,��E6�t���kS�W2��&�b��\;R}t�������>bA+?�
_.Ưu
��*ც����r�
GA�Ɗ;���:F�A���}�rD���l��P�F�Q����b-I�1*=y٠��� ����o�Y*��ũ�a�.��ȥ*;p
i3��C�#s�ۑ���3Vi��	�C��̻]��Ͱz�"�+!�䂮s�"��pԈ������m�:���@A��ŜZ���_��HS�]r���7�&܁�V˞����F�;SG���%R��Rg,�I^���R��g @�a��3���ѝ�
h�7}�,æ��
�	��X�iՠH�:�q�^k��0�?8���W������K��r�(_�- 6�w��Gd��u��:q��I�/�Ѓ+�@<���%"�v�0,0-Z8��>����m
�D����������y���!
Z%�)�n���t���@rg����
Go�'	��S�>����Cp�����`�43w�:�']�}�tf�@$�tP&c��8��Ҹ���c���w$q���Z3q��t����G����Z4�B�gmo�n���JdI��R���*L�q�Z����9N|}iF�R�F�V+���1�a�O��}>�[_f��3:*�����[�h�4�CR��yP��(�jR��`���� �Z\nð�T��M����̕�_ �
m�3F�;��'��M�4��9%"�:���tA�i�~� � ����MZǒ\�}�Zfe�P9Ξ� ��Z9�yO��]B�z�w>�X��Ip�*݋�M^z��^�������
iK�Sz�S��-�A<]4�D� �1@x�,�w+�~��e!;������]9��F�t�&n��C��x��O�#�2:a�$�.ϛ�t��?(^81~m�ȁ� R-�K�8��������h�^�-OUP����A�eN�چ�1(�Aȏ��.;���2*��֢]Pk���K��:�%ǎ=��F�$�|
>�H�J~���2������s�'Eg@�m��.U��`H}W���x�>���m���:g|/3�@�CC}B���beޠ����(z��*^��K��{
�<m˼�Цq�<-_�w6W,���a#JWИ���@S��ID�cA�'�11�u��Z��|m�?*M�K�@�MB���O�.�Ѧ]�7���h��;�I�5n����T���nG]QA���H�k�VR ˵��<� yӃ��[-��^pԯ���Ζ]��C�F���1�q��3�㢠ʉ��Ɵ�b�g���l�#�=��9���P�O[7��<�Fb����������lb _�[͈��qwk-�<�(c�	$�Mݏ�����?u�H���#y�� 3-�/��?+��pY����`����ׄ,�d�j��u�m����������f]�w��L�A��=�kP��� ����P�� u�S|J����+�f���\*�«���r��©���,U�4���'d�ĕ�ٷn=���r�٘~iCt14�q�<��m���	t�T�S]a~��8nO�.�k���i㒗���)��j3T{�<���U��4gެ���g�vT�?�
��J��K�	l���Z �Z���_+������%'�7Y�<Y.,�f%���I>sK��:�y�g�Q�P&Sx��{5Fgc����}�;��l3i/Y�u6~���/�;�B�0��� W	�[_5�QV��)�|��ID�:׌��V�@b{�v�؜�՜�3�\:�u�����:��ۺ,�N���4ֽZK|Y�s��H�CC��:�h7H1 �A���_�n�N��	;�Q��6xC��ǿ�XJ�i�����dl0�����	o�1��o _?rD����o��q�{�v%6�-4������:��L;�z�J�'g����՞3�_��K7u��̟k�ؿgL��@���M\I�$�	e$mo7h�DjR�`0�$�+�ec$S~*���``Tά�'5Té��L>W��P���q�yoEU��n�T�A 6Ȝ�>�ZFr�&e�B�c ��}���Ӄpwo�!~~��౹����o���E���G[o�%�k!�<�nM��ِ��#�A� ��+�j���dH��6j�|��1$��Y���xS4w	
�AU2�t9+G�'Rq�����$}6:5cU.'��K��1g�6��r�:y%v������O���#T}���g�׃�,&tIe��3mfMrgezo��`~�䖽�M\��o*A~��R
x��;����Km�?��}΁���6�I���r�0���H�aj^���^�v�*������m���p9"�� ���<D���w�>b!����5��#G���xۋ���%��q"�m��Ƚ�h��Yu���[�n���T�6���	W� �Di�ߠ���GP��$��f�B��,xѳ��Ӥ}����h4s$6�ژx �K�-G���0�nϢ\���q�A�Z� �jD� ��f�ffolLg]jN
)���b���*_���+%����Ō��}���dVrE7,�tu�c��ct+q���0fx�c����1�fc5�y�σ�л[�J|\}æ
�؁�㲎������E�{~f�6/?��Ҵem��<{�P�DQ�ò'���W$���l ȩ?7&���Q(m�V��������u:,�{ǐy���S��RCo�"�s�q{�<.�[�=
�T���r��cnM<���~{j]L#x�<��1��k��t����XXE�/��������.��Мj�8�_����q�e�uw�"�4��fd�p�����N����H���p�=�.��Y�ag#Tu��Nx6:���g����Jxp=vwt�GTn���
�����{F�E��z���nR��Փ6����I��ؖ����4�k.��Ld0�������R��7�%3��+[۷A�Uȳ0��%ч*q�'d��j"���:;�������(�T��ޚ����j�����6���4�(��!�_f�f�����P=�Df'��g�D1��1�ظ��S�4�G�N0�p���)�v��[��,�F=����z�r��"����/��y�P��Sɣ��tYy����n�B��c��LE�(���9e9����N��(��ٯ��IQ�b~�oLy�.]�;���?��ؤNwL�uϡb6k�`� ep#���h��A���[ܟòX ��5���'@Nt%J��N����nqҲ���R�XȽʤ���x�/rw:�t�!3͢quȊ)u��$��B1���zH`_��s�;��,�/�	8��9�y�Zpq
�w��N����̧IVJ*��*`�	�yB�������b��8BFN�T���c������/�ד;���d�͙k՜�p|��7(_;�	��Y�gk2���
7��C�g!��9~9�/���i�8�`�v�I�d�':l��Eb������4�G���׮ٱsJ���*�ږ\2�f����X���0�1{r���M������7׼&��j�L ӯNߩ��j
���w��o���^D�_w�
O�w-qqz�K,CL�
V Hr21��^0v	6$�)s:�i���ׁ���R��u^1t��
DLW�	p�ْ�`�������7X�C�N1X�:���rc�{�_3r�TO�i�vf������ȀU呂���?,��ֱ}��K�t�o=>�r�o^Р=����7�Yȁ�X� m>�B H���4)���|��4Mkt
_�q]w�=��z�W�:;/��/��r�����^Pخ����/�\��~�đYc?���;$�l�h�Nn8>`����Bi�ù���R͏XI{`J�-�c������Z���r�h�0�����cm�_:Yu�����=����Őc甏p�~���Xk�<9H��Ϣ�C�}�r>�h��M�k�F�[��B[��1.KOU=��13h{J�c��6������<*�!BA�՚�Z�,�w���S�+̝bH����C�>*�_EϹ�H]�8"ξ�1�|eX�W��*y����q��?�a9�� Pt�?��Be>e��z�}Փh�gwΠ$v�C���&,�X?����@K�v�*$���}�s���Mܕ���jU
ߏ2�|���	�|Q�k�����v���R���<�v�GF+���'VH`Jh&#�%6�G#���v��<�:AF��~G�]�?s�̞���G�upYi����E���)���?9&Ë���7Y��H�I��:������rN��²�n0"i�X�S~�!�6�n�*<��9�P�f5VF�J2hY���h��f$yH�>��D
\R�����o1@"u� ��fb!����J��Ej�j�k���{(#�4IC�~7F��d��]�2T���֞�}aB��:�}�K%J ���&�{iuu"G+�DZ6g�`*UZN��>d���U��"o����}g�F;%w2gn�͡���vCZx�|�	��3��[W�1�/��wx��z�VG�6My�:}c�opCt�w]F(i0��x�3$)�MRj;���߭f*�3G�Q��+�6ފ�&�ʈ!�]
8�b�4���&���2@;��*���/�y�m_/ٛN��j9��2������n��(:�>y¼�c�]O�G�.�~��R���� �bT�m�]����)�/�V������(J�S�>dYp��P:l� �ٻ���90\�����흔�&���hU�`�?�hx�h��\�s�gy�f�l���DQ�mഥh�V+�r�x�h�m#��-�a�Z������ |���[������|��wЇ�Q�_�jG��Ʈw�Ha� ��#󤯤թO�Z��A+� �����(?_��oB�_矲`�:cȈ��z"?>0�^MAI��Dj/�fe�t��d�sK�i`�[u�yf_��%/�	A�F����%�Ԭ�p�m$�l�1˰t'O�{��L���������t��m�g6��w�1	�bq���\O��>��{�l�_ƚ�=9wn q�_f}�2�`�Ym*F ���40
(/G#V���ʑk�C#�� �����Ql��	��]�
S�mP���ӫNf��U�'̤c3�fwtL��J^er��Q��"z�����:]9�8�:��;�x|��@��v��Qs"2��$�v[v��G4�ޤ��Xh��XcR�3�d�J�5��ܫ��xt��9��j��v=���/'zYuU{��Nr�[���T`R;I#�ibd�	���NO�����op왙�a[�?�a[ie�]��
��tn�B ߨ1�s	���r���^̨W64��MQ3ԥ�F+�(�{д�M�#uZP�����8m��5���)�AtX�_V��D���S��6j�'�	�����c|KIr4�k��ڂ�Zh�U��hQ�D����8&���p���T�F��)RC��$����,�8�~��UJ	4e���2�@��1A܃J??�bF��t䃕���f�rU����}H���	G��V+���XOۜw�!AJJ-ߝW~��,R�{�:�V��֮��n�S�U6A�}��}����'��JktG�k�NIǣ	j�A�ƹ���WG�����=%<v�-f�O��Ay��YRDF����y)bE1;pk��K��ӊ�o䂙d�F �s�Ⓙ�H)t ��h%�rLJ��G{�S�X�?9�WH��2O���G�^�+"�4�cxq��#�k�m/2�U�HyU[t;�4�`��Q�#����Q��{���0��Y�������F�5!D�r�"}�m��j��!_�A��KƹpO(���5��4�
3j7p��?%$���M�H�E��H�f}9�V��J��k�J���V��AR�����VW�u2�5B����׏���z��6��?0B��U(���^cMM����ӶqĢd|�4�k�P\��u���J�س֧0mcZ�N	�%��k��U���iM,���ʰ���ݰ�p���Za�����{��.�E:�58 �H9��w�{�/��,�W�)ma���p`�u�t/2�$��ܕC o[q3�X�pmt���Pf;��"R�39��e��Y�D�\5���>1�����׀<G3�m;P[��� G5�CR�bS�%y��ɸ��V�*Z2K�Z��)����:5+<�ʵc�>j`E� w��� .C�MH���8T-	��O-C��U:	h��1g-thߙ�=-��.28"� ϲ�'�(eE���"�[�iCw�^�%/@�#@�+TC��[cy>Ў���m�d�|!{�Ӓ'6>��݇�U��X�5l��e��>g�枾T��zf��mV �ߪ����{����m�
|�5��`|A�M��,�('�Ǩ��_� F,�`^ga��jf۴�1
�Q����I�#٧ہ���2H#��SB]�*6�%�6 ��Li��P!wĺ1�����Uј�V���~ڠP�I���`��8Mn��y��i´��d���S1O���O��1���̚�vr�?��*�+��p������]#:8 �	{�&��訹�x��85�f�%�V���ό�2Y��e���$�5q���m�$�_�R�B3!g���j5i�������+j��F�ؘ�1���͐L�a�T�p:Ƽ�?���Q�R`�Q1�6�m��X%��}&(�N���$0�p�)0�P���V|�̻��M")�'CE'�!s��{B6Iܦ�/l�;���j�*s�e�R7L�|��\��u�M�]̅u����a�c�75�IR�ӯ��úQ��!i	qzJ��3<m=Ӫv�V���B�����0R�T�_\b��)癜pr�@;˯��_�O��B�HYVXQ�oE�2� �j����xA ��D`C 9.�gl��ݦN��פ�ǺC#GI���|s�פ�
ڏs�VJ�=����m�������Gg�o2��'�WG���6�L�o��'��{o'+� ֺ��Y6�~~L��Q�<C�R�
�J�m�YN�:|�)ʓ���a�r)�=��Wt�����
nk��I�*A��KR����kn�Ĕ�}� ����*�$�w���s�Z	��m�=E��E�,Ksi���@�Y��K���<�3�X_�u"�J�ȿF�������@��&��@/�i�/�"&���9�)g@(4pLQ�J�a�U>1��=�Hӵ��@�#�z�n���,G
�\7\ ��rǩ��.����@�;;�( �ޒ�7;��߻nH?`񲕦�Q@���
�p���V�5�֠&�کԢ��|%�@�}��
!���%��mx�%�B�kB[�δ��
f�w��vu��9w���|�8�6�'e* ��x�K2�L��6f�$�(Q-�E?`Y��ɲf�1�1���Ql���5D��.��f�i�oE�R�1�Uf��yfX���pd5���L��y܎ixN�Wk>-��Ó)��[��d����|r�SC3����L�p9�H���"����,*zv@H�?rO��~X	��^iYZi�q��eA�a�0[�� �'�Y]��ӠȘ��$��5' �s3џ^�H>��ī�c'�O\�=��L[T����0ћ��mڍ��!�:��M3��o���X��s/����l�N0sFHt��A�=�kʊ�O؀��tHpB~�.�;}��~�"���:F��߾���S�p�/�V2n�������d�n��:�Чn�lEK�*|�3J'���`%��Lb���7�ު�������R:�����tQeH O����Hb2�}��c�͍������Ş*Ź�'�����dp���;��`�T��M������K#c�:�sBA��݉�h�=��uݨ��4�1�{��٨FEm�d�:�d�������p��Ŗ!�(���]�� /&�����轈��'Nn���v� 4�Y~��@|fk�ԋ f+�4:�<z�R���=�L8R�ᄬ/�KLE��Q��'�ZH	)$�:܄Aɀ�^!X�5d�f��"�&��� '�d~^���elt�3,W�7���˳D�;�;,����j?�1%Y�	Z�K�U��(2�#�bZ���|��k��%��/uӛK�p�*c���~=Ô�E�F�wX�z���t���!o\����`xĒ��r��:G$�\�����V�%zxZ���E�ƌ�`nk��n6��d;;��ƃ�/�M�H����e�>1̙4��8���4
,�|=��f�u�Ud�ܻs%1��
��Ki&S���=�n;�m8?i��wr����S��x.�䕄mEvCC�Y/�B�B��uĔS!���JC7Dn�5 |j�'3�y,������Ls�P{��K���t�}R.�PjQ�B��]�i)"�/!Ks즟��z\��� 1�j��'x��%�GJ
	�A_ø��@���a����3~����c�}zh�vN��#=�b�־/�~����l¥L}���rK��F/]v[�r<�&y������Z;����+����V���6Z�S�5�5-B/�����D�������F�WΉ+�����a�����a����l�.�H�
��zN���k�M���$����0�cT��w;��Pl�%��,�nU>�-X��);V���	����b.��%2w�3dpڔH�ɬ4K�*�В?��H;C� ƴ����#j��YK�nL��,��m�(m��{�%��`y�7���iVZ�"ꢨ�+�<V�hNi�C���ը�	��;�����IY|�������%�����7�� ���9�3�����nз��vw����Me�a��8�����0����s?���V<64R�/"��A���/�ߊ	�ٳ��.��~t�4���K�o��5eʹ�Q�����n&�'Dx�W(�hA�ph8��#��i�wI)��mv�2�&]�����.D&j��X�̦)�zt�����#U�A�w���d�G'�� f��X�o���{dƒ|��U� ���=�T��sH0�-r��yϟ?���6[����r�{�k�wJ���O�aS	JdE�yV
�VlX~ƌ}�O��C1'��=Fu;�w���&�0L|6 ��#-)��tKR6�����O)
�����+j�e��L.T9�<%YT��)���K�Qt�\����&����־��J�3WiF�'= �Ֆ���j�!m��P����#�)�b"�Ԑc\s��&�5l�X���{�^��l�ˆ�W��#�y#-Qb�܎��F�ق�A3��j{�Vǡ.��`�묹�s(���L��@�(
����@����, ���}�5=W$g-��cL�Y�����X>\�^KKC�;X�����n�ָ$�ʢT��%�q�<N������v'��|$Av�۲���fY�K"��G�i��]����h#�DM�h�H{ùC'�}�ߟ�!?���֠�뿂���}/������i��(��rN��E�r�<������y�[A%K�,��K��k�Lw����4��:������H�ލE� ��+q\����P�n�����HL�w��ޘ����xl(��5����f���3ІN�yĨfh��.�Җo�Ld�w�YϳB�$�Ғ���n������Im���8�2�/Y;a
ǹ�F�${�E�mAN`���i��v=۟b��(�󽝞8��q����k8�c�Pn
y��V[���ɺ���a�R 揫�+�pܦ,N�{9�ּMqi��W�����>\���%M�a�����Х#�@"�:���8�C��8�΀�<�3�nJ*EM;,�n�{IOCŖզ8�0��&!�0��{�����BY=9S�-�f벊@�腸h�x�@)tX.8��(���8��N��;|,uR�)ӏ�PE��ɡu<ug胣l��9Y�� ���+l In�"}$?w�ό��3ThNÍT��\UK���VA��%��[�L6V�P�P�ץ��� (�(=�J:O,<&/�,�{�I���߅����G�P�{` ���-����y+n�$F-łs��o8���

�
6@�Jֳba7{\y֐��}��]kK��,���{�î�|�a��g�����_�/Dذ�X��B�Rχr)2�n�Z�J8��_B�W,�ҭT�G�v���n��&�I�����A���"lG��M�X�s�7"\��t��/m��Ѿ��  1����D*�Y��@C�ctx ��c=�®��m'��ms�o�+ ��\Y-����0 �����(�I7|��4lCKi8r���.~��� T{�zȏ��<Vw~�����/.����t�9.x�A��!�}����.���$w�� �^�R���`�ĸ�iJ.^�B2GmVkE��Q��6�����ZWY�*͊�r%�(z�r� �U��g�`��S�(a�����GW�6反2"�XO�r����M���\O���i���?TB
���v�� ��[ohq�F�}�Bم��c) /��9B�v%Eq�"1V�kH2Y�E�=sM�7�7l�'3"u%Wh>�S/�ۄhjJ�w�L��X��şZ^fQK4?�������Ȯ���er�)E���������y�ۡ��H�����CiZ_
B�tfU�8��ٵ;'��P�s�&��D=Η���+�
8D]sl�cr>#!.TQ������V팩�k��j�dHrҼc�mE�����p]f���N�ⳇ6u�7��>5-�F��p	�ݰ�nc)��LYC�N��B�r%xvŇ�W��2�_�h�~����6�͜�
*f( wK��0\��m����?�$b��'�۔����~�8�6�gW����|0S�����=R�qs�iw;@��&Mв��"���E�����]B��a�>p�	����H慎�W����q7�Ǡ��,���on��7�U�x�L`;�&L�\)�o>M��>�2�}1��9�6������Jq	�R��ݟ���W���<������˃xEE�XeƎ5�w��Sb�R-�ͫ�Xn�L��(	�����ŕ~�$�ʵMv�煄��ld�^[3�e��S�!����ֵ�`#��7�6�a��^h��jI_�)Q�M���� �w�`m�����~�;WS\�Q eW��� ��q)�M�=�:���e,��.����I�(?�<�� �8�5bN':t��㰛��{W��8&�ƀ|�V7��>1����0��q��c���B�S[m�p�f�l<��kc�_��Uo>�I��\��k/�@�pDԁ6e��a�F�N�����2V�K-�0���W�2�W�.I��
��W��y`&����S�|Q7Ye�!�?z����)�e�Da��)��n^<��Y�I��z���Ź_�	\G
�aONJ4���u]�7'wnq�u<� %c�-uDon���A :�b�N���ī��� �qE�b-F������V�xO����D;nۀU^v�__�S�����{�H��sg0a�B���Frpݥ�	q��	]r�K�D[\#�%�)��.$�f�v�z�F��{0��L���F�"@�^;ʄ��=:%�+)EO��bg���}��9��AL��>͜R��!�1�x�وx"�ZCq�hrh�§��:�C{f�J���*>2:Z�]~�G�`�)-���CG��A��9�Nha�Ά�g
�%��7	�qD�N�Y�$m��Y�_���GVc"��֫\����HMi��N�,W
2}a�zE�ZS9�ulnt�[�
[�3a��H}�SW{�P.�gD���8N��� k�D��6L'6Jv{Y���+�]�0'L Q�$t~e`mt!��TP����='Rt���"��/���
�ȍ�Baj��m##wg��Z�M�W���bH}���li`�	�8k}��~>2�'��6n/s����i�����2V\��֎�J@D}	����?��絛Y������<K](��@�˺��F�
�'̡/*},T�QbuD��C|���DVbp�r����-6L ��LHh��˾�}�]�
�|����$����r`/�����q�y@�W��<��41�G],'���t��:8B�ѥyUOt�R��:�w��]�����q��6�||���a2���ZaFcj.W5�|5g{&��g���.�Ga`�q9�2��{�%ݸĨ��QL�	^.C��L�|Z� �C�V���u�)=F�B����X��]����p�߉�������ÃB�b-����y�M�N,<�ZDuA�ut��I���FS�E�U�ɳ@w+~��,��%$�!fa�L��w{O�� ��'u��F/�.=�
lp9�u	3����ցf�?���v�+�1ͧEJ�K�#��Y,�6�]��z�O��ɒ���@pk�	�|� m��c?v�g���@p��rl������$�vO�g�g�HW�Y�FJ�0p
��(����ۚSA��W�;{�q�>a�Bv�� ��+ 0�Q��\��滛��9+�z�.s޳s��"|w(�f�}a%���q&��0co���.꫗�4�@/k�t���Z�V=MFRB�4kQ�w���5����X�ݳJ�f&��Ɣ�A���W�+{ �p3�ܓ���r�VG�C��Ph`=�(�.c�WN��<X%��~��Yt��q(Z�&�-,����1M>0 ��l� �#�͹c�MFXV��a{*z�����YKP��ra�|��[�I8֑~C�Rh��yܓ��=����0�P�����q��T�\�5	�"�U;�j��m��{` �31��\���C�;Go�٩��4����Z?Ӓ���IA�B�������m�����Ak/@=C��a�з��]���p)��尓X�{��9X�߅#�6�A\��6���>T�}/�#��3���x�Z
p��:��x�����L>@�.���a� �~]G`�{	�z��$����z�AI<��;��m}�$�#an?72:�ryj|�'�i�1����cUTj��n�OR 5FS���/q���6?����vqM+�|�5��ӻ<m!(�	�"�!*:�9�"5���f#[�w��f��ٟc F2��u���U���&+�_Y��w�r=.�z˨pJ�=iH��Z����n!�� #�2�H֍+��su����q\%�H
��lG�cw���2���^�f΃�}v<�{�R�|M|d����*	��[��ŕ��ە%���m����b�Nlr#6\�a$'�䷭�p�ʾ!�]��o�	`6h���Y鹝�u���f2YU�<".��`2+(Q��=��]�F���Y��K9�<��]@�Ku����X���׬�-�dWR<�k%�:�<��v!Ǳ;/qzM��*������/}�Ż�^֘-~���7�\!�j�˓6Ֆk���=����?�yq5��E�1}���K-TT�R0{,����Ѣ��b�Ų*�k�2��c�q���;)�>������yt�փ�@��W)��[�2�Ɩ�)�d�Q2��Kq&�P���lctZ#�
���^BB�0��p�^�C�^0��5@��t0�@�Y���'��r��n�k�߆��C�id[�����q�~�i����CLE�F��E��
���GdoQ 1�ԤŅ�ϝ6�	_Y�z�#�s���:'\��y$˶�kp��B��feO!J�AZZ֮��{�P�/����@��(�UG���#�`7��R��]����`��s�3��nz�뢑��eZ؂LS�JR��)��X�����%�H��k�D�
��o&|>��m���q�
�=zs�,����H� �{a����p��/�$z��C�X[@wf�4Z�q�V��Է�5���e��Dw�J�E�|'� ��  R���nf8�P��}ŊaQn�]����p�g���J*j{�M��L�y}YD��A-��yI�����mv2�R��~������0�:8���s�	<�*lctK�E0�Mv�1��Kо`3@��@ @��JWۄD1��QfY�B���~�Z�!c��y�e�p�^�MG��,��;�f�F�'�q�n)�tY���]��KQ�"����7�
ޏ�s����Ų�i_cKXN�.I���lX�+�������� �_���5V6��.��@1�a]s$��W��O��lm���#/K5N�fL}�e�.���|�4t�M]=�"I�T������ð)"+եe�ʯ���{��Μ���V�(�Y:+��>,Ͱ�"���(�^��+1W��<,W�$3��۪P��9�{X���"!���
}�mgu/=�7�����"�~����)�`}�Ut�THh� !_rI�����6�{���|%���m�c��5ȨP��,hn����?�%k���h��˷k�������_����L?�P��O�������VIjRmn+N�=��7�����aŮ��q
�
1�(������y��Q@/��Un#&9Xn���Vz�kٚ�sslR��Ji�W*�������ٱ[�����יR�+T��$��yH�2_�$lF���I�k̋@#�qvj�$��I���y+��X���7���#}I�׬v�݂C�'��Ә�k�i8o �ͷ6~h���Y���/���*���b��{�[epW��@uZ l��DT@�Acj�u�nuoP���[�&;8���8�0�n.���K�R�1�s:���~w�1�D��)&����\ޤ�p�(���#�:AYpl�zH����Õ�0
����0귥�z��1����������͔�ou������j�2��}Z�Η���Ώ$|�jvu�2��s(�>#�����|�3xHKM.�x=֚=4�T4\_:j��
p�<��*�H����\@�ב��<��W�Vx��A񠝊���x�hw�`��0�x��{�Y�ߕX����8��&1�����XA`g���_Z�.��ګЏ���,����a8�ش�g�q���!�����\�f�z�0�\�(����~�N��ӎ������y��X���5��	��E%V�,wO1#7��G]�V
7.��t�	1�������cX����l�`������׀x�͖�/ơR�T��)0[���i:=��=���duյه�N�|�ô3mӅ�޷���%�����8�u��I�-�Lf���mak³�
�[?��'3c[ڊ�n"T�
S)�ݩ_�%JzL����>te��Ϣ&��rx*�(�\��䭛����u�r��_l�8ɽ�,�`!��2ux�Y1���˙�aV����z�Ԛ��eAW�#zH�ݧ9鏨
�R�������t�0��?3�X���&w�	J�͑�Ӟ�u����\s�oB�sr.�.`Zj�먅۞���ǄvyM;����z=o�36{�>V��}_��;d�[��l�#���ڦ�n�tW2���T:��� w��H� ��ݬ{��]N�ntGm�J(򤇡?�}?:�2��r�w�����ĆU�ohL{� v_�Fr��I;�w5�x���.A�	�����N`X��!����	���T�ಿ�+���eVW��vҋ߃����x�v�h�p�Z�)�������T1���^��A�3�/D���x���-�va�i.S��:8��Y[�����*B��!Jɶd߷�|�ow�����n`�΂��&�>�����'�i�r��SU�eL�h��;�������Ӧ�k`�x>�oS��]�`�����]9 ��Ƅ�#3���.=��6���S~�=�Ӽ�6]��^e���5o�]
�M:�'�j���R�@G|<���U���Tf����X�觮����G��V��c�@zէ�7�1��X�N�A�?�j��z�co%�g��֗R���!J�G�����tᐗL6!�݅�x"�cD�b�¿RV�
��B�a�s���!i�̭Cx\��.��:�'��M��\0>1_k��0O'~�1N��~�j�m���\�`2WK�5]_��?�����r��<_`|��J�����#���j��4-��5��(���3��L�T�ژ^��X_W��F@X�����1�#�H��k���X�"W�nT.�&Ӽ�s�%��Q�8�P^Δ�}[Q�2ԉ6�)Ø���I$�����3y����h 1�ؤ��E�Ѫt��`���p�I�Q���G9/�?�]�����~Ya^8��y�fn~���} �n��~f6.k�ݽ�sY@p°H0CfrW���
�X;)6i�>.�Y9���"�=��-,*�9��O��^�u�>d�V��j=�G���5�t�؇ߙ?
k�S��Z&ϫ���l&O�������+�>�M���|�D5VZZ/���I��[���OQ2]"H�%��R�ҽkܦ��.z�Oci�"[�@�e�1�(#Փ�:;>��C��@'��a��Z	�̥+����N�a��2�x]������r$c0X_�S"��)ٽ� Kx 6�8�y����8��_A�j�a��çwk�3j��4(���9?��ﮱ��ܨ-�("*f S/���6�rMH��M87���{U�ҘW�(�e����\9k�B�aV�5���!t	~(�u�qמ�~21�^	HQ�������$֊�)�-�K�J����n�P�Lq��63K�U��7�a!W�e��!���A;@TF�ES�? �#�S�nEբx������,w]ٶ*�Vt��1XоeHsV�j��Y�5�����`5��� r�ڟw�vX"�~%5�w2���|�z�IW���c�Շ��rX�3�Sx�G�bpzqi:��FɅ+�u,�#{�x����"�I������{�p��I�yF}����$N	�t;�!ct�jg؏�=�ڙL��6���x�Sb�X��	�ˀJ�_�Żl�(9%T�����le�7n����q��� �:�meo����������w|OD�79f�����5���6��,�Z>��f&�� ��zi�*�MI�.�#�w��m;p�B�d}l3�ې�:D�S�;����c���P�x��e�;@�p7�_3e�H��z�'b���ڛ��-�_��X-7�8η%�@�l�3=�ƾ�v*T{������fi�\���F<�G�zF:V�Q�8G�W[��E��uO�����������2���v�ya�xk��)�+l<�U�*��7�`�U�2��NN��$�&����vzb���䷅$@�V}��udt�}r�3aAY ����A�����9C瀱d�H�S�y� 2-�:6��Mon�#i� 4e=<��OA�Ṕj�!W ��v+ŌڄJtsW�"�Dß��&X��'���>���ߔ�q���%xK	9*��6e��;ٰ���v���H���:ؤMy��W!���Сb-�u���o�"�3UC�d��ل�Ds��̈��ff!��F[p��?�U�Լm��@�1P�y\?q=<���]��x1�He���~[�E�@?˱]�"���	������=/Ёِ[X���ɻ;��=j~p�1~�h��4��m��ʭY��#�n�ӥ��܊�G]?��.b��Y�J��������ʼ���E'� �G��U*�yj4{��[:�l]�'��i��k:G���"������V�KZ�r�ז��m]����-�2��+�уT��B#����ȩ��C{�}��^ ��V���z��'�21 �/#:0���~+��A�A�~Az�iR�_J�#ַ>E7Wn��#����ݸ� ��̖��N��[�w�N��ή��@2=�G�XN5��7���|S���>�T;����Mh##U����(L�̌G5%��D�� �<�
b�>^~��m�J6���pS�L���)�(6v���f0�}^�]Up���>T��N���禀���F�I�뀊�R�a�=i�#�\�s �EV�����&?��\����jy���#�v��_F�#�p6
������(�w@�+Fq>�}��c��~�����M�I)C&
�$��(Ӥ~�<�4��1y���d��jY�=�KA��!A�H#I?]���v�����gec�=�Tg��\�����Ue�!�LN!l�&I~�h����5��+�~�c8V��e�>VT����ak55RS�4#�Ž\Ρ�n��*��z���4x�DG��P������!b�\@�䀿�_O�Yf9�ܜ���s�Kuke�N��D�\S"PC�Yq��d�5X>ts���h�U���,ڛ�/Sg�Ml���U�y�*@6ɍ��������"_�*�LCA;��8咑 �5J8:��+t���'h�|۲�+�E~�R�W�?�L�:�|���Y»��Hl����k��$�~���fK�3t���S���W��7�o(��XӫX �,��,iI����F�
��(��οL�Ō˼�A�.�IZ��hm&�Q�(AML��z��a��b�%�e���<*�7�/�fk�~�g!4��ߩt6�t$]��k�I]l*Ԫ� �����5�0���H�*")as�_���Qᴻ���tRgq����OZ!�T-�#�F��J���Gp%�(h�X������3
PӨ��`��=�q�C#�(m_���i�M_žMxMp:��l��8�`��x�:s����U�t���JE��i�k+�g��6�w��;�lE����@w��h@��]����"-��ُ=�YɔR�|�z#�TR�P��y��I-���=�.-�)�s�l���J��ƣ�Z<��k�?8�M�?ر�4Tw6�S��_�h^&q%?�1,��,d�kCt��R��G_'=��y��D��X��C�-�����}qʩ�R��y��U�����?�Y[��H�������@M�͡j�d�>g�hS��\���5t$�1��{�!���g!�Zw���w�l��Ō���?h2��q�I!'��b��B�8Z43D��P�CW��<�]')Ԉi�4�,����[�MT��#*S~����#�����֡�&�\��a���w�W�I�S=�1}V�T�2#�����Yy��m�x]��k��'�#��&R������Wa,T��S����V@qc�U�oJ� ��Qi�]}qp�-YY	�ᷴr*���Fс'����"8�3�3�Z�-�_�|4�����*�BƆ���"ԧVe� �_[�X	�g5F�����[j�Xѱ���Hx�"!*{At��޶��b�-WN�(?��/�Sד��!e��(2jBq�<gU�7p��p)7�dU�v���<P�c&&'Ӵ�AT�K%�`�kB=�5F������;�w0OB�O�ce���$��fi����3�0�3�$���\���A�6�ང��0�z�3�0NA��Q7�w�'ۣ﹁&�|�$1�W&g[��`EOjy<���VQ����':{�fя�j��^E���k�ƹ����P�����!�5ӵo���/��u�9�SZ`J	q���m�zVN��j\r��:Ex#.è��}L�-�=3lkL�_#s��ֱOb�r���g��:�q��s^n���z7���_:	#�:� +��ND5z���h�I4}r�Ca�(�j�d8gE�k:ʹ�>��n^m�d�cľH�F>���_�Yo,��|�E�($�>��v]����6��,�Ր9�9��EM�X5��OisYsup:T�Q�U)����=�,���v��a	�M�]w&�`�HOІ�NUON�x������q"�����K$7���+sܚ3X�5�1���ѯ�*��R0�
e�lE�H�	!'1u�P*s�_�_�)�� �_�����W����}R��^D�p�˱:Uq�xڣ�&��
c�q����G�*ϱy��b/�D�;�`\����84�`HlӮKUY��
��|����nb���GӖ"j�ި�=6�P �_+/���������l;3���I�s��)�\Nt�*O�<WXd��ƕQ^4�Y�E�.m�YSKZ��w ��p���P��8��0�Ie�{��v�h&���D�\�ʃ��O�X8��dem韾#�Mh�a����g�s��Ϋ�����[�.Kj����	�m�f6&䶵:�AÄ��7�S�W��r]/�W��A�]"�J!	\��;��P�~�)��Ij���	9�N32�Rm�T���̐A0��`��}8Gx��L�p�4*o��P	�Ą\r�W	�?�x�ɽ mIQ����-w3��A���/�y18)J��}�*��pD�uŉ�������-������>���኉3�x>�v\C)��(Qe��/NA5Z���a�)�V*ݦ��&Rep��g�g�	���T�F����ƴ�bbAC8ҍ�|q
���:������4i��������Ƚ�[��?I��q0+^D� ���G\�)�臏�O��DO����結�~����!���yb_�!'K�1h�U��!S����Tm1�oS�6T@`�8V�q}!R4� 1 ���b�z2���6���:����RGh��D�j��q�%x)\��q�k��I0M�A��x{'��zF��ʰ`��o��{�r���S�%73��W�R�����������,�h)�_�E�&��a��a<��c��+���gP`\:+R�chB2�t$Y�ɦT�N�t�����W��"�C�2�&"H��d�uPKQ+!rf���>6.�+�U�na�my����vk�!�OC�ߍTA�]�����gI)y
z�d�;���_b��Z����P޶�L�1�TN�o��̪YZx	�#��o�0��+�~�H� �D��`gL��?�K�XS�O�n�'��"�T!!xj,�Ec*,��0�a��s6o
�!�p��w��ˑ�u`�>I�(�/�s4��E�=Q�iJR���"���R��8��3Z\�l�U%�Ǡw��r�o��C�q�v�O����ܷ�gk�c���a4K��kB��cp��Gd�=r__6��t�"/>BQ�8��� 8+D�b�<��?��p[��"�P��)�n�/t��X�~�y���px�k���s ���'Z�U}�9��~äZ@8Zc�Z����#'�r]$׆;�>x���W����~�.=�#J}��H:W?jթb4������Zt��� ~��A��U�*i�\��7,W|�y�B{-_E5k�	����tWNu�?�L����1�S�ʭ���O���+��j�}U��qS�G9P/ں�BIF-Z�aP5E��|�`5T���س�v1eQ>�yjȨ��>�L�Ĥ���\?� �-�n�`;�SF^�"V�A]��|��_�Cj3����nĜ�`�&БoMHb�HF�b�.a{��;���\d���uRʘ��F�U�I?�+@N�6w���.����8H��-rMh���\oe��o[f��(�G4��m\E~�N���eGCi�\���F�kf��`I��osKV�e��c�#�D��b(�4(��+ �a���*�U �yeɥ���k�:0ij;�x.K�qT�� ,*|4����m�t�{�T=��
��c;	h��<����
��H��h�{��#�����2����ҥ�N��V�7O-��ۊ7
���c�.p�U7{vk�gڤ8Bk������ Kz����7�"���Ʉ�7���0>9by��|7��AJ��&�V��c�w����~k��~�/��ˠw�L�
~����?{�E%���;C�ۅ;)>		ex��dufъ�Z�ֶ?��\����K�hQ|Nt�-EVH$�K&Mpq@.Y����CǾ��$g�1� Z�ɟ�͊�����-f&E7s������Ԅ�y��w;XA\�-=���r;�?�g�����F<�;s��ն
�� 聿g�kf�4/���0���"A�������b!'e���񩰌<�;`�Ovr�h�]t^co�����������T�l1�j�?;3z�#��3��PG��.~��tXH�5���=I���g;vc���7El��8�I�h	�j��H	��+\E!���.��J�0�)��"7�2N`����G|�U�
H������G����J��H΢���܃���lD���������-��8|�I�4���Q{��mN��7�Ӵ wQo{UT�Lee��OQL�z��f~TtK�S�D�`rh��.�����%�s��[g��)�"����7�mCsKHd�P{®�d�#B1�g�3��=@N�K�q�㜃���:J-�S$Y�́zP����.�`*qA��C�twC,����5��%z/^ .��nJs!S�u�tt��֜'�
V�m�<81IwsT���I�w�R���m-O+�2��������\�SR�Z�a\&W~.
�XNe? �y5���t׆⛂���mH�*.9��������E�`c	���IJ"?�N��7���A��3��'�d�T �\�;|n�@P�,��,�S��K���,	����9X*C����^C���c&~w:u4�
�\l���!��ڔ#Z��@*U��3��� :��f�r1��/)��0����v�h��G�����7M�[V�<�m�Vr{π�u����C7�p�JIT�l/m֐bs"�:���UN�v#5�F�8_g���6kI��Tf� �*�'���p��w7&(ډTtڼ�2��x�΄*�S<y��;`�s܀)����C�6t`,�J�#�����xm�$�AߟV�8��/;\��ÆeϨ6mŴ������&�Jg&��a'<�򔩷�x~��ȳKE�C��L�7
<�':�r"����hv"���sW��1RYG����\���[��������M���(�R��3�����B�'�ō�|%uQ�N�zuR{������	iwC�Y�@5S���t(̘O!|g�(΅ʢ.Y��Ao�����BM��kѮ>�<k�O<�H�j(��8�(a �'� ��A8F<Sp P�i�/�G�~8�~Hdא1=b������-���u�!�@;�fN�c��5!�J����+�4`}$�
����y6.N9���{��r{��<9��.x%�<��󹣢ޮ'Hz/b�vK��7�����_j#����8�q����td̿��w��lD����0"�u�Y
d��Rj*\A��5��I��3U�	�s�:|&\ꉮ���$�v��W�4��x��BD�@���X�k���vsR�ĽA$���k�tn"}��t��EdMJ�<$FX @����PJ4����Z#���$[�w����}�dh�X��&t��[�ɗэ�*Q�K�w�Y?<��`vlC�Wyo�@p2�G����_ ������8�������t���nœ�'�!����G������{E� 1��vY�pU4D�Y*o)أ��@���5�a�4��7DƆ�珢)gs�v����\ra��+gV�Ȱ������W�h?��r�5#N$�I� q�1����@2.�A���1�I�P/�6&��j���bNG�r���w�)y{^ .��>���W��*0%��P}�G��i�T��Q╖5��؍" �Ce��Z����K�/�R^DY�l�hFdo6#I���7\k��J٧�' R�5�*<xDk<2/;]�7�%,�5�ŉ��v� \�O��-m=����5UE�c��q��2�*���Q�
�P@1�DP�o�u�_��r,߳!hI@e�%ͅ ������f3e��	ľy,����X����4f�@�G�~�J�zq���1Sx/�oO����?�f
���inCfH%�z��zI_��UM�%j���VHљ����)*��� ~L[�)��0[ZSwH���F������<�pm�L�1f���"�^x�C�J��QuNi�#M�5�i���Fɱ�F�J�k��)�`��E�����?ɖ!g8�yN��8�@�.�Ӛ�zc>�� J�� vK��Rv�y�dv��dk���[� �kD�n�h�z�w@���u���z���p�v^9�w/��yRF�A���<m&���A^���9S���RIg�ؐ\������^�yT���O������!���4/=o��A�r�Ia����ܛ��T	&W3���ۦ.%���/��{!H�^�]�	��,�ʌ�t�U6���wbC��Z(�wNh%H��W�+�k�"�m�����c���GG�g�  m vt/F#?	\�'�A�f�l�d�H�t9a&�m ������A���N����d�=��_�gy�q�z�M��(� B�R`�Y�,�8]^�,n�2�Ǆ�%ލ�����j�1�a���E��Vki-Oj��K6o�*���u��VS c��ȩ�m���b`��e��9�~?=���u�ǬA�t�3J�u�������dUꅀ�� ���P��A4�Œ��/V*A�"�o�߆�=�S�Ylz%$�;��f����M�+�'m�mX�;��]�6�Y� �]�?m[�ߎZ�=�D���=4��{I�{�t]��+d��/M��I��B����\��yX�>� �z�'���>���Y���@u�7I87��d �sy濼a����-m�r�m�"a�$^j�ɜU�Y,f�_��,��4��O�ؐ]7�4d4�
ᖪS�gKW1�ʨZx����`Z��8>߿����n�|V��8뼮Z��ɮ�>$��^#�
�����U�I�ʵyw���cv<�7^w�C��BA�J[ݴ�j�+E���^�E��|�%�M��^�8N�����%�l�k�w҆����s�T2E�;��77��t��Ř{���'3A�&
!2�~pK9Y��m@���)�8b���|&ԙ�:��tEO{f��*_��#�K#�@�J�HK�a݀urJR�hU�}.���#���c�H(s�Ӓ�JP�c@M-�J���F$��)K��W��ڵ�j&�N[�E���ye�������o��Z8��$x��a��cl��k#.���Fz/�&O�o�SW��dc(g�,`�X]KD]��e�\��j�&�'�uO��C�������_�����)�.I�O���u��%�����×��_d���� �3�o?��Bw��I@��4���Jܟ�"����~��Ŋ�N��e}�z�!���.���B>�Ր�n3e�݄[� ���-�������bQ��|�샄����l�H
�im�o��"vrtT���u�.�u�c�G6-Z���ā}��_/�]��� 8]�*f�m�~g�bG/=�T<�O�ŞM(F���z��*�%����` ��y��y��R��Y%Y�C7�ݶ�u�n��a�g\��)�P���wv�����ŷ��B��@�����mH��#�l��q  ˔�$r	��ݳ�5�;x�'�1A�)D Žh�e�X����>�K��D?g�g��u2!���v�R���C_��B�/��8n�w�
ĪcF�?�oSc@S�	�������@_ap�������k�J���k�=���ݥPIs��#pЃL��A�z6�v��'��@$������zj�g�>h�,��u�刊Q�J���)ў����m�ڵQ��x�S1���8` &Ŧ-`W�e���{C�0Z#ZѦݝ4��WOَP�D{��]�-(U�J��:����F�:3��.U�	��2����N�;��Y^=�e"����u��eu�^����r�P�H�.�q�Ȇ�\�;R������6=>�q�F�=]b�h��n�w�C�>م.��`�c��#�����q2,����=���F��>=ԖE!�=7���2e���ʘc�
4X����6y?�P#. �4{��8Q�FU%���{xȹ�+F��o߅����f�Z����j�t��!�U�f��Z�I?OB�iN�=�B��Z�:��ٞ�1�qF�5�՞*1�JT��F��j��!Bx^N��/��bV�n��1&���"���b�R���O��(I��G�4z-��Cu��ūV�(*X�����fc�C�)����ŮCy�^7�2*��|�G��m"�6���ʆ���\ze��9)��O"���}3xE��
�~�Q�Z�G�E�Ћ�d) ����?|���@�s�b�-�Я�-�V��VT����H�V����'�>{Y����i�gs�K#gHw���{��m�S��!�D)���3Dy����
�����s!����K�ȣQ�xǜ�gR2��e��ւV�Ў�߂'-��D�S�@]��;b@5���ׂ�~gHm�d�W,!���W4�=��������r�*u�"����2�yZ�h�}�ɣ���.��f�+�9VH��ǧG�׉�s;�kz�xC�� ����u��7�;��Z~&����W����Y��O�W�B1��)�����~g�"��h��O&� �.\<���8�Z��L��+^
ua#�h�)Ka�גڅ�S���[�gdU5C����f�z�]�?&#ӗa��l'����e둇��8�:�cD4�d&��z$��G��^h��K�X�7�N��'�"��}-�<bU��=���p��d4��R@�.R3C��/S�L���I(u��bND;����:E�E ��{.Z�� �9���^��D�U��UP�8���3=�2������\��j0���k���!�g��i��3�h��81'��3e,k5[nXu������r��\�N]�B�g��^aazVc]p���s��A�|�g��90OT�� �����^|< ����D5'�wX���ՆVϥ�i�qpM��4�D�8�}�/]���/A���Җ�hbs�(�J;����l�D_c�8���[5��O�š��^��n�h�0i�MλՑ���o���\�G�hd[y_��>F�q��akb��zS$Ş�?�����r�J��scb�����5�1e�hLM�����_���o}#\�th&m�SC#Q��Bt�˼�.�I�� T�liw��K[�r`�2ٝ�uB"�tߜ��o98{�ᾖ�D�9�/�N�_����\�b�iV:b|�%�֭��d~Os�#�s��k�bl,�[�����z��wsA��Q�ۄ��-wY8*zeA` �6�_�(k^��}��#Eq�k��1�$
�«&Zw��dc%�l�L�B�mUr��v/C\ĭ��&�;a}�Z�%Q+H������y�j�*N������2��O��e�F?PKVA�v�M�]�z��E��^j ��N�veB��+�� >�m�"}�f^@�zb�2�}je-;�8eƸ.ۿSx�iD	�ja�����=��S�s�{e3�⯅�����d+A��yXn�xn*#�`����W�3hV��2b����YO:�v?��v��'�B7^��
vi�V(*�v���b����uEx���IR�R���@n)��*�����]��vLp^�=1h�J�E���!2��y*�����@��ϐ��n����-���n'q�p������x�ҡϰI�A���gD��R��82�vznN�#g3��A1];���.}2��L����d;�r�����lT��}x{�����ԝS�m0�sG-�����i@�&��n����o�����Bg���x���x�4�g��(;�ı��-����/p G\�ua�w�����,���A�@,V'�]Z�^��-�R�n��r���[5�����[�:�-ˤ;Z��1^���ץq���#2*�"yR���i�����S�'�#ܸM��g�?�w�50��Δ�ͪ����&fB�ī?x�k,���
�\_��K@�~Ƽ��੺��dh�2<B�?A<nw���@*��h6l��k�m��inT���}�����4Ɋub���#����.�h��ɴ�{���a~�w��gN��?+c��������l�	Z��v;~*��"Zd)����vK���.�����d�̘8�������`�� nV�i��+�S\;�h(�$J/����&@w(� �����L�qX��-��g�v�5_���HK��aNP�}d�v��I"��ӇG�+�f<��x���g�+N�:�����S+�3�	�Pd�ŹɪR��?	�� 
j���W'
�� �x�
<�����'җn<8��F�[��S+,s8U�׃`ŋԌ��,_�6��Js���OW��_�L&��j��PmjYY�P7B��os���nT���J����V;p�������sS��(��y h��c&>5=L�B��l6's+67���8q�.�M�}����QzJ�p�Q�KC�Qd���i|�ǒ���DP�����
NK:� ~5jNk���&G"e��z�����?�o��i�T��cdB��8�K�0�)�`�[p����nz��U�8ׅ�{f�?�*/�L W���&7%��k�#az]X��3U�aᎾ>�*�<a�x�L�B�GJ��d;��t���6�:}�Zl!�B��܃ޝd!AZ�D��Xk��?�5�O�Π+0^���ë�=KI �ZG�9u��OڻZ#�\Y���KR���=mOyM1Lǲ�}��Jhg���?�.�
?H򼜇)0�_B껒4�&1���B���b�/��O�\���Xo�(���P ��
5���=8��b�\�P7#�m�)���%�
0�����M�C�l+r�
i���ڗ	'�_ڨШ�3�(�ʟjx&��h3z�v-q�v��u��Vl0�n5fF�%�!��LL�j�]?�v��(�}�� jxS�Q)ӟKy�t�Ykw�],��/"�D����u�;��K���E�	�b���}�R�����o���_d�衮�Hy�n�PYn08�Jt?VC��Ȱ3�
�R�`�
%�xpT`���� "O���'�)�h�����jL�C�
��fʳ����^
k�׳Fԏbj�Ũ#z9��W.��		�2�Pz�}♆.�Ņ����Ȏ�s�l��b��Q�A�
��<��[��*B�Uma�nw�� o��q��f�/}!P[i ���BU�y=�-�a�~9���oE�ҽ�]nϷ�t�:XBxCJAަ6��]٣R�gX~��Di�A��a�Puމ�X�V-@�9�t��w�O��ךn|͕ǷW�c��(��E���Ŧ�%יZ����*�.��������Yh�і笥�_rj&H��ϥ���G�vdLL8��{��<o�f��,c��z������o�s�����#��<x�ԁ�g@ܐ�r})t�V>C3����|���I9�-���,�o����hޔ/��)Z�*6K�n�m^�)tPc��S�qe�b�?6M�YI�t��ƗQ�ҿ���0I~�I��,n�����Vfr�$�p��X�7S=�'/�k�>V�_�Y�ELsv7�=�0�Ը��ИM�^��ID1�l����6���w�?�#NQl�h`�?���^��VA?���>�y�5�*i�B�� p��tu�j�"�ꅟI��b�6[;���!+k��H�:��צ$pKL�B��,6�/ �p�����F�ly�32d��x�P)�v]���<y���l�.]�- �;V�%������}9�B�΍�}�P���o��k��>��U���C�0�B��s]�T��z>2�;׾�z�g���A��#୚�}����:��Jes>�g7��x����m�Ǌ��p�q�,d�3��{ [	�����a�|�0"��O�����<ӖF�S���	NU�e��NK�˨���~GB���m��Gź�8�����J;;�ZS��ff�;7�ѱ�ֺ��k��FnV��� NR��wzOQ�ްE,�Ct�J1V�_c���j3�2��t�y�=S�X8j�X����u���]�p�k+(�o�=4���B��ʠ���+67���וxbׇ0[���,��؊��ՠ��˾��JJ �ll�ŭ�>��l�c��P�j�|��-Ig�<��Z�X3�����aM�M�-F�i�Y�L�6���m������zу��ǯt6%&bRaw���O7���԰i=��Ԫ�m�@���n����w�7k����uS�E��#H�����sY(Ȍ�U�Nt����)���B��� T϶�#u/���Y�1��2\���qX�єtH�����*M���������%��kލ���W+xʜͺk�
3�T+y@����*u���U!��,rz3�(�#�UR8E���?}ܙ�(k*� ��.�-�ھ��(�����(qe�<���~��e���h����¶N�a��Kϓl&8��\�d.59��B��=�z蠝w8�������������:�]s��C"��0��A;bb�Nx����QsY��"Z������Г"/I�C�:���R�I�$:Z�Z.��Y�MN�N_5��S��g�W�I���4C�`������0�G���\�z�At��4У.6ޖ�M���=�V�́��\_<9���E��`����!�99�;[����7���lw]�v����^bt��S�LYx��x�lkL�QJ=�}����r��BA2�h���c�N����	'�#����w{�v��a[��Oջ�d��R)Җ��zp�N�����W�N�Ap�v���o@����8,���=y�P]�R���F��X�w�D������5�45Nv{ޡ�	�eVK(�ʞ���|ev�~U!�|[j!#΋2t7M�/�^'Y0�����p&���6T��3b!N�ۡ'L$�؄��'��5S��C�T���B!Ork�95!�i�ɚ��2��ea���*%�x'�Pf��Z�^Y0GS��H�r���u/Ao��Ze�&���w����I32��R6�� ~Ӱ1᧰����y28��e��$�}�b��-��L�H��{�0aC�+9�{k�ل	i�"��Z�w�x��%�;�ץ�r�j3f���j��""'��0n�C�#�����	��uM���[2��֞@0�J:�,�ZQ�8|��*Wv��Ԕ�:��@�-X�a���� n����ЧEAtz��c�&\2���R���+K��+{Az�Y-�q@���uH����: ^��5�_��4�� ��Y�!)��_�Peyf�s��o���£ʂx�3��)������m�ԗc�K}��	�:.��^٨��z��\�e<���(5��ē���@�j���@
X�}��U|��������1<~T>���,r�Z���W��+okp�j����O:���'�eC�}�ӟ�[14�����Wᄺ��dC9�/<�PSp�˘%NS0�/*?�_����-���]+v�b֛Xk���Gr���A���֒D��sFj��),Tk��U�����gD�~�h���К��	]v������}d��o0p�GL�������]T���f���)j_�M���%������6	`/�����v�[�cӇJ/�*�"F!�0���i��ǭ �s��;�dÿ;��`0��G��c�<y�&�!��6�RT���!=���xH�������O�D~�L�N�y�`5�>���4�rH�� ܧ��9��E,�#���->�7A��׌��E�L(�}�K�O�aM�~�8%�=@�o��o����9�{qk=gi5��c�.�&�H�.y�8U������-�b��M����tU��N��M�T=��|�J,P_`�Q��ξ�R��t�Z�Z��)Rmi�t���C*��(=�� 2qBx�|*;,֮v26�oDu�3-����6G6V;��K�w�o�$�͓����(#�|e�q����7 �HɁ���z%����#pG���Ald7HH{�e�'��F@ +Τ�����H��W0x	O�_x��"^0i��}��BmLF��Y~��2�����r�9b�Go)l�L%eE>YN��pynK����\�8�!�Dr����ą��gj�c��F����N�7]cgi�e9�H���Ǻ5�=&�Hx򱰊15&�Q!�n�.��zJ�) #��V�>�d�i?%�ei_!�݀Y�汰�3ͫ����	l��)��:��б-O*��*�DW������E��l^z9�9xi�_����Ed7X�Pm�T7�Y$=�,��H�R��T���8��ܗ^Mh��i�C�a�b�@n���Yp_˱6����c�k�6B�?2���
�X�"x�����|DJ�	Eǲ0s�
u)�a�p���� K/GÞ�� )��P��g���\&I�?��IhE�����E�_3���&2kSL��� B=�ˡ��~�A����s΀.�����I��I?�Ԫ‑+X%��~����j����- �?ֆ�8/�H�����2U�&��F9��+�)Z�,��uq�)9��;"�'��y��E�<�X��!��콍z~QF�h�"O�@N8���Fmm,�U�p��rl1!Z]����@��ley~x�!��H�-!�_��2��	ٜJ�@O����k�B�����F�W�Χ"
]�ΥU��PV���}���&_�qRR�d����J��E�$��:�ᚩٕy����Q̡Y1��(3߉$o��*��Ƹ^�zz\�}D5%��Z�M����a��LD����Ƃ��𩛘���%7Z�Xw����=��Y[ߪ�ڻ� �Gv�:~�������@<�8��8s��+��=t�����}� ��k�[Z" d�/��%n����ؠ;"�,'1�>�;"���/8�RWUq��!X����)�^R?��b��7O��Y�%��c��s���N��'��]� ��7!�� ��Dgp��P�A4Nj0K�E�����ݐ<D��~�^
Ȓ��P��[�[&R�,Z
(\����0����3�'TWgi�b�pL�3�����·��q�Fx�*�E&&C�:��"�$�yC7��8~;	��ʹ�4;�@�~���,�'?��M��)8����2�l���������>���CJMge�}�T�J�߲T��ۻ���I������ǂ@�7�Α�(^�G��ߦV��Yck�`l�1�ڀ�����/;��) .?�F�[�.a˦|o'G��3�~�t��|��ӿ��R�]ޚgLon}XX���S�6����f�8d�<�`�rA`�:W��4g�frG��h!,��h���%�$3P��)#�n��;��;������7�h�In��uz�mo�K�=l�m�M�6:�ڀ��S�U��x��D�L�������%j�0z�p�h`�T�n�6wl8��eݹ"s�e���m�!�-��[�cT6#�`�49Q�&l�"�=g��z�v��a����ʬ��-�d��RK���.����to�oP��� %�
��
�,����Rԅ�W�R�?u�?&�+ZŽCR�����TX��&���1�jFdJ�Yzɣ���a;4쫋{o��('���r��a��^}�{�l�[����5��-Ze��^07� e���� �u����ۃ���ak��\n
t�Z9�t������3bVc�R>���sP�0B�H,�@��0���,�$+XS��uv���L^��LV%)^���L�'����&�)T6;���>��n\��B!���B�����yJW�E�����R|7�h@�V+1��C��I;��P���=���[|B���e.�̏Ӓ~��#��6���~-׸;��Y�hA�M�J�D���Q<�9�Q�w���b��c�pG��Y�w��g(�V���z�T�E;Q��j�ć��q5�k5�4�)@�'�4D=t�2���o�[�#[��`�4�@���96�Ks�#�W����	�O~4L�E��iћn_Te,)�ίC��o�:U���ߖ�i�ƪGj�[��{�Y<��4�A�H�
vb+�Ae���N*�г�M]d�H�9X��.B��8���;@�ї������p�'v�8�#�D@�����x�h����go�Ϣ5VC2)�E��7G��<���a�>����I�բ�)�P�$m5�&���#�b�^R9��Rb�3ס�g��'sb=9c���	P+��wI��8�):�e�$�%�A)�J{T|������>]��w�h(�l���G99i'�����h�o���"�5�%r���;�[�`��.�S?�4��-LSp���z ���FZ��;�椀��9�,�N�暡Qs���Q{\��?j��h� �p53�1r�������C�
5ZL�a�bR��d\vZˑ�W�4V�|#'��eB&Y��l|�᷻dp�jGM+��)�h��v�iw��B.�H�7�� 'ϧ��x�x�U�E(�@>�/����K�b� ʏ�@���xeh&����Ⱦ@2����!��JA�q��#�}��n�o
e�+9Ȍ�0�7����pxdR���trC:`Ђ��V�ح�#��wDjŷ'/��y�J��ačkdlZA؉N�v�sL���Y�Kʭ�㔿��2U;��ؔ���[4�����8��Ad8z��M�q9�u��_F}���{aɁrM.7����7��n�Q�y}�aJXlHI�k�S;�ym᜜Nx���	ݮh�H��S�Ԑר���.W^�@N��)W	�:XT������(���@����k��F8��M|�=�S��ND�D���&�ɆX�"����"0�)�o���������K6wu�]0>ɚ�8�X�SI��v$��������3 �X�B\ɝ?�,�c�QV�G��48���,q�����.f��&4���r��_t{ ��2��vo��W˚�g��(m2�V'*X��T���:��F���ђ>��f�����]Z����ߝҺ���'���%��"B.q�ty�NN���R"��M�����D��5i4*��y�%�~�T(y�'���?��^�v}�3	:�u	���ʛ2�I�X�%[ �k��tN�i�$c�1ؑm�GCL���30��R;  i��!5���r�b���mhF/�i�� ܊��k{��ڹ��U����9�tR�l��7n%���q��D���Ŭ� �xd������!�;!��J����@���|G("�''�� ;ڿ1�f5 �
�m��C��B=�|�<���K�XT�أ��]�����d���5ݝ@�G{}�-2��|�(���OR���bq ���[�|�w��#�O�t:�V$���7��c�65�He���Q?r��		�z��+Ӕ�	���X��
_b7�PD����A`�Bq_ލ�A}�>�.�a�~�D��toeE3���%��س�ۛ�B�b8�Fp�RU]�E�\h�L�����8$���
)�G�Q��o�~�ā<b;)#�)T*�Ӻ#��࠳�x��Sq��2�t���롐���D �o0ce���r������:�x 5{Ę6��P�6����s,��F$x�zN��-�^��	�]�����"k�f"9
�w'5�\�֠��kbf�p�h5�7�Б>	�F �L�ݽ����4v��=e3$�4HK�S����ֹj�qF��3�����z����rv�B��1>��-(F�D`�uj��p��LC����aF�w7��|LH�*E���F�&,�O*]��^�Iľ���k���s�Q=��Y��y�L������o�E}0䚋-m �G��m�O�|65�#����峕�/d�)kXS�Y�\��o�Iˬ-��iyQ8���C�!��Sه? ^_�A5���� [��x�?�ĚTq`E�l�˺����t��\�ko���EiO;F�MC��=�!n������}�+�&pk����s����5	��T bk;��$dix�(���u���A�pdƵϡU&EQ����gQ�u6cڦ���̮����1��*5��]\	�O���n13�]|ࣦA�D�o0�&j�k1����H�u��n>qɡSY�ܣ��.�G�r�YQM�/�[MRY�b:A�|SM}��������A�l�1����Zx�W�08�R�x�]�mr(x۳!Z����5��q|1��M=���^|=S��'߉�ƶ(k"����f,7����TJ��>#��=Ԁ�e\v'ɗ��� `���H�����:��	j�S-���~1qdZ��[�=�B�4���3�4ٵ^�υs�翹~��_�f��+2��>u��0��;W���Du����3Lvd:L�3�/��ka��p"ٗ8�N��*�̋���g	���J��M���b�%�����ц5�,M�4-�7EI� ������\�K{��Z�8aK�P��d�qu��2��&LS&��E
�薘Vm�u_~��C����L��b��@��ɇ |���(�9�5�dNNdh�a�4����0r�2�g's��Q����5PQ�^��`)i�ѿy��{-.<����Ip��"5�,#N� �
��0k�� ؒ�m�Sks8�E}�ݍ��S�=m�9����׽��c�����An:7=ۭM�!�ذ܌�9I�=s�C�X#����	g�Ψ�j&U��q~6$:*?�*��B� �ʒPr�Er��^2�2�?/kx|��$�#�l�F-���1(L@�Cg�D���I'�@����D�����JW���:'Ǭ�fV,�����0;��1�e��-��'��z���2[�>uV9�ch��>�ǌW�qQ}X�p�M�e�v�����V���"�$�/t�m�5ղ_����w��.�1��
J�PսX�1�μ/�.!g��$�m6j�3.�;2L��,7�'EҞ�ރ*Q�J�WM:v�Wu(���"�'{tS��?��g�ك���\L"�?n�@�=M�M�m�L�o���3L@��_�;u��S*ִ�QX�go��=�R�^�ub/�(�����])n��4>���0u�~�֡���Řx�yr�(@��,��k����䙚����HH�̓%H�o:��I������.UQt2����S�y�E��Qw��'a'�j��-U��~lU�Ik�lo��xՀn�ޏ�t���R���[�?Ϥ����~����uG��<?������Yz�zwx�e'�0e���E�$!��
�R:�g��^� �)�sU����"�i��3K�������f�x7h��pn1�W���z�sz�ŝWB7����7YŇ����	
�=���fCT�#�8Z﬿�*O��,�x4Yj�HN�u�i�5=�F�Ȗ�瘈��>p9��׉g��l���0��e�X8�J�U�0#!�*�^��&a��͔��-m�WKi}F�ǥ��؄[Icض]��/py������'��_����n��E4<л����������ןx�d�=	�ˈk$vU!���r�t
�?u�޹���H�-L����0�hpbk�M|8�8q��7@�6Ӄ�;fV~��GՆ? @�����w����%�g��FD�.���o�ՠ��>JinZ�j��%��|��:O[K��C�8�6�(@������UPG��v����g4d��E}�����.S��o6u>3�5��I�l�`����߉��Uقۀ��v��AӾ�fY��A��ed��(�x̍�r~<
&{��?>	|��]����7��t�iaǵy�J�u,!����r��[=��31�O��^�r�3x�S��}eh�rkti�R�}l_*��}W+}�����)6�;��5Ly���j���`7�AjS���$ɶ�oڭ�Ra<����+�l.��K��O��D*�O�d�0. ��s4� *�{Y�D1�GH��ju�3�ZL�Ɂ�9��mv6Z$��jR�w�E�b܌VX�Ⱦ�C8oZ�oba!�݉�j�7vh��^N���)�0߫U �/���~Ŋt;6�?�]��Y�[�(��
7�FD�/�yxH=Q�WR��:<$N[��L@�r��e���&U_�?26�v��@�<���0�C�(�8��ZW�c��I�k�^�U�Rf��f���f;ӱ�_?GEքI[I���Jxrq5m��f��ji
�c+�U���aUi�U��M1��0+�4���-��c]���3�G������k�d<�����Ƿ�k^RS�(�6��1�=M����#�r#���8��nA���]�����,��ԛ��o��a���xʺTP~8 ]$�ξ�1�6W`�4ݓip0<����?�v��u�<�ͫ�b�ܠ�
���6�u��뎿���yJ��=�O�Q�ƣ��x���}����z�h�����i�6�a��'{�a a�I��辠�	���N�Csv�_��$Sb�5���_���e�y�q�� �`�2ᵪX@��n�Ԭh2{c�;�M�������`�'(�ev�����G-|�%�L��U��#Z2��D�Nޢ��:<nW��H���Kk��4�Ê�K�7����R��e�u
娛Z��n�OQ�U�Gv�z��,�:�1�4��j���-D�������KF����$ ���v[I��P��D#�	�o��$
w�7^[���U|U@V ����t��m~�G{ve}�y�*�}9 ε*��1�11k�!��9��&��_xw���}�܉��ǲ�D5��G{6�ը�z��OO��H8J7�sL���s��' j.�5ǟ`+���k5/�[�TxNչ�jR���NVU��б��9����9�6*�c3�������"�+E�M�I��ż����KR)I\���"P���sI$ֹ�Nt:���5��,����\r�P	���
�5��he|gT@�D�,O�f�S+בdui�Oh���70!���_�_����c�ŉ�1�AO�I��a������1|�T��~������	?�G���Ifz�[}\$��>�\E