��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���}AW��l��&�zZ�#F����e�i��j*�z\����1��8qvY�������B��
�>cs�I 4W<��m��#L�&���
�t�j���i���n��5�9����X2c`�|_}�h�
_��K��JG��b���fq��z3�H{ΘIm��>�$��E�Z\�w����Bt�?����%e���x����Y]PI��W+!�9gxђ}>��;㡨 �l�o��/�=�3�o��Eq}�e��2�PW�a�u�>.�7�����f��o�G�b
o�I9�ǾU¿t�YV��=�[3v$�a����xT�u �;lK2�(����$��
C�d�9��t ��K�m���wb�p��� >e�ݳvv�H�sh�bks�/�3t�D�Q�rк�3�Rz���xtx]�g�$coTf�>��E�����_�%D}ڟ�E(�N���1A0��P�Aô�d�3l�i����u��o��)��{��Z�3�H��Z�4������Aͼ}���3Jh�G�ɱ���?(+�,E�:����j�&Ud���J<��R���峄�ǌ�7a1�Ƚ#���c�0��U�Y�-����O8��6�a��yN^\��|]���0���pO�\?��W�ȃ�yiP'�(���ߟ�n��[f����Q|����?�j��F ��a��%&�~���0$!�,�� )��o�R>����acv��\3�q��������=�f?��az'Q��	����5\��?�G������m�T�~�__X"A_u�,�`H�fp[��p4�A�����p/�
<���O��T��&�]��V����w�Za&Ǧ=��R���/���
�z�<���X)��ˡu�`O��~��B�W2ީ�꯿)
a�� F�HA 8S���B�t�TlU�ۜ\Ϸ�o�U�7+��_PH�C����w�����r������&N?5�wҾ��٫vl���A֊k	�����t61�$}�V�>NX�ڈ�&G����BRI}��ۘ!3�>i$��C��fH*��bT��oq��*�Ө��0#��f���p%�Z�2�J�ڃ2��X�m��׮��G����8c�!S�`	Z�t 6�ڟ0b>�.��N'X�űÇ���"g�lH�����Am?���l׋7��>�m?W�S<	��a�WBs�Mj��e~�d���4Φ��s�Xx�;��3A٭�m���<H
��8���9�F���[v*�p�;�)k�Z.đO��2�!�.�}pN���)�i�۩�yg�ޥ$����d�Ӓ������E�EwU��c��:EN���T�+n�V��3N��z��ga�7c��F��)E��"`�NUk�B� w2�Wޠ0��
��۴��a-fWOҝ�Z�J�(�Y����vC�yJ��� <N��)�2�$4��-H�� L��N=@s��0`9장_7��@5^�m������-���.nYYV��X�`�٥L�gV����ŉ.�ߟ���X�w�6.��.➩�����>y^�**b��6;��Cn�Ł��
K���X�g���u�1�FV#��)�Ls��ҷ��HA�ޒq#Ԩt��*�XA�3�r3�t?�@��Zъ�`
2�,�@��:�D#Q7��.�|��\�ӣ+>�Mk�h�Vn��A��b2���t������.����d��4륿��~_�ڶE���?]ê�G�����L��j1{V5W5�,���;��n����L���M�����s����:	�2�F&���)��GR���Ku/����ϠX���1i�ɰ$^�9��v��s�`�(pip��}�楋E �GL�Z̖�t��8՜�=��~ѩ.P8w.*��g��4�HbZn����x�j8O|E��|����S���]�b%S���`|n��鸰�z���j|�����_�[P�
.��6���y�n-�/��I��	���*�2�YM�^�����ryG`�Z^�>�6dc����M�Ok�Ҁ+eְ�=��I�p� �)�wֶ���'�O�}��*�Y�#���އ�Ѐ���c�U��թ���sK�^��j���{[���"�o9P��䒹����_3FAJ�}?Y>�