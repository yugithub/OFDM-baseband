��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ��t-�Y�n�.>�!ɸ��r��a,��x��h]�����1�g}_?	xm�
�f���yG�)���H�^���Y(����&�!�&#i�ţ��YaÈ6��r���^��()	C����O�B��N�k��XRS��-�*�~j�������H�_�"��k�����c��妢Jm�]l�4�Ne�"ů ��," /^��f�e�D���>2�F��_���ӇQ*����[ż��BԈ��5f�@	��A��F=g�[^�� ��Z���$�����\5�}e]Cs[�UQ����~���	L"��	��.��_z�+1����=JTv~�L�/��t�e��(�;,`�t7n,��U�w)�P7PX�u_�f�%�����[���e�L�V��u���f�����x�x�_�~]�di�|��Ǫа��R��
	�t>��	�6
��t����>QF��ܷ���cV-��@f,h|[\��F��ױ�����){I�Л�E>�|:-�>��=�0�}D��PLE���B�e&֓jǖ��R��۷R��(ױƯ�K�K>ܩ�z�	;�"y�9>М,L��0��J���y�6���B{?������j�Yr��"������4
���oĖ�_�޳'��_�e��aN]�m��eJ�;��ҨyZw���x 0���C��W �� ���dx�q��s�$�ވ5��.��O]�m!�4�Q�W� ;K��`�'9kg�o���ra8�}t� S���| &����E�@�x�yZ�ݏ�=a|�"ַa� O�]�����;�������w��%`�
F�N]�r1��҉�|ڡ�s�ݐ�G���5�!�B\=��C��[j��$+{�"C���4K����MqS���`I��V�ɨw��_����g��e<n�s�b��_�Է_\�����XǱ�%ɶ��G�p�.��/��F��E*<�f��k@����[��[�D��kW�q�zx�$j 	��`,�P���P6����PR��M��V�3J����g"�8����V.����_H	ܺ(��7��l2R��P�&8D<�[�����6��$I������z�? N��o�0�0�3�0���o��wxҾ�o�Kl��ml�@� ��S F����ڰ2;�o"ci6�#� ������쁘�>���J�p�������\����a�y�?���W�#� D��7,
�KA�/¶���!3���r\x��o�A�y�("�-uNV�t�{����vI�TX(9!�38��3x������!�7(�2O�U3vq�����n���l�w	q,�9�퓛��^[M��-���`�Qr5��a�Wm�cy�����s)�Mxb�zg��/���?S��h͋H��l�ϡ�`���
FF��q�-/����jb�l���)���o�26-�E��~�xrj��������O\쬿�8��<͈9fu]k|������w�2I.��c��/���>.�9��G�M�	�8�w ��Cڕ�Z�se6�?.
|���	��,��9��D��&��ɳ�W.��6|ײ�tD8:A��K7�A�"tϫ�`��OOc��y�Lɛll�B�b�������d��0-ή�{vC'%c-�gf���/���	,|V9���Ώ���d�|v�]��yU�''�;&�7)v�	X�i�w�/�4l������_��1e�N��¥o���H3�KwF;@����7� G��b��`;�a%{CHC�Sr���f%9'�_GPH��YD��:q����T��q��M���zr06��v��lZ�fb�694{�u־��T���N�SC8h-�J���-د K��	��5�)@l�cMax��n���^���a�j����^��'l%���>h:����C �%����N��`Q6,eVHG�I'[��y�I��� 1X�O��ʃ&ZR2ա��a�L���@�zs��W���d�׶Tv$
r�2�#{?������SM�7�A`�y֤Ü�+Bs�^�(j��1%H��~|� �k��V��B��I�D�q���!���ψ�����_��v����~��5���iY�^��;]5 C��y�2]��p
����H3��`�.�4���,��Ъuz;��8����\'���V!x,�[�'��v���4g��J���>�k�⥐O&C3��b[e���G�l�i�~�kZ@424OD-���%�������F/z����;����!E!7�V́��)uԵ�(�t&E9��B�����a�,��(Y"���@E��X�q���.�	؁�����d��m���@j�RQ{�/jλ�y��<�8�MTh+k��ےKs?�u�|	�Z1���
=�\*ƣ�J�s�|�%�zo���R��N�������Y70N�6"ߐ�_s�|�������`�i�R���9 �HVC�ỏ�ۊw$�a]����Јȉ�bY�/>��`Xi2�O�mcq�rG�������a�!|���+��̡����"��ൎB��ؓ� /��9D_9:��Ahbyz,r��{nG fA�B2�����z�snT<[���nP�o	g�.�������6��,���SL:�2�3p#�R�\�����M�![{��y�/b�1%T�S�(Eo���s{*$$�M�����)IVv+��ݔ�
�bQ����l �����,i]�J�"�&Ws2)�n�t�Δ(��u���1�.T4��?w)h�~A�>G�j�d����'�·�(*��#��m��6V1g������k^/��`Yz6��0�7�'��J-�D�I��2~���\&g��Y���������!2�f�e�Obk�3�:G�MC�$^����T��6���;�����`�%0�
��{p
��v�����ͿV�Kx�B�/�H�;Y��Uu��֒֡F@<���a���Z���=�������x���9���x�����Kj0\�/:8�ݎ�))�b�IS(M{(����%�O��༠�-f��/�V��:O�v���]/�䛑�/��/�9�vR��6Y��.���7�G���N��ї p���B+��YP^��7q��S���b�)�|�<��{w��D�_�aTtSځ�ɭm�zS/���bq'�|���2 �>)���G��5�����i�uŷ��m;E�v9 :A̏|�Z��CMy{t�x���=��c3��p��j�e`C�̂f� �\<�����R��Y�3��[�9J��J �{Z�#��@�p�JM�+��s;���;ɨ,t��k>�K>�W9��~�M��Ӡ�����x�9�C�l.xh7���0����y̍-��3�n<ޣE ޺��٨Cw�aW��N��FEN�Q��0���!n#���X�y]�gw71!��;��a��CG�n�*���|��+Ma�|��ļŷ�9��d�sE��&b=��ٜA�(�P ��5��b9�~��E����z\dh~�WΧ`��4A|�n$�������k{M!ZbO��`�;k�4�&�����`��P���5`GP�ݑB>�TC��.Q�_�_�7�@G7'�y���m�l����y�lњĔ�����H��7�~i&$��������U/�.&?Sor��U&Z�����n����>���E�r���$����&࿼��q�N��y�ٵ�F�Ê�����A�挂���r���$��N�����27�Z��\C�Z�c:��Q?�����e������WH���a]7ޓ��œB�.�(��Z�=�ߎ�B�,Ͻ�N( wFt��G���vt�������o����(�S�ff�|�p^!Ax��P�^ܩ�A}��-MF+ �a>�\����.���	=O�i�=��V�.ZE��j�	�)�-�SFRwDm��Yiu0��p	�R���ǷX>%�]@�Rk���f��"Oz-���.�� ��\�wg��0\v�_јͯ�]��Oچ�������oW���W2VU~ڡ�Ól���$������@�b߀"��p���� ��-q�-k�y*�ya;���秸�ט�PoL��í0A�	��D�A[Y��Q)�6�0�}h�=x�;lac�Z1�͈���7x�7�A�~�pft�Zjr=շ"y.�2�pt�,�&f(�²@e0W�#�ڻ�Gލ��5ls�:A@!Y��)��61T'6�ӵ[ɑ���~�Gg|qf�(��-��Վ3
6�,
�q1Pm��Uµ���p����*���gD��,k���u����@V�4������ЊN&��۲��8���/r(��ɴ�\�IоXٕ"��K�$Ǡ��@�1>�|��A��^�#�.Q1T�)y��F���e�;���GW��+DTM܅!�9���꺭���w�#�
2S=�?*�����)x�%����O�Aa�D'���:~Ww�2��I�o1{��HV�T~�Q���з�m��^b��p�U�7.���u�|�ѱ��nJ�`\��!��$n�|٬�hA��)����0sx�`�.X.N�?�o�������\i�޿&�lg�'�K���x�y ��g��b�,IN�̇����-��I�-��D���6{Z'@,�?�ae̤�+f/aȞ���|L`��ɀi'�c�.}{z�2��.'�Q��A[o���ah��e]l/��?�