��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ����8��x���
~���͵5=��@���62Pb���0�x��!N�����4�K���C�AHC"&X� ����D$��O;�l+��d�w J�۞f���;4�$��l	�lCN��4+��~���TL����٘��Ȱp��nax�撠��_��"���0���I�g� ��>T�p�k*Ժ6�l��P2�h��%��!�/���t�աw����e���M�{X�	F�N��{N\(�h����>��P�Z{jLc�i�,��T([J�R�к�	���IU*e6��@�5V��KWJ,�hX����}��#4�g��&��N^(H���}L�,��G�M��>�g1շ����ƛ콼���!�����"�;3�1�),��ћ�W���:�|�3/|[*�v�s�竀Ak��n�\c]G�XW��X�u�1s
j�������"
��4�չ�ˁ&�YG��0����5��W�y��[���td��@#��_��M���B6������H�h�oL6Ղ��k]�y;%�r��ǣ�1�����v�(��h��W�f&�A���Cd�%q賞	(!U^R��u�Dsҋ(}$���s�;DBH�n���.V��& 7����9���0��w�W��r�;�ҥ�u6	����S��6�@�Oā���s�`aU%�ڭ�������0��"MN4�[�w<`�]&�z�޴ǟ�'�?
�ruT|t�/*��y���o{�Ν,��|LY��@؉��ؒX0��|�Y�5�Fs��<��ǌ�^S����V�e;T�ߘ[���C4���[���2U/|�R
W��n��r����eP��u�9���$�F�K%����E|ߛM0�gT����U�@���#�m�z&l�
� r�5��F��i�MZ������`X��E���c�3����r(���߾L���R�C�|�PM�-Ù��+��ݠI����v�{�������FN@C鿏�?&gk6�ߵ޸��t��"
�te�����'\����ˬA3Y�p���}}ư�~�B%�[\Fq�5��2N��h�;"25��埚����U��x�b��� K	(�-f��1h7�����b$���Lcs%p�g9����Q�5�߻�zoC��ό�&��!�l�%q�F��7�LR��iVw���J�Tr����Gw@�|�F��c�����z�;�����;U1O��
e@R�Љ�d�;=:CC�ao��0�,��F��
��jk6�B!���S�B��؋	8�G8�̊��F��c2y�����vOQ�� Lb<*z�ΉnN��P�Ӹ+E�^>�=*V�3g&'�a5�9�\�x���5�L�P<ǂh����"�iׄm���m�=�qmH3������I�Gc�&?��Q�6W�����y�#@kK�S ���%��רbj�0�u�@�/|p׽z�\R����0�y+�H�ʲ�#�j�Bl�(�YUO���E
1o�6�Z�NLb� �>(=�	a�d��EG��K�ӝ�j�u�)�1�u�}��wDM�O�ޔ<&�����[��cS1�͜�^��o"M��)�2��V��Q�p�p�J%mC`BҥZv�qd�;��i� ����E���j��H�5��[DJvY�&�<��p�00�8��7Y�z�K�V}:e��F�nW58r���GB�!�a���(�uI��>Y!:H��B����5'd��НkdB�Dݵ����Q��h�����V��A��^�oK��p1:v������@��sz�3�<v�g���v@݅�]3w�"�Q��T:�ƺ�!&oOM�5��p.@%�E\Ų��&I5fV�!�v��r�FՇH*����;��'�潫����;7��eq��Vy���mӪ?�:�����	C�ח]�'�؏œl6�@g�s`n�s����@�͉'�9���C��Wt5�H���JR�o�;m-^�Z�x�>�����JQ_xU��n����;8����ר���ټTJ4`UziI>^/�]|�����������-�|d�J|�$S���]sb�n�h���Zā!��V%��5�ޔ�@/
���%8���@R�z߇�����;�S�	�i$��-"	<�P��iL_AZ�ݟ�"!���F�"x��פ��I?�l�)8���"Lm@����&���B'*���sc�P�M\-���\���y�\W�H���{��oI�}�5�+ȦgZ74���1>G�a��3��~��h�/�(�f�) ��u .g���0R�'�E���W�'�����0�˫��R�����qٷgOȾ"1�_�+��L�7AniWZ�q����F�21A&<�������4�h�����X���B@��1��be�4��̝��]	��A�RZ��>�P�a�k�⍄�6�t-�`p��=��ݵCc��?|m8L%��ٯG����Vl��&p��\��ZJ [�6����_4��=ܗ�g9ŤM>�!�������M�j5T-V�e������>~�>mg���Wj:��f�)��q����	����uTkgT�=�6���	�M������G�W�>"4�f6^a����R89#��l&��0%m�Tz�L�X�I޼�,CݷZ�g\$�C_i ��R�C<��:Č(��?��W�`�M�M�P�f��}�%����ۑ%�j'�2��/t:}�ou&_����e�c���C�������2�q���cIc��֢{�<���� ���x��˯4b�l��O�GaR�a��wy��|��I�Z���t�?c="Dt��!)f0{&��/<spE�LZ=%赖��N*n\�5�9�]'�{(ï�%B�W�y�i�����[�)�@�FKڔ�H~e	����܉(��&֖T#����P�]R�?�sV]6����3�'cӰ�b1�(��'� ����#̳��l%&`>T
*\�y?��xj@F_xD]Ɠ���;�.'�dT�4��e M	ڊ���^U��ֲ���r>5ŗ�6*�R3v!�C��E�@E5����kO�#���B?��zs����Ft9�����|.���l^w�}_��P�O��������%<�ڃ4���9�����N���=KWu&F��e�%���s)�,+�{��G�/�GӞ��u���׼_�Hd��D��? �_%�ᡎ��شR����%n��w��v��q��:H��F)�ı�[냴��z�wV��n��EJ��Gy����㸠F��K��:�8�aH�Y|OSٔ4���U�D��]Q���|f�<?݊.����{��l�Q�x��P\$y���Q׼ő��hV��5'S5#K�#U���e�û�L��V�sB�͖o9�
��ٞH����iZ��\�0�;�4?6���`� e��@ U���d��SfN9.��ۨz��	�<jr�@�@�Ob��v� ����uZ/y�`� Af�Pb��OQ��҂9�/�d�-���2e+�OĜq�?��]��� �ۃ�UVL0���$���J�`�����JV
Y�+>/���n���7�hv��Y��PvYƵx%�F�=��>Z^�nV��̈䱻���*�G��;�	o�_�M��Z��JBؚs眰�Z����X�x��2hޱaO���/�1���Óɴ�w+m^��s8���q�G��ua��1�Mw�yi��9o]J#t|��x̜jه�L�eH��#g��dw�1
K�D�1�����y�]3��x��7�	lT��u���۔w�2�,����ƪߵ+���;�j�f۔T.ܱ��1��S��څ�y��*���mw�m���z�C������su��>����T�����U��&T`�5=1iq�d%%fDp�:���ϧ�-�zp�ܙ^k��HH���=�/��ϐ�	ki;���!V8�EvJ��F��k�?|�#SX�:{V@*́�f�L��H��(�M�������H��8���|U/i_�R7�4�g�唫)J��vr���4o���6%�(������틞��������}�#]Utx�"|����� �E��?��Sl�wy��WM/W�����T�Nmv�6V�䠝m�����l��4����.�kw���I��e����J���Oֲ���0�o9����YbQ����/�����r�T$��%���5{�E7���+K��a. IS'�̓�7�QI�FA����n����\i"�]�t�t
����^�ͨ�#Q�Xs���Sz���F�@��/A�k.�%�~q�{�Q��趘����O�k��T�T�.�,&C�%#�AG��j���>�i��W�Q��t�ؔn�&Z�)��� ��{�����Y�S�,�w��v(y웾��#�ΤF!�aG���_��)n{�h9X2,?�^��R�y���坮c��/�h#n�<�+��E>m�d�(
��Z�cX�j�l�<�d0�"9���a�(x�́L>#�V�Q�.�]����Z��91+Ѯތ�e�c+Go�H��]�P�J���;�F�=�s���[E==��`�l7O�|� +� +7��qd���P({��k�1��w.����)(��U+?��羥/�����C��]�k�XP�o�s/��s���,i��KkY�v��$)�l��X��e3��`��H�r�FW�/�P~��\��s��4�8�<a�imةSY�������.�n]���Vox��m^O�l�G؀.��:do�I���*���*^�s�^��n�v������������T�(����Gl�[Y,��%�t/7����V��rZ��׫��|���O��y�H��F�� ���j=��V1��(�˩��Vmo�Z�~C#1,�@rm0�\05Բj��s��2e@���D�	�Tܡ��O��u��뿡Lw�/��5�������W+,��4|�*�,-hT��<5�$�C��ܢ�<���,��?����릏vk�5<��	�r�4�n�|�%ek=��P���抙%y�^P��J�b�U�3�I�|�gX��_~���j��Ba��`�+>F�:)7���M�]��o ǧji{k���{&X/��b�q� �V��3mZX�Ct3�2k5m��o��xH/��[�(�U��=���*�-�aǫa���U�QD��^��j�)A���uw����ʂ	�����q�IS�PkƐI$ۈ�Qt��D��CM	����v�(��e��,/��$lן5�Z^  �@�<��(B�����Z���$g�$����Lj�g��e�&�5����h�)��Q:m�0�+f��%��#�ɓ�<4;-����V�ZS��vS��b�?dr�L�tdN��,���4�e� W:�gԩ2J��d,H�4�eb���TJOyFn�6'�q��'���ғ��A���cg���q�{�YN`5�(�	���b ��U��w^�U��ޱhu��*@^�ǭQ[�	o1����&�U"Q���.K�}~��@*�o�)`��C��%1\{Z��7�<W�������kߖ�u��г8�3Aձ�~O������4�N�����~�����d�~�	���}�5Z`��\�1�Q� ��y�,�I~&��#>E ��K��a	o]���@��m�����}�{b0��1�o�`
�����;�R� Dw�5-t���q�6�=bҌ���[Z�&�Co�F�m[}+��5�R���X-��R�
�P�3mZ���2%Fw2��ISD`	>]ׅ* �$ˀw�9�E4�أ!tϨ��t�J�n�z��n=+i ��U�N0r1�י>	e������b �69R�Ɖ�M��>�w��p�7��d��7�Q%�ԓ���a�߀R��D�����9��vwpn!�����R�O�o���R�bKv�+( Ow�9M3"�>�2��i������Ԗ��F�3�LR�0�
�gYK,��v:�앪
-�>�e�;+�v��2�%w����6�h9*���-�l����!��ʏUh6.�3�4�c�2��zN �
�$b{�@V����W��*r�����۪fQ���bKf ������FQw���9R�1_>�Ѭ���Y���ƣ����r�Ȥ0)�N)q���X[�$�12�^�ؐ�x�V��?d&+i�,��D�}��ُ��<�I�*��Z�j.�@��@F���,�vr�"'�b�6��wP�<�~$iHTs��#�d~Q�����.�
��G��Ws�2lO�V��Lb�6>O���,�z"���1���Q9[��o�܀��]�y��o2���9� ������t�f��~��j$�r	�����9���Г�����h�S� ���!nhNRK��4ВoE��85 _�Oe�r|L�S��� =���Q�=x֙:��M�k������W9�� ^+N(��]�p��Y#v�;��^M��n�~���ռ�<��bng�Z����#�F槝!��
�(��H��Ў/-1�T�̉����y��e8��"����6��D�h��j��b0�*F=�d�F�n�@��L�J��_�x��gl/�y�31+��"C��z1�#����_��y|u�+#��K8��d�B�������I@�LUk�)�x��ǰ�'%�WDnά�יb]��B��4\G����j���A�)��n�]���8"�Q����j+z�$89$��Bb���:G*#����m-�~�����SJ��p����2���$�I!���hQ��j������Y�p�d�H)�˚e�2����ެÆ��m��0g��Y����|�y�W�3�1Z[������ҁ=ɽ�T@UG[��7�"�X�g�'d�@j����Bw��U�'���F�܏^,Z�v�P����Gt:;�Nr���Z�M�u���.}a�!��m�B�08|8qG�;��~���Bd�Q�F��ȉ낞��ك0�Rzy�,	VD3� }�b\E ��[���C�Hݸ�G��h�[�Ƀ��G���c�S���$�3�L�+)�?��r�n��yg�Y�Oj+�,e����8����h����m6a���W�3q
,�"�N	��O׵�˿1�1�H�����E>���P
�T�t8)��(^)Fq�q��Z?�F_ �XP�Q��/���R�rU_LQ*�V�M���iIj8��qΉF���S��q���El�k� 4���b6�>1'i���������hX=��>�.����$�3�Ar�c�5HK��s��>�<m���2k��ʲmg��Y���]��4u��8��߾w������y����?!�Ǽ6+��iMf%� �K� �@B�*�S9��n4yS'�;s}4�x��R�M"	r\d��ʹ7¹�̂���j��D<0լ�i�<8�^W=(�����Pk�*[��]��w�����0�� ��%k�^TNN0�V�3KY><��P��:�|?ʧ���3X#�l�x]F��-E�����ǄX�~��)�����O��-.�}���AV�)&��x����T�2L\C�.3���r:D�I���I�'Nk/VOI4!�f�l�H�:ʭfb�T�~�\I�l�޵[n8�]��A���ym�H�GA}�^u��(�˒���-/i���o.�<��LP|�a3��+��HG����KT�Z��.�]�ĲjX�#���L@B���=�u�=���5r�$�#�H��`!f_��
^;���C ����9:/L�Q��lA�"
0�J,Cܐ�R�U���2~<���U�'*_�E�~�q
�`ך��o��`$�@$*��H4�����om���+�A47)�y��S_��,�=�C�W�T��s��&�^� �Fɝ��6���嚤p��p�X�Q8��&}zo ���G/k�	���,YG.��Q8�bs�f"�C~/Q���T'z	��)�q-&f�)ƍ��;�}=F8tD#V��
�O��~4�O�U��@�s����Bڅ�DW$��Y��\����wb�����h/�������ʇ��9Kȧ���p�č��d��V�;XkN/�Y�,�!G0��Ŕw�TM�����?�z��@��a��D��G;�S�0[R�Z$#ǭ�
4������yt���I�w��$��G2��Uk_��MDŢf&~�Eg�f��k,�x����^#Ro�{�a,���8��9B��c\�GٗFxMJ6{�=f���_�`5"�Lӌ#�Q���C���v�� x�d�AM���o����sh۾��	�:v��,67d�������֞xZ��i:ӣ�i�
j��7��`>�?C��	¶sJ�:��d�	U����**��ѽ�ʮP.ڇ������Eͅd2,�6۫l��{�W�� V�:�I��B5�G0�m��,o���t$�cr��(D��b���,�o� ���9`���I{��1�9�U{�`P���VTU��H,|�M�<��N�֚xn�0eS���
�r&/����n�8�s���~u`s�Ǜ�d��[�&0��v�Y���F�@�-IsJm��n��޼{"4��ʲ0��}J��v���/�t�;���v�����y�
:��HDsr�b~�͊�j B�'?8aU�+}A��[5�C4�!�:p<b����Bo,�ΤeM-�֮���odm�D#M���:��12��(��t�آna~>=��u2�ȍ|6���k���CO��;�M	_OuڽM:`N�;;s�9:�ކ�{�z���8YJ�C���^�;&�<I"�P؜��ۚ(ڛ�q�0ݡHqsM~Q'��C!x) mT���"�jL���t��&*���~Id��]�ȋ�E�%2�p��Q�c��"P�$��]�l�-��%&�)���C�$2g��&J��k��fTU˿x�����{H�m6a�?<@���?���v��ؖ^��8�w�pQ�h\8�����CS�.�A�D�o�QZ�)�˝�m�h�f��Wh��<D)@�)�yA,Ϫq��<���}�E.5�繰���v��p��bW�,�H{����"{��:d�Ҽ�>���PH)��pmP�
V`��hڑ�?0y�