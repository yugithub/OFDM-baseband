��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ'���ugJ�J��G�m�����	������)����q����G^?jt���ja(�Υ��Y(0�̐<�.� _U!&�-�.�5�!7����>��(��C�:1尃���J�.x��'�c&��\Ġ�}�~E[dC�~L&0�l�n�gǜ��z�v�{�x����e���F��a�PІ�TeMņJf������n;��wL��#�ccK�?'d�M"
��V��W�.���8!��6��H��gC�O��K+@��'-V���5�fq�h��l��{��'7����31L����ɥw�P/V9��,��.RN�>RS�T Ω��dd���.��U�|���I@�ơ}�����V�?NЩ_~�%��:{�V���Y���2�Q<`8B_S�Y@u&y�u�H9V��:k8$���V�=�-%7�Q[1�q!���|lG�3�~ǭ�8���k�r���~P0��e�C&��F�G�%��LW�4�0t{s�����~�`����SC={���ElJ�I�Ԙ��nR/�]5�Q�V_�>d��pN"��)��\��@�\��}~Ɓ9������O�pz5���S
29����2�7�#ή�vf9�*G��y����	m? ��%�4�������Pċ]W���w\�Zÿ��AΣ=� ��Rɛө��ij�	?��6tN~���\�����xd�#T��?�wM�x����VXs )TL,�e�U��}*`���a��	���	���z�QF3D+�D웢�@�f�5�!J!�]��H�)*&���A^Xs6㯂T!��Ut����S/vxI�}�4u��X���h�ýsw��Z˶sV}��*������:(��Q
mw����'���Փ\�0=9 3A�qd^p]������mfI�y�_�w̪��?�O��CEr� ���d{�,t�)���t�G_����E���ܘ�2T��ř=i���Eҷl���ZB
=s
S�I��FP{D��<�C�O���
o�����f�4&g���?��iS�I.9j
?D�0�Dŉ7��p�7;�7��ڛ�pm7���7�]�Uz�!��z�3��Ch1���zɶ0�����>��h:�6�Yw�"XY�{"#��_�]�����0y�N*ZȅU��z���p0�LUNZ��~����Y9Ga"vh��Q�(�#���1�BJ���C4�6�m�P�?t����~�?���2���2�x�f