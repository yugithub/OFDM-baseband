��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ��O'-�d%#��Pi\��0C�x���*��IR�~ry����x�wJ����,�$ ����f0l��L�kb���<�rPĥ���f�U�j����6�$��dF!���^Z�ҭ;t�p�B��Imj�r���.����7�/�"ǩ�9S�5j�YckQ�G��?
`7�xjs@d�PRV�$V�c�s?�1I��U="��5H*8����2I�|��l�&�S�O�v�<�6:%9+HN���I%�m�,s������'�Ⓥ{�ơ���0��u����_`,����46� �*���ߦ�e������
"����,��-?��#�H��d���HM���CV�Px����b� ��՛��[{�/��my�u��|�U����a��~nؽ�GH6��n_1Ϳ̶��6~;b��~ֺl�=qxd�D���K�T�6�6dO��EI�������:OY�8D}1��-Xr�#1;���d���~{����`�4l��Z��0�mQ�@����N\g*0=�:�\�%�͂��e����]�sT ��A�(��4\�ۨY�=W��dD�&4�Eɻa)�ckO���M0��\Rn1P:�iv�kq��ۖ�V���a��S)����ў����մ~��fsI�x����B��L�/сgB0=E��Fi/��z�B-V���� ��S�Ͳ$�hQ��������.O��C��H(�8�/\m�c�`���x�;*LN����������4��I�����a����������x0k�Hk,�䎌;�K���-��[���}�~�Z9NFz����5ś����i��T?�'�"����Z�ݏ�]�3��\xwiZѥ��:D��}��+���w��W6�<̮�����m��|i0:��:ߗ^)r�lN7ۏs���:9�l�Nj����<���V���� �)�պ�f���pG�65nv� E
6],\9��G��ȃ6���+HA�2M�#��]VT#�WJ��i���Mc�w@DQ�i�o�z4~��;����Hm�/�J���SR��τ����I:����D��x�qK�å��:�_����[߼&��>]����������5z�D�3�I�� ��#z3'�y�rθuKD��?fV/P
ʛ1fɌ{zݶ1^e�kZB�wo۰L��p�^;ּ�����T�zH�����G<<��c�	�o�-�2�����о|�O��;�'Ls�&n.7k2�ˈ�GM�V�2]���.Iv'��P,��u��L7�$�r�W�w6{�#r�,�0�`�ed�.��an֙����`��Jg��ݒ*(C��1hg�ֹ�m�tRЗ܉<[C��,:�R��9�3Β�T��h��������y�xVc1�,��1���L����ӱ��|��5U��mHۺ���1�m_�%�}�%�D�D1�Lf�()�S9AQ�.�&��OQ��a�/��?�8���tUЪ|k�9��R��n'\�R@{�W�0�T�9�`AU\���q�6�o�Q��^.Ԥ$�ₒ*1��dUw�^��G8cŞ!ʊ�S���w�*<�e��� Hņ�MWly�"jk��V̔/٧Ίm(bc�p^��1sB�� ��txb��4��_泖C�T�> �	�]�aM,�z�٧"��I5�9G�����NKu��4��Pg��z��*
|*Ѐe��heS�SL�H,u��,�YO�=y��h�mH|��������K��c��ky��e�^��eп�Q�Zr-so����&,`9��U-�hϐ�j���TfRly�L����4�Lo���A���ch�"NK>��, Lǵ��K1'!6+Co�b���r�����\��FNys\+m��x��Hz`�ΰѠV���5�jt"��ك�#��Qj���ś����/�x��:X� ��Qi	S�P�c���Vt&`G�bxs*ꋈ���F
�U#e��_R�����)q��(�,f8�S`�t�N$�I6xA�+���?��5��C�
�o6xcyN�w{�j*"|G���OT�$�W����vMd�e7�g2��]T]�A|v56Ց9 ��
��ǂ��1����$�1�Mdw����R�}�����<�s_��%Jm�V���J�Z��Ÿ���)	[���B�Q���e*�}ݎQ��ڟ!Flj�급���`a�E�h�h{�L}��z~@��[��b�3�,g�IԲl�'�li��G|����#���D�1?Ց��E��si������̶��~���sJ�k|��r��Qn})��^2�)0_�I�F[6Mg4�+�Ё����G����M����_�וO>��W63ٹ��x��L�~x���W`Ɓu�t��|�t�)�*`�T��,K�±�Q_\��Mu���	r�����ݑ"�it��*�K�%��]v�eB�����|���Ĳ\�Զ�P��@��a6@��[����E�U������p=ݟ��Iw�qJ���8nO��w't3-�c���k)ƿ>�A(���E��w�C׼�O>�51�Wp(2�G@�i�sàea�T������iCk^����R�/�8i&ܪZe�t�ƱKzl��V���@����/`�Nk�}����A�c�/5��F`��y���o�Xk���rV��k��-�5l[�9KlC��������%�C�%3��,����Ӊ� �����`�0�M� ��f�����B��T��D��L(����/��<�׈m����]k���.�� \Ĭ����nױ���R�u²p4��Z"�� ��:]�(-L ���&;�����R+oɶ� Fj9��X˚3P��Z�C�Ң�UR�=�'�jz�H)��[H�ߠ��&{��ӫ���Σ�����4b\l��Q�4	�0;�r�6�.Y*��6��������Ex���<~zU����D��j*vkn���m�%��]�{1�h�:ꬋ$�+�O>V�}��"W�(�4}kdd1M����D�q�����F��2�{��� �z񾖩�U�Q��R���q
_*�p^Y%��S-0h��W͌pe ��U�ڿ�i��q�8&r/�X~M�I�O����iȂS�"��*P-\_����ߑv�n�?����t���D�w�pt�P�>�I��]��w���s�1k4�_ʔ4���8�1���ן�OOq|�]�bV\�s�?�L��=���b'@1�4�S}����CMP1��3���^h��W�ޓ�3w��#	o�W�C�6�L����)s*ʆ
UL��^��?Y�"�XGώ�r��Eݑ=p]�	V�H$w�p�%g����C!H�����8'v._,�$�KA��R��c����?ha��m�1:I@�q�[ڠ�|q�ڛ�f��d��4�:�("y���)K��k���Ь�G�gB�6n�Y���Ԛ�����z����Ox��bkjʞ&�]��C�)�R�N&�!���*V�8�e}Ny["ϒQf94ǽD�WtZW�[�9��C�����
��e�73E�Ɨ�BՕ��hӺ���fU��m!��Q?`�n�x�|E}H�Ox �k!�V��_�`(�򌂴�J��N�����t�Dm����N���$^
�g�R�_����H�����!e��s�Pț>N�)>ѴE[T����W�[�ג�Zc���3�����tN�8܋K�Ɖ�E�s������P/D�f���1e>�/LS��|Kf[.�d
0@.���(�m"
���~n�
}��L˞vk���N�W�n�kڮ��YL#���C����I�9:��
4�}��+�d�i�L��<F��cs�S+s��z�oQ� �df^'�D.�FΨu��8++j�I6�]nW�L�Z��q�R����a����n>ä~�$SGm��_j��u�`��
�/C�'�� QC�n�&=�z���o��,�M��J��J0�{���.�V�P���!v?NK�y��-��9�#���R'��9n1s��`N p(����,>f���9V�]2�;X�3��"]x+R	�WBː�qd�b�j����^w"�f���'���Q9H�x8ߢa�it3L�M������x�{���vM���Z�|~=|H
˜6h��Yz�'<
3e����5��Y�G~wˌ��5+�.mAX�,BrP���M��7�$7�X��'�ی���t��s�����u��5���Y��,���M�J�.�C �q���9����h�"���P6ۦ.�M/��W��F=���s���nQ�v�qH�v,�o�ͭ���l;PgoQT\A�S����;�w� Ie s����KR�c(��/��{e&��� �丁5e�m-�� t'E]���H�]�EV͟h]��Vxk4!QD��j��]zc�'���B��^в��nG�gц�����J�O��ǰ{)��/�%�#�~7�K��g�
��p���t�n���>?;�, 
.�w;�Y�"�uZś#��:?1M��!Ak���8�&tZ��?�fז#����K1�UK����ԓ��F�*�M^�D�5	՗��n��0��I��|��l5F�Jm\�Ք�g^¶Qq��y���j�	����Tl
�2�v�D�X���ݪ���ȷS�1?&=�����/.��O�u�x��ƨߋ����5�����/�D��֩ �� p��Y6}rU���0�DkP��=K�����SB�]�n�˼�g�|�)��	;#�ȃ���@T�-�t���]e���Z�.O��3�����m���`��r������Ԑ��!�����I��VG��i�Dy�=�߅��d% ,t�a�El`��-���r���s���Rfڇf�cJ��G��ݞ��NSM�A�JY�|���5�bb[I| @�@0c��d�%R��w�c D1B�V��u��y�d�����!e���T��
��ܴ�E��&ڦ��k��a$.����Q��I�M�c��'�w��B�Z�$j�i��`Z������!.K���SE�ܡr֡3k�㆕:�d��璣��:3.�t,���,m�������~������.~�\�6�E��\!0b
�����9���z|�+7��N��D}������%�/� [F�;U+ޥݮ�^����		��8 di��ҍ��#.ΰ�����ԣ.F�p��q{F���i�fK�\���cW��������5���U���O57�;$%M���J�&�Ki��XU��,C�j����ȿ�-���l�0]����1��紈@���a	7�xh_����Q��!�]N�/��>�k`uys��������*|`] ?+�D��M�A��4�� �lp�L$ڒ�bi�p� �VȦLԞh�v���	ī�"^����g�=q��h�;d��uy�T�\�z��h&b��G��.�n�h��yv�nlE��� ���}�Zk���;SN3k���C�On�C�I�pq�"�<��wT����~�h��6��R�2���[�H那�n�y�]�N��,*1E`��&�](|��0�&�*cA���鸄ôDP�"^(,{вۢ�j���n��szه��br�붋�=0cC���Dk��T�M�?����h��a��y;�ζ�9/Iv�9�M����1�N�Y�̺��W��1�^�3C�*�y%a���!;ϿkϠ��b�Zu����c*��䜪>��	��Ks|:��[/�S���`��7d5�v�[��Y%v���Z�Qf��7q��:+Ӛ���E�<���T,X>mfA�pZ��i�&3��O�ը���ߎ��T�R���$4��y[t4m����1��q��"�� �ޒ����P�\o���P�X���f,#��/տBR�j	]��#k��Z�L���Ma	F�w�=��]C=z�TW����o4�N��F��ˀ�d�@�ևDio��}��/�.��GV��)8N����S�B�ᢕi�8����_�ԴOx֩��i���>��;˗y�t�xB��� �7�ȓ�?�$�J��Gg,Ha�#ȏ���"�z���ݘዘ�@�y8~��q�V&v��'�idD�\�%I�ɰ�f�ׯDY���-�;l���?��W�1��?]%�+�rR��Uk�-�q�J���i�� ��Rأ6�VF�C`��X�*I�I4��f�`�ٔi��VX�lW���{�ļ�����1Y�7
t�YB��+u�h���q����t�]��S���{������'�~��T"U��S3-�����Ġ���.�@��$�	�5�PgȆ�a[X治t�m�qr�t��&��/�u�Z06\H1K8@�TϠ�#�I���F-������YgE�ϔ����A�<7,�K~��#1�N�����)�nU?�~��As�|��%���]��l���d���2����!>��Pc�t�bۯ�fj��i�d`�+5�<"X�9�+c ����� Q,��)��>QoұĨ�/�+W��@С�g��~y���G/鰑��:��f���O	bD�Q���AO�7�������]S�rV���
����I�
�%/ZHC��u��Sޘ����D��+�3�ROÙHnZ��`����%�K����)|>��?.�l�k��(�]KM�`�D��j5%ڷ{��@a��xx�c�Ĝ�I�@��S\�}#�#��w���M�ꡩ%�����`IfXx��w���4H�����!%{\͚�|�[H�d�c�[u��K��^B�^��P�2@�E��f�Z���%I��<�z)�r&���ض�{�B��x)oNw��a�����������L�6N@�����	8�φ�hKV����h�
99�+ԉމJ�#@DW�@3U%ȯ#)��<�����y�L��
KLV��WW�P����t_�O׃����2��T�)�@я�p��q��1��`G{ؔ �c�����X}�緓/2Lݑ'�e?�����C(EB[����sp.*A�C"^Z߹�ᬓ��$�}���3���L��h�
�]�,�h��2W��!�#BfS0��]�p�B�$�9�>�m�
�!T� �kL���W�3�� ����|�[�������3�8j���n9�p�l,l��A�/-���j}%�\��Ѯm��m�9�hv�˪�#|x�6"
�<|'���'o�|�woTt�	P@�P0D�Ӆ�S�7�&��)�G�m@�?R�q��l�;)oX���T�E�}'���-���ݍ�=?-�g�Z7��fz�;0P����f��@ф��K�������W���%� 8���S�|O�`fh�C�=	-N�^�+����-�B �b�VO� �7k�>\(�x�g��!���X�s��+w�L~\�Z/S~ʹ�0���hS�b6:���?~�r����&�_���p��P��d�&�����T���뢕 �-�̭>
�k�<��P����&B��1����X�4�"ns�}��Iq-�	rfI��Ύ�c�)��._����b��)�#�2#0�'�p���΋5�N��b[�@f�8�^=������W}+�2��Ź|%0*�G�ɪ�z��~���XgҎ��|�=��t��?����es��,ܷRo���h����XHY�(��E�
G��t����r�]VZ_	�t�\~Fs��j�ޕ�fȎ���%x'��%WS O>@�,�5~��®������51��(`<,`̤3�=9�G/�`.v�z�c�{M*2�F\ڑ�T�i�^"�
�0�����d۵ֹN��#+��.�`DP����q�@4sL��PK�œ�]H���.4[��Ü2^�E� ����s0S�I�ܬΜ{[ݠ(bc��e���ą�>�XA�
*%��-�����T������(�M���a����g�j#�������e�S��H�9�9�R��$x�
��f�����S�W��@Po�ܢ���~\�PZ��@&���:������C�m?	�P�������>9с��D�6�� s�(�s�W+=�u�t���7	*���2���|������R����Ő��yj�7f�J9	늊�a��&�Qm��rlQ������K*�QJC?�'#���	�S�ĉ��M��$�S&d?�7���Ji��\�� �'d߹�ᬓV���~�AȀ$0��:5�V��՚;A���4]��U�V�+{�����Cj-d��J�b���#p��)ŽsϹ	.#�X�Jb�iK�)$�������ĥ
���2SZ۪�z}���
T޶�ʌ�����YO�l��*�bG!"����^�c�(y��d\3�T��υ�l��M�Z�Fw���E6��_�6C��X��K��w�Gݾ����Z��<�ȁt���YhI���q���	�ѯG;X�������0��ݩ�l9ѷd[�f��2_3]�q5Wg�)��$e2��$UR,�ՕG���j?�!�*����O��F�D"��";�>e�d7�[��K?9
wV�a�	P@L�z�cx�C̒�q�ҒO�E p#�{��1���dn��h!-N�
H�=(�/xӬ
<��K�]#��92�q�Kj�O h�+Jۄ-$_�f#W���Oom�-d�(|?|c�����d��Jk&^�P<��n�=�1:aۛ8]��TPZ៻]��U��E�>��?�	5*8�v�q������������z}1rb�w���l� ����Z��G������?`�1��U��/�Y�'-c��L���8[�b0��V���i/�3J���r�Ǝ�l>�N����ӟ��x�H@�;�*���]�J��/�CpͅvM�?�e��&7:s��yD�"P`����5�:�|��_��f�?�ն�����< �V.*-��$\�!8)'���k�=���� m{C�4P�Q�������N�A�\�ǩ�/P���,��i�1�=$���e�����l��իq��2�X#sB&K�%���<�[�
_��ov�U�&�����Zͥ���pd/=D7��9�`�Q�E2P��G��SM+�Iy��9ZΣ���Κ���� ���>ʦߘv��h��B�~�ȍ���l)�o�����ڻ�64�i�i1&�nQ�<�Ө>�#(�`�Ҧ9� u�q�$'���цSf�=ӎ�|��$�����|�㌷�@��'��d�_����b�&�8�/E�i	�~+��8_��z�S�O������T�N�Zl'Q3 l��$�Y�^�{�_2*�Lb��� ^�߱f���?�EPM����]�hnb?�1����t�����@�g�1�����Ry�$N��<����#t����4�I�����L[���v^��0�A���K(�2�����;�>�����d���+^���	`WRU�v(_(�$ ��e�D:����)�գ�eV1�A�u	�+)�ik��[~����ݼn��r���|/a&п��6P��I�r��H-1�=~|���5y^�/6@�-:c^�T��-�X�Ꜫ�n���;���|j�ћ�+*F���p[h=1m8"*��U7������� �����yN��Я��U�g�LI��I��N�D����,��`�V�]�^��4�␚ǲ�����@�,AXs5w= b���l��<�+��%^T�{�YO|Eju�{��p�����wIR<�	W�Ai��"FN�D�x��S�����b�y��I�Yū�7�+�Iz�(8��,Vcۭe��F.���ΥaV
�4>~[Fn�����j�m,�[��\<��S�2�0ɹ�V�%��Q2�Q����]R����6��� ~�0��Q�j�$~���o���]�f+�ስ��u���a�/�aaK0�6�M?(W��$�ha[&�8�������{G�:+����q70o���.-���yz+}~��|����U<�r�P0��䄹�w'5Җ
�]%�(qGr���+�.X_��<N���=�c꓋%�9(ɺ�'�����gz�ց o��?|�����nQǬ+� (L�����������u�Ż[�2m�c>�1r�n#��B_%9"�2~�9%�EI��'AN��4�0bS�'D���KSNǥ�@�(��?��}n��XW�y�+K^.O�ɛk�ӆB�{������x�:�� �~�:`S�SB�e?��s|�������T�Jl"�Vg���JS�Y8W�H�ajP(�ɠ�2�d�Mx��
#�XB�jl�	0Ir���L�3�e"��vJ�O�Ȃ_w]B��l4�;���u��=-�����S֫dt�n��E8�Ro���믦=����Ղ@�r�/6�B��۟��xs��|���ґ˃��O����{,�7�Ս'�Z�g"h8Uf=��'���Jj�b�����8������f�GG]Q����p'q��B�ӜEW���s��8[^��n{]�1�%���9\Qb���Z��"��r��/��üܢ%�~Q���'�"�jy3�4Қl�`�"�Pq�N���C�m��AԊi�g�����k�7��X�,�X��Wf'$n|�y@�Is;�d�4� H��� 2�a	�S����ࠉH�U,~�������K$���sU�"d �P�3�Į�����gW±���!kW1�f��k���ș�W~�ھ�ϖW�=B�Lӷ	�.x�����&�8�� �HI49Rye߉ �TIpiF�7j�{�Z�Ρa��IV�i=3$�庰��|��>���ë��K?0�	��� ���$�j�҈���%MsMU�Р�CV�{���$�n�l2a�#H�%����lu|ù�*?{���J�}?kzIj��mt>d��#�p���\�9!��7�/ք�fb� �G7^������zv��]�?�|�t%T��~W�H���
ā���Le7Du�s��)��G�Y��1x���D���3�Ø]tN%�u�JhyuN��V��ݵ���@�_kX4�q�x�_:S����Y���&�����Q��SR�/��NYMnsHU��MA�s�r->K/��~����Z��Lp5�%�ƅZ�5v��7�;p����m`-.!�	Y�&�p��7^U7�L��Y|̂�u�K��Q�CabI�MƉ������]�3�&�+��Ec����D��UϑR3T��$���w/HQl��d���e8���D޳�e�D;ثg��#�fV������P�Ԓ�v���'NN�?yy;�!\�H}[��u;���47v~Q>؅׽S��Z�^�*P\��9M�~BD�ȽJ��7�~�Cɔ?I�H)�V��{N��Qz�PR��P��.`�~����t���/=�0��]&�*Q���A�%��5+�[�W*�m:�=o��H._6^1�xn�-z��=$�N��X�[��%�.ָ��?G�ٟ�vl�>ɜ=�},�
ug�sc����2��4�^ˬ�ۡS����M���]��3��M�@��� �q||���gh��ۮ�V��I�|��x�c%ZJ�*gũ�E�[�H��%-�
F'��0:F��I���?_oc���b�+��̪'Zx}4��/��I̩��� >y�Kk+^��֨�ȡ҉3ѕ����,���4�}��������Y����f��C�;���NL�"���R�B;�GIl��sr�]D��½��aef��zfE�U�������[�"&U]U�.���Y�v���*��{E���",�*62&�9���K3@���r����4���ӫ�Gۢi���"8��U��j]ݲQ��s�{;:P=�6�m��}[
�hI�vFP�m��L��9��+D�� t��R��7(s�iup;vOv���6��n�_�Gz-�2-�[%��G�!��8jZ	�xO�C<��Hu{¸:�7�2Hkܯ�(<P�P��z0�v+�?��d�'�uG"~,&���&��,/�O��|��n��}���䍱���}�ݛ�u��Gˊ�?�y�'�E$ڻl끵����(n���{�Ï͗�f_-Oz�+q(}��Ɋ_N�}�mؕ߭�(�=*���Wl�"����.|�pg�u)�l�9�V/h+�'����̋�c[ްV��9��9�4�x�v=�"]/�,�f�zՏ�D�H�	��{L�i��#UR���|���ΥA�R?ޞ�J�wJ���}Ic�{��,��1}6nv��T�GЁ��@P�fsV7F���!�7������O��ú�����ȍ�,N�dru�>��ϑD��5%8�V����<4(��]h�v���W�e3NRa4��S��pM�1] F&2���eI���$5ٹ��@�u��u8.�>-��,W�g��tEf��0�����~��L�wZ<v�Pz?���?��Ht`D�:9�Bյ�܋Ƌ�]��ĻNIl�Fӧ�¯���%t�����ߤ�eވ�L��������S��<+�`@Wa����[��	���#)��d(�d�3y����D|��c�k�&P9M��@����0�D�Nrڛ�^��)}Kʧ�D�j�li�d���
-��n�-���=<0�]�ye��L�������yp�kviN��/=�5�|��:�{[�k�*e*�\5vy�nq���D���O�ˋ.��'5���q��ݏ~$�����s��bj�c#��!�ir٫<�<]O0q�Q0����Wq����$��n<�B�BAo������?�̚�x1���&���g�O�Y���گzJP�va��W7,~� x�t�����q�|R�8�%���Jj����3���V!��=l]�{����>	�6�E)'F�rp?�zI�m����>�n�0=��rJ�����Ă�¤N
C��8������m�}�8)�֚6j��fj��# ��@ �\7�H#��%~
L�eo:�|{���Ƒ�ษs�6jΎ����6cy��3��bh��@=G�A��`&3	�����(?�Ȧ�E�w�������#y�}�4[I�ƫ4Y�j�G�d>nP��$iY���]�N�jr�C*��~O��� ϻ��ߡ<G���0�핎�9�[�'��֩�_����*X�*�|oc��d�Z��P�)��g�J��
V���rt����-q[�~ńĿl�������@0���������t�TV�cݪ�7�r[��)=�h԰�h�і�Ky��<w-��������]}+����q]Ȥ|�d:�q��IH�diH�ǁ�#=Ň�s>�QAs��fb-��rPXm�q���n\���g}�'0t��tG�d6��t��� ��i�>�բ�O��v_h���zH��c�DB�~�T�cw���2I3F�ڏ�P����� � �v�ѾdO�9��A��A�E�O[.�{K�%���`Т�0e�G���N�N��;�ᵬ@7_ER�4BmM�
����k��rۃ��sZ�k��]�8��l	�$b��n�}��;PXm�5ؠ�ߤh���,�,3�jI]�`RV���B%5.]l��s5�2r�C*h~8���������c�ӕ<�+�"�>B�Hk��sR�Z3��U�}�=y���E��|�:H��YO����;<�&�������e��bk� ��|P1��G��,m9�/�����UnL��[��A��?���'�|�u�>v&&��k�'�ѧ@�bO�ş�g�g1�o(#9B�7%¬�N�̎���x���
�d���0>����ݬ2p�_n�%����I��;1�����Ӿ`
�����|M����w�ga��0i��"ф����B|a��;��C�va��עv�>M~��t7��z	���{�0{��PV��s#������E��H+
���s�W:6N>�c�f�9st���IP�,s:7�Yv]��Y~��m�;��u�&���p��M��O��9{{P)N�+VR[�M �}Q-V�)��5��ap��~�Z2sZ�z#�W`�2"`��K�)Нe��_ǅ����9D�u�/ȥm�Tvc���%*֊�'�/ .�~�X<�e���h���#▟u��ku�)��n��(���}��ҏ���V#L��¿�2ʼz� }�6m��
�4�;���x�����򠓸�D1��G��i���o��v���q�5"U��m�s�=�K��������^�Z���_$�P����Ǣ����M@�!,�D�:lz�N�!�w�a+mM�a���"�"��3S���z�a$�qh��/�Р�B�33f?�g5��ȷ
=gJ%<$��w��)!�dw�TkT�ں_�%���'����.W0�tH+��P~���L= �5O�lP3Dr1���s��v�s��T��6��I��~v�,�[��"EmS�2v�h]THb5=�"�_!\�r��y?�� FT�D`<6&�+iq*��*7�����[���o!��ȾW�7}Q���� �`�:�0�"���;UG��E)͆�}�8M�^���K���'�{�S����9R�}Jz`K�CB�n��Q��L��c�k/I�]��ő�S���@�\�z���t����CTѸ�11#��J�}��'-��X�A��n�˼�+	�V�t����� ��"m5���%���JgWC���2�A���kZ���.�킺�hb��-¿p�P �<��_p��v8{1/m�'�"�?ᒯ�1B�΂G 4�2U��m�����;p`����Wf>�p�=�+�_82�_�vV�8��(՚Y�]
�V2�;�H��gZ(q�5�K���:���p^_H��X3���E+K�u����&�#�ft
��j��2���b{`4����Q�W5$B��wb4 	<�����4q�%���$E��W��t�&���� s��.I7r��;�K���U]z�T!5������<YD��=����&�R���ݰ�_�ף��ͦ�H����|#��O�9Y�n$�A��ru6pn�>|����'�z,���/|=��q��p�0OBB~�q=mWּW84���_��IZ�o���| �*��<k�ϮQ����r�~/�n����W��_���|¼�{����!����U��87��T�Q��~=Z�oS�f<T��Q�u��Kg�u����_���3�fEEI�Dt5�#"Yc���|�����e�u5��'&�l0��/�xW�ύ�vn��CqC>�M�z$E�1����пH[-	`�E�/4�=L{5�h=d�����(,����˔��)�zl���O��K�)2���\BÖ�%V�������!�>�T
9Y����)�e0A*i�����L�u��� ʡ�����/��e�c��j����F�(\�&���tš��w�O�.�n��o>�A��4�>K@]��%<��i�Bl������Y��v�$��|���p7�̃	,J\�^�yp�gf�/�0܈у+ �f�D	�:�5N�+J����Ÿ!��ّ����j5 ������>-)�	%�>2>�F����IǍ�b
+�揮 k�wެFcG�W�����Y�>)�F��� �K]�]�3^�i�Γ��6+U�>ޏB@Ạl%њ;X��RH�4��j�ٰr���p%"|^2C�Gs`msT�u��~�ۉQ�;��+�X�s=�1���g���Z�׎�/g���S��Y#����m���;�b�!��c.�NW�)"+V��ÇSMɑ �~C�:A��FL>�}�;m>v
�N -����v'-�o��ƭI���@m��J�RK*�c���۴�CX��z����w�Cߧ�v-U�W��Y�Z�_g��xq�7wla��,��� �Jg����Ȧ��t\Ȓ�0��K��a��5y;&3���a�^�4�U���]Z���L�x�c�i�3'$�5�r��BbRϋ�Gt3����2��^��~Mk���4���#-T��Rj<�bA���t��������V*�n&a"{P���Zv��O�AcuTg���"	F���K�F��\$���[N��oy�s�zp�ī�,����ַq������Ȣ���
p��=.�	��q�*ß�������2Q�E1h��l��������N��"��.�}|�/ͫ�RD���q�Qp�Y�Pp@�}t��X
�4^��nH����2��H#�3����'�_)���V�ِ��<��;�������6�^�]<F��ᖨ3׫���OO;����Oa
 �{���@��z���(~˄k��>J�@Ѱ��uGH�w���]@KὯ����&F�%4�AcH�,NI�p��R��aS�VXI�A17�r�y�Z߹ʐ[GP�&[����V�ϙ�,O��
=�$�$�n[G�==�����ט�1�����������K���U���R8Z̅a���"G�~=q����I�B�c8��ejE�vHO(�2@��$�y4��{M)~gn�`Sb�z�:�ºfx4.�2l/���b���.�b\���.S뤓i�D�MXn����̦�*��Zb�&�i ���;�$VZͻ]��Q����C�y��
���ʐ0%�;ۑU.Dx����aE�Q����d��:^a��=��s�y��{��EM��V����\�UyvU��8��"�3"�:ܾ Q�򃥳�)��"ìRG0��M+p[<��8��Q��#�BC0�y����V�vI�^�l3{B��&]ϙ�����xʜ�xO����������ȍw �x��h�Vh��,���Q��;��J" ��!+�]���jm��jΏ��Ȉ�*Ws�����5��Rd�n/�-m�&/��{�
y.�&/�UTq�5
y(d]�-��<��K\��r��y>�j�����a��������n�㈲������)\M�`Y N~���9KRQǤ
\��գ��z����F����iJЦ�!�o����{5�R�d���*f�d�"�����h@^O����PS��a�������
��	�x�q��A�T~�fj��z�/��x�:d�tI��/�1�[6gآ!��}q�%ǽh��*�����[��P<�w�� �%FeP���-N��ٶx-��Z�!��TK��o;1���U�f9������b �q��J��߷	��$�,5Ĺ���*�J�/�?�Z����(R��6lW�1ǚ�6���$��1h�Ka\U)���lV��>�y�Ԍ��� z��v������`��� 5�}�!X��!:I�p&��������*�{Se�p�G�:0��l���/@<5* K��y����n�?���_���i�� �����U;-����\�`V�ɏ��ɭ�Jɨ:#���Ρ�\�	�@6� #�-�Ñr�/Gx�8�坜[�C���B(C֔^,�^��Űh�7�B1�Rg<1H�!^�\�0ŗD��h��=�����3�׾����4JD৳�A��f-h�D�W�9����4l��t�V,��0iS��Lrn(�Qy�nx�F�>�A�ةl�*��
E�L�NK���䮂�5M	<_�6e˔�ʳ�}хPg��mT1YSX��)���%FC�#��ў�l4���/���h_N8�qNy��m�."�<p���F�W�lg	I�k��}�`r��4�Q�SCfZ���nI2�˃�m��93�;`��;�� �]%��|"v^�ޝs�^p�8?��yb�M���v_�#-��E�jU&z��"An.q."#L�����3�L�e3q�VX����)1����fc���l�O]�5��#F��}�7�|�C������
���Ĵ��]
����{qV�Q�|"�����Y��[`+tgD�%2e_���[oG:��:`��*�6�:k���>�X�!�n�8t���������	�*F�%�,_F�PM�=��"^�.�Y��G�?� �B�`�81U���e��ߍ#��9+�2����W���8�o�$Ц�� Kn����R�N��ѓ��fѣ������@��L
Z��:;7<\��ecZ���-4���"g&�� ���IGg�"o�Jde�"����[Z3��Wm6�<�@Kx��̋��e�mv*jS/�g�M�����On��	�.�*,�����C�>���P~��z��<ߠ��k�Q5��E=m0�������gO��N�^�����J�t�|!>h�����'8"�Q�wAѬ2�#���g� ��Mz�&zG֝w)�D�>hR�
�O�t�HF_�/+X��Gin譥�1����(z�:�C�58P�b�7�;ĳB�%��+�����jn'd�%#�M�F(5�_������}�����87�b�U�{�n���Ǌ�Q�ւ!����*���6�$M�U�"Uܬ֫�8�㆛�(�m�c�3����Dm�����@���>��qB'�V�s�DL^ky���)8K����Xw��T�o��ZG��nroQ:��@=B x�
���y�>���(F�IZ�gVǂ*�2boa�����a.����wf��X�Zl�(k�P���� %��%4�$ԧ�*��B��ڠ�1ڔ P�\�YBo2��j����ٕ��""�dK�م����:J֥������&�҇�;��s���tᠻ.,����d�QF4��a�f��Ĝ�}X����ceQ��P=A��3$Y����	�����E�S�-��~�&��QJ��~��
L��e��a0�D���Z-�]"��N{P`tg���(N>r��+�|*�e�&����m���,
G�>�^��b���ʌ����y�v�qW٠��V}�yu���?'҂����ʭW>�, �W}h��V��{��^A{�@�[�2pϕ'VBf	GuJ'��c�"0����$�&�~���2���s�����wxE��/�':��(������S�~�ڧ#��L�����Z)~*��)���CX���mj9+J�Ru,�@,{��y��n�h�\ۀ�-,���͢;FC�7�9{��~� M���3p!��id�Ŵ���a�ȟh�`p�Bx��o�j�|{8q��ߧ=��z��\��1ORQ�F�tEI:��
>u��y>Nw�)��Y����x�~W�L���K ��gx��Q�\��@ȋ�h�m�A�>�K[�6����&�`V�Yۏ;����z�M~|S��8�_��N�@���N�v�/���wy+���V�֠k���JD.��X���ea+�N���H�ЮjefH1j	F�9����!����G���rj�e���{ž3�*9r
�i���o"���lcd��?O�hñ�<f\Z�+��\�y�ȩ�M���]=�pƶ�����C�w�`>�,+)*��#�[5�W�{
�h�kt?'�IM��j�h����_���aC���8��e��k���;�)��X��k1̸�P�br�:�fs��^"�+���m�!�Ӏ���g0y%�Rء����)�#r��j���{e�Ʊ�2����/����j��͆4����cvN[.��z�ۈml�7�,-nT�N�ndd&Ҩ��Z$��Q���%�1���&��RZ#qA��Kn�X7��Aup�g���f�d��L���^��1�K�v���]�+��=����W$�-:�����%e�+��&=9��l�ƞ���tz����zY-�(7��H�w���T]�8*�����h�apT��`����J�T�~�.�ڷ<���?���{V�<��!�p�/�+u�R���}�w �c�<�{�鄺�2O2Xm�u�4����hw���r+Z�ț�#��=��`(�$g�5bmb�6�&%[����0L�tWۻkVi5�6�n��x ���R�6�px��|՗���������
��PxK��4K=�3XU�:�Ԭ��)����Oq{:��oB��l�U(���f(�8����Cw��.�$�}e\�������:��_R�tV���Uhn�`ꎸEp�5�<[npe�y6��a'��ڑ�B��>���!"��&�}�?�RՈݨ	�I�)ə�3Z�#7~D�uJ��6�i�{����b��_��֟�(N�<;��sY5����u2�Ŀ��b�	L�_%��J�� �u�J���FL����{x�P�G@�Fz�V�V/���~g�]���3VN���#���%�R7Tf����{9���#�ܭN��Y�àA�Q�������|�=�2� ���L�C��̉hG�@��Y��C_����L�����S6�0���� �4�����ӊ�ٮLYɷ"7���}%EG�	�/��/q��G�4�����?g�p��[Ӝ�=jd�N�)4��[BVL���$[�w�����M��^1���<�r5��5�f3f��	#}Cn���d�'�X�O�����D)	{ʟ�눺�}�\Y&%�^���L�۸��w>�s"f�T��y�f�d�gU��.�>����-�qS)̦���>��C=P=�\P���j������Rj2o>��^��u�k������$����D�F���t��d6�@a	4��~)����?�M��D�N�)�͹b���4��mX�L��\��ٗ[�jXU�h��Z�wj�獩Z��x�e\�A}K�����-qG��,Y~ȡ3p'>�����.WM�w�v�3��B|��`͚`l�GR���@Fmg@���� ��t�\��XgW�Md3aH��6�B��!���g�=��8�ZO�ux��)tI�%�9U���Na:� [
+C�~�=���T��J��s������ti�x.7I1;w����-xĨ��e��C��='��Dx�={280<j�гH��6e#��5[U��Ĕ�3�-���+�o���PQ�s�O�ŐCu�^��f�2�m�(>q��(����H��(�z��L&���3���Y ��#N��(<oȔAY�V��3�e��Y�S6d\��V�/ȯ���ק|#-q�@�9(uPC�  �-��2C��dn��9L<C��t�x�eKӡ�0��IkTM!�q+�
4\e�8Jg'�u1ٯ���x§��O�P�����{��/�b���Yj6�>uG��0�ŢG7,�>R�f��:�('89��R)�\�J��F�
���^��;�C�����Ӊ��A��f��6�Yn���G]C�����ȱK����<��U;ݢ�D��/y���vw������ۿ�?&X�Rڮ���-���
�"l��=P�ܳ+��P9L%Sv��e����+(��l<s>'��c�*�rkb��N��W�_i��]��k���/ai'�%|���ū��j�"h���hՌ��SCPT�s��d}_SL撥u��F6]X ���I�8���Hk#t��Ƌ��\�1P�D�q���.�� ���S![Sʟ��]��`p�[evo��1���
G�2�V��������6��M��
Cx�{�Ñ߿a�{~IǍ�|��jQ���Jx�w��A+�[Vއ�~�c�*M���l��%�E � �������_z�;���2}?0�ӻ�3bH�Hf�	q�$}�h�c[7�*ֈ*+kJM6m��H߰ �t�ӼDS�@;H!�1�� M�4���Ɩ�S>�W�\(;t���]�"#Ɓ��_@��]B$���Y�,�l�j"SC���=�F(��}�Cb�z���)��T�b�%���ݮ�F���=�Zt0�C�G��{�F,�ھ����7�P����h���_�9>S��=��!����G���Н �[%G8Qg~�'�=i�9�,�ꠄp�k��@��{f7���l
���hj��`��Q����/��!�aZYa�oA��i�_�3����aO��6/ 튳�򡤎���_E���jBR�:V�_s[	�H�1�5���[�� G�4�n��.9������[�b"����+IX�����q3�j�~@�����(�Ɠ׮M!�E|M<ly�
+d�XFM� ���g���>9��lR~W���4B��=Pd�H�3@�$�g#�h����>ٖ�Â�����m�Q�Å�������g�G���|p��z��e�н��M�����7�G�ͰzK�x��_�}��}�� ��K��,4����nm��HV����1���xu�G�3�9 E�mmr���uPd.��8��
�Qؓ�Wŗ��0/���Y��W�\|_Q���'�K�دϠ�К!�X���?�[�+g,7c\�AC>�yE��>�?��V��>ʭ�5Q����#ML�n�������Q3���P*�O����������a���I��5&�K�Ҳ�o�2`��6 �ܣᾏ�3�i!]�r<�p�����I��迺�zU��̶m5[�wv�A(����Eq�r�Ζ
k�i���q����ZI�܅�@�1�u��z�4k�t?��I	���R�2=�Y��&��9&����;�8��=�E�P�|/bJ�b's�yR�ɟj1s���?���7�SOG��|+j��ԁm�s��N����L��m��h��W�v��^%��y(k�i��$�p� ~�m8W���&�{A;��2`�w����ed���5��RkM��
���x��s��X뻹���夃�*�\��ϒ �z&�K�-�����[�/�~���ع#��)�$�� �,%<��a�Nh��L��<c:�B7�T�����*	����}����o��d�7��U}�5�w;Pi	˥i��,�'�{&���3^�=(_�$����B�#��G.s��LVoʓH�J�ɫl�Vq�FAv̕��	+sCc`�|����
X`M��}�I�x�]@��˖��x���o�����a'�X��!�<���1��(�/?�u�̫׿�8?�Zni*U24Wf�:�R�E�3��&=���!�4��� @�6�V��DR�v�C��ca�$��h�J�V���~�	��J6K̜��D���Z�� �5Crj�љ��!ۑ1��`�M�e}���K�f��1�ϳp��)
��*s&Y�/����8�8��^�:����y;{i��6b�ԥ�g�N]���N�G��1����^}����-}��&��g#l�hM`�[ť�:î�x��g�b�!#2�� a�K�Jsh��n��Gr�@�����Hi$�s2 2=#y�_a{X��N-�lJ�k��I�ӓ���<{����:�K���#.1�!l9#�'��@�F����I�U1ҖH9j�nQ��&CP��}>	O���c@�������F�"�PB\j�t!�<��Q�2w<t毲�?}�{|���/m��[%��I�5�S\�{X}�_����D�	�0
�ybW�\�r�5��.���C�?JV/��<�ڿ�<C�&9!�5b5
�8�wi)NqBc��<�V���N\΋�\@/f�3=(�^Jg�aԋ"�9-��>.��E��0Eg�gI�� HN>�w"���[B�#�"q���w�Yd��`��K��;�iK!�'�H�������<�׻�"�����2ۣ&\N�	��vB��3���MW
e��7`E�β;
·6����H��c�ѺB���]�E� XsQ�.Q�`�Kd,�Pg�湍:?O���I.��n�	��VI�2�v�z��|������'�o����], vè��[�{���||F�{V����Z;��lk`5����n�%�.�)g's�9�����6�U.e|��*� X���t燘E��Ȉ�"ؐ��J���T��vH��)K�"����З�rȾ<��p�[:�,lb���}�[m(rpʊ-¥f£��KY�ۭNK�ι��C�IF>ֈvo?2n�:� ��=k��f:<��½��Αd��$?d4$�h����^�߱ �I!7�=���������p�&��U��J&q���"��2"��{�P���N�:����Dߠf6�!0�^K�̞Z>�f�Y�S`r�FVy��M���w4�;��;�i�#B�/�k:��۟��2$!�H.AY��F�-X#}�kFm>�)�d���mVm>`=��\~�C���G۱T��T^��H���Z\���B�޸�{>���G��8ٓ7i��:��Q�MhuP�wE������k����Y��i��S�G�ސ�]N!x4I�?�)��md��(��I�tR��P�EW��ނ������i�ơ������؋��V��-w��O;�������(E�y�fi��|^¯0�2�F��fgl��v>ð�[o��jF����*:�KIE~㵝�R�n<�P��E&k�}l��	5�j�� ��;�E6����8f2�Ť�/0X�T�bĹ��� Ԭ�õz�u�V�'Z�J&�i�+�$��S��y�<rZ���a߬�n���S��+���.J���7}9ƺ3+�,�	:��-�6�_A��;dGeE������4��Ei�"[��6���[���d�Jv�x�������4������>�2��-��*º>�v�ӷ3 #�|�$Zbwʲ�}�`+�G���U"�<F��4a�^��/�X���k�oi�O?,X	�-aLy0k�c���|���w*����I�K)ES��s[%�ջ@���+lLL��rA��\*z���m_�gA/6��/�q���'*�^Q�LO�[�𽞩2\����[���^���q��J5>[puz���-}�6�Dθ���d`�_�Y�3�g}�����+%"moZ{8�
'L�l����8�S��o�j!s�!8�����&��;Gt�jǫŗD8&ȃ���F˃D����5������}�G�{날�a��R�n�G�m�	ME+>=�]U"m��������ݶ��v�|w��!;6P�y)���		�Ǔ����������&;9a�G�D$ ���K��[0q��mn���9��1�Bi�L�ߨcX����Ӑ`�Oް?���l��)��2V)�����~��5\d,o�������M�����uD����h�������j:*ͯpR���l޼����T�:\�R���`��ra��;]!��sP��U^Sci9F��J6�F+���,?�R��Cg�~˂/�t�9�^�[��D�&��OY��5/Oe8���"b��F@�؜+#�[
?I�g��D�C4+if�X�,$}��g)�gM)��ì��* �6K�$�=�����͏��ۢM�|��:H��Od2kCI솱٤���q����Q.ؠ�y`]O�K����<([a���r�t޴rOk~k�n �,U�$��߭��c��f�� ��fz�Y.�Zb�ԟb�A��&O�Waҧ�g�i�% ��#�޳��Ǝw��?��ȅjX�#t�,��@��C����t��_%�r	�ǆnT�,���N�7��S�5���J��ܩè���D�y� �������ΞQ�a�������]Q��p��r�oJuH����%K�/���1T�Rp���p�Sc;)"TO��<��T�F���7�%Q� r�E�ҍMl�p���E�("���c�����x+~@�x@��#�gm�l�f����ǐ�w�K�MQF���\ϫ�F�h�keWE�C�j�5$�N
@�b y�y4�6~���b	�^Btx���䳧x�qﴍ�MGuN�}8�%-���[[c�{k��~="v�j[����!_�1��S[ʾb���$��f�hԑ�Mi0�r�?{I)�g�l�{�!Z�8<�#<���<�]�YY�t�2�E1�o������=�㚲(��L�δw���{��M&R�M� ��\��ힼ�m!�g�j+(2���@�.�`¹�b�}��^�o���< ��b����L�h5	WzQx�/���m��ž�b�2a�09QB�"�O��~�x�	� �>P�!ԹX�o�sm����v�}?�d��[�и���M_�g<,�ڝ���ؽ_�,�����f�
�懌|�|��Q���Da�>��['�+h#)[�7��������uC+�O��0l����a��ʐ7��^�/�9��'��اjS������E�� ��)BF��fH}�q퇹ƖC[f�u�	[��BsF��+7mW��3�\|*']�]���d1��nُ'S��������"���w%���x�d�f	�=a҅�d�
�Ȝ��^>�kߥS�M 誣�~�u���{8_�Vt����X�X��/��Oܕz�n����C�3�k�Zmܭ=Q�`rzI�"s#:��Wa�~���%08���S�'~�_!$3��f5����p��6��܁�CM �m�G�u���>s�l��C�9���;O�}>D�lzd�W��jO`�����t'%;�g�/�JUe���9I�cT���>{젒@��j�N�Xڳ,~ ;m��a��M`S# u����e�_��wQAxOҐ�6{��r�����J�M��i������_
�E�ʐ������Z
m��N�luN4�_.b���,�aF���/������z��"��p
o�Y�[�<�D��2��զ�0�ѵ4 ��˪�p������㨗�i)���Kwt���*.F�f�8 �C�Tt�"Z%{Tk`�#F���0�J���F�L���T8��ګ�d*(<�rh�5Wj��E�&;Z���젒n�xH���\�Z�^�C�#�y	�N�b;�#M��/�	yj�q3��F<T���x�*��B�}��xf\ܼ�5�p��lu�K����#�Ő�m���:^����n����>���_V�0�:��#^��YPi�={������ڷ�'�C�at'v�����Ά�H�[�C����ŅYN�%�Ӫ�ٷ�A,b����nZ��>8��P(l��IR�U[�\p¾�?�����f$_)߫���_'������]�2ĶJ
�x������n�H|=�+w��^�kJV}�*����_�,�_T;e�w�e8��G�pi]pY�8_�3g��&?�Z��'R	�2Y��> g��6��,�D.�$����r�_��+V���kE�N�Գd>l�����tW����u`�?�\L���|>F�jm�ɻ�k󪼖�Aʓ�`�9$��3��(�|GL�8���`	�ݸ~w<����͠]�=���+k�?��ɒ�}�+|*�ཾѸW�/�΀'ν4�������H5:�E��v��r�B��x*�L�Uv c	X��ĹҢ��ء�9�IHb��gf8�Oǃ�oO���1'N�$�?�Y>SV%��h��
E����<;�4��n��7FOH%����k�ЁҜ�V�!�ל��{2a�E@"���.���K�V�ݣ ��J]��[��D�Af���(s�>ڙ>��ߡա�k��c�i�4Ȳ)���A$�z�yR-����0����5�d�&�����o���ɇ����)�����ҬN���`�Bݿz�aml\]���j�I�ޝ؃aW}(Xy \kq�N͸H��秱5���������s�T`EAO����WчL7��,o�N��c��T���rZ`��9υ�dO=����e�#5�AM�9�'I|yXH5�u� R�ކt@#��âb�� ����=�^�Z���O#OoUT�x8ܯ�[�ofS_2�T)�lj
Mh�欧���)��\�V(9lLM��[��ϛ{4�����r�<�cſ�C�a�G�p7�L[ɜ�u=ځ�e�~�*�-jg��ʎ� _��1\��a]a ct���#E<�r �4�l��*���^�j�"��C��g��g�����/d�?���攽�p|��>]��?!_4����s���L�5�+Q��l�ƽ�EfA�b�5mf��;2�N*�����Z
�P��D��#1������^�����4('���t����ʸ���6���m�`S+������WYn.�a�NQX����v �������xU��:!�Ѩ�+ze�q�FW�$qVG�}\$	�N칥�7���O�ܘ���x%3W�?��6��D���k�	r��9�ﱯMN�IE��׀�Z=Tu����tT^<�0��x� n3~Ц�ƏU��]:�R�;/�U���^f��0�)����.�M�Y�??W׾�/iti��]mF���A�nŅy6!�.l��F7
t�R���?Ԝ�۠j��V~�P�7(篅w�MX���زUnz�߬����V�h��gB��<��LnB�pO���j��YK���:ǻ�m�y8���P�P�X|��?>e�G04j*w�nV�5l��
�$R��z� 6���4~'�i��Lf� g���y�c�*A�'��yb�v��4r������_L�E�Cݷo2rd�'�2-�)'�h0�b�m�F@-����>/pK�^�]͔�8/F�l�Xp���\G�҆��K�c��_�R����o�/^�.m^��4�f UO�3	�!x���t)�Ck��$.�zbJ�@�\���H�9�s�b�G�����R�C��şFמB�0��u!:���6@#�sEoػOM���n��#�C��e�ts����۰�xO ��9�+ٮ�a����~~�G[�&k��Ͻ�^ٝ���#�,�����ݔ����{ρ�zz����5����a���|M�;��2&�pRw��ݪ�����r��j@���e��s/�3����tv�����3�}���7O�N*3�flN�n���ac��;۸���+"�Ԝ1�~��1;�)\�\ǂ��+���oE�֯�v���ӽa�ʜ�A�f��(�}Y��z����ɳ����绾|�s13�m�i�Dɰ��c�1�Ү΀*9T��jh�̲\V�'�*�B���y�*�c�=Zq��Rpt�t15���/Ub7W_Kf<h�^t*]���~�[4��.XFL����ª���I׋O�r�3i��9.��Vx�:�����ykt��j&l�FF��Ϧ���c��V+W����a?sR
a�~AU�+1�[l�� �p�2���e�ęZ,nq�yi��s'J3�K�"�@l'%���,�q�cB�-��ySk�8J*�#�t\СFC�+c��f�Ns�^�%�	u5�, ���]m�-�~vX�:^}��� k��1&w[�+��N~�~���,��Co+������jQ�rju��E��i�O�a~�7�"��
:<BBB���E�m(���/���c��60\�X�<���b���tG��onALUi6iuW�������'�a��U+�\������KOHL��F��o�j�[���ì��8�Ia;��XB��Q��(k�m���a!L��.���"[�0�	mr|��Dh!�,��0��Q홈��@@�~��E�eo�P;Z��/��w�i���>�����vp޸ӟz=�ݼ�z�Y�(���=B��m�@���hٞ�b�a?CϚl��r�f#�]hЯ_��uh���c��ˆ,k!��Yc�ź��X���7)��nE�c��/��� Pҕ��m`�["�X�P�L����޽ ��P���|}g�s��b�Q ��z��^h7��j!?��x�ː���B�e�0�*B��f/���9'~b`˼�a��ۉ%rb=��O�װ��d`�8�Bb(��W)�Vz��h��2�kMK�E�*��[�V�A&-���~���ۗ~w+�*?z�s�]jK�������;�ֹ�r�SB�X�]��0=h�&dSnV�y;�~���$r��u`'�-�DZ ͈LY!���_1��꾛�% ��2��?���R��H3|ȕ��ػ�l̀��O�L&����h#�?~��8`�*Ԑ��B��u�3����^�nx���xD*8C� S�[
���R��!�۟���;Ν�����&����e�\f�h}�-��K����y|�0���+(�Ϲ��ٙs{k1��z����� ���
�&�X�y�E-[�}������NO=qm��m�Yu�CTzAXO"�fk�K�馞*�qk	�44	��(�	��2`�]�v��u�:69٭�:����̧G�N� ۄ���Lø_Ra�~�� �9�m%gk'�1g�kz�tB��a8�~w��Q~�?+�2h��),k`����%�"�Ie��"���x�pSڴ�����d��k�b�l�����д�CQd�uK�����$]��e~�+LC�菓%/��pD�>2ԩ١N�T��f!�~�V��з���z�M��7^|tc;���7�ӦJ�hB���l�I+�����nm�Qq��a5�S�J�<mE-�	K(Aq�ez=������!y3k�z��m�_I�F�~��u�.Z3ԑq&�{>I����D݇;�7b81�A�%S�S�����?&�\vuu1L��ԃG��֑�Y�U�nG�uOe�� ��U�z+�K�Z��l�}GK���e��yAVË� �,`��_cD�뇧�X�w��x�����{$��X2�$�#��6�0G�?�7�f	C�mj�x�yao���^��~%�O��i���9eV[�����.�`�n�}j0, ,Cp69��Xb��#m��Ё8p,��Q�ۆ�pj����z���Z�	 �v�*�8�[)�k(>D��Sǭ��ʮ�>]"��C���8L�t|e�@6T�G5���5S}��+o�[@Y���P�]��DQ���n%��M*�$�r�I��Ff��<X��Byn�}V�*�oi(`��J�%e¿����~4g�l �2:��53���)��f��g�^I5��_f6�:,P���?�-ِ�l$�ڪϬ�C���N��V�J$��;%�
;F:�:E7��<p�2Js�4�'�Y7׀v7H�F��������+@:�����O@'�1��)�c�^���9V��F��ÚM�2�����k��sO�ٚm8�����0?�)\v����w�A��iC
k��3�v$�g ����}ؠ�^
�s"��:\�M��>��������ٿ�^=RvځS���ߥ�LjJkf�	��HA�ח�ƛ�`�{��`ٗ��a��PԬ�D�y!6��1����H�R��Ag�����?ɆDc��?������w�c����C�1���@_�-)�Z�)��c�7SnG�Ra5�8J�a,���.�m�*Q�wd�=mE��U�g�v�u��OJ﹦?�����Q�i�E���#̨]F��"�K ��>�LH��-�b�J�|t� �S/�ʱ�d����{kIY����q�y�~�>�ݗC[`]|xZ��0ؒiO���,잸� �OF�Y�+�s������@�����9!�,�������46�����dP��R���rڔ��͒�Y0[�9�a�����`��/�jD��n3/����{۸�����/&�m>�~EƄ�V�Y�ѫ�h-��4F� ���M�RYU�;`�Z�}6Z!��v�e+I��g���W%��%EU���W�9*�\jz��ƨx���0��}4�xJ� ��	�Lm��ʙ5��3��ۀ%�*��h���8�EH�ϩHς�m����Ck���0��g�}��%@lQ��-���
���TU�T&���Lf�Ba�`�����+`�w����ډ!]��b�Q6�I3+[�%�K��
Zv��U�`���Md�2A�Ͼ/0���a�s͠wB:f��q�"�E���V�����/�\=���V�p3^�Fι1i�vC`{3N]����\�k���;��,ׁ�g}C�Eyh�L1/3~';X�(�	f����9�_£06�p����-C=q�Rnu�d��z�kʬ�~�4��@%���������L����Vu���#M/ۊJV���LV.8y����_�e�����Թ���=*�;�r�58I�R�*�a��$��n?Ân�0�̯?��ؼJͅ���PQ��]����M��q�.�(P��7�M��$��'|΍5�����]�{���B3DҖ�ц����L��rcAM��q�ӄ��:+2�ߌ�eX�i��=	��[���l��kvLE(��C�5�g_	#�%䷦�u�Dv�YV�{)[�2��	�
)�M��e��"��A
�Qz�L���h�B̈{B�-+B^�x@P�5����lp�>�y�
��+�����=��<tFq,��P�̬[~�`9��v��9�dU;6�n�f��d�����C��@���.��y�;�Q��f���u|{%�>�7|'�A=&'6ҧY�ڶc3(\��� ��n�M���=#���qsʦϖ\��t�-��\Oc$&h랋ށ����5���w�+V,��L�C`w�lMڢ;��{�aA�l"��w����ٱl�C�[g�Y7/�|��.��ϕ�=�I�i��e��'�	j6v*���x��EF�*2���T�y�NZ!���_rV�@Av��OOLD�����e�,|�X>��G�Nk_�K>C&İEJ[簄2ޜ_�Q�F���W]� L���?�h�w�T
�����F�g�y��s<lc���;c������ ���d� D,�k1���"�(�L*!2�q�v�N��P�H?⬶�6�ei�e_�������,�cٝ��`:����$lY�t�O�9���ע�,ŝ}N�ڪ��5�D�%b�h�yx���|�	E�&.��WQ�]e��\�~���Z�*��u��=7����;������NN�U�VgzDɻ���X)e��D2��'PT�i1��˱1{���Nԝ��v�:ҵV�XY�b=��#<������K���<D�y(z&�]V���K(Td�����&-u�S,�T?�y�y�榟����S��JUDw@[���{��o�v�5E����@Z�f�#7v�_\|c����Ơe����4ҾU��>Ny�X$�e�ѳ�9�4,&Y�2�"V�e��{3d���cB8w@�,�mk��j������ȁJ͸O���7[�C���uL~9�:���d"$����Fq�'�ʸ�؄'�
����M +z02�NE���<�	r�y>�6�OL�٠~:"W@��;k�+e��ww��󵦣
p���:p��?uGŴ\�H�=����re��҈)b�B�-7��I@�IJ�|�A>I%w�i	O�� �%B\h=�s�wU�Y����k�ߑ��,���X�U��I� �x�������.b\z��4�`�n��}�v���fn�OHg3�L��¾���R�4�EI�5e�-�������~�T��_:|���(RE"�Z����Hg@��b���%t�UÎ�7�>L|
�l[+A(=,��,��Q��k��p��mu��T?$�h��D�8��Q�'BI׽��c,�m:x𰭖�xlm�l��:׎�'2A?*͝����ω9dԴ�&�wt�Y]Z�}ۻo�ք�_�.n+����W�Ե�e�?|8n`��u��� �Z���M��b{�N���Pf'�}�2iD"��Ɗ'Z�P�QЋ5�/ց�SaD��_�72Y�4�C��|�%&ɡn�R�H�P:A͉dS�A����|� ��AZ���VBYtR �*<�gǓ��a�dF׳Pn\6��*������oWhL�M
���u���r�����u���$eK �ٝ����8�@�+��ZlɹT��� ����9A��Wb�Mz�Mt���J��a�D�/�EG4M��$!�\(G��&f�
.h�{�#I����`�*�49�N����hѳ�������SZG�k���/���q`��c3s�ЄB�:}�,�8���Q�_4��ڽ����AXh)��31)�1�!n�qm��5ӓ�Mi��uO��â_��B ���9| ����g?��{��(�4@D��۽�"y�=��бƴW����>����8�z�*(��X$0	
*�0�%��3XɱYi�N��h�OB'bf��}А9��n�N�O?��I �T�^�+�,l�O�Dx�s�DZ��S���,�J���r2�K��Y�=�J�墙�f�"%�66ѓ�(P��q�T���jdl���V��Uf�Y�J	L3c��C=��������*�ͨ�#Q��?KV�$g�2 ��율�����3x�n�P�DQ_X��&�d�~P�=A���&�!XJ�Z�VG��w�@�R���c	���
�ӣ65,�nġׁG�R7�*X|�̄Q4IlW;n	�����Wy��3F����gȓ���7Fk�3��5�,*=)�)��P�*~��q��p��@�V^������^��`���ba��]�{f�l��U$�a
�j��K�
�E�*<��qR�vFqKk4�Q��R�X�e�OP��z �ܑb�Q�]�է�%�����#_)ռP��3^�:3�2 �c2�5S7��CM��f�;�"�wpU��Y:�(ޡI��b��v!B]8���-ܣ}�dT�f؊Q�$��C�}1~4<����S��SY����SM�-h�x�i����9!l��l��P��F��4w䗾�]r��=���d�m�zP;|޿�`���@��5WD3�Q���z���<�2�nP���z4:���Sa�o���<*'&���K
��bb$$3�
��*)YS�0B<�?˥�MJ%їoa�\Ņ�JwDɥ���9>Lt�����c�*l�v�")D��n�/����l���ǼL�������Bo���G���?�Af�w��.T�݃����-X�#Sղ�O�M����%rs��<8E:���������y\�Ո��fa!.��,\�9���[�|F��j<BW��Ʀ�F��g�g;Q�f�A6_�h���㕤�h����JfM�BR��Ax��3綔]�Z�>�&�̼��'�����	 �9C�F�`�zI�(�u���d�v�_vܸ��;��&X�/)S,���OZO��u�3n$iB�`�^�3����|����WZ��U��,\���ˇ��6���8��c%�h ْ~���,��4�"�����ԓ�˰�i�Lj���qZC�Zq�K-��M*S�	5��C��]�ZC��.���Ķ*�"8���{�C4``Hj"hs�[���9�Uw�uq% Q����\�55^'h�2�V��NT͟K�5c�=�u�y-Q>�Ŏ��r��0���v^�Jx)�Ds�	͉N�6k�E�@:x�*�~���|oQ�=��zQa? ܨ��&�0"� �^Tq#X0xn0�і�MN��NZn�:�8d�B��܅����مtZ��:[�&�7'گ��pa)�̷�sH����-]"_��p�^��o"W��~��@Gl�#"��B�q��t �	�Jr��La�/��U��b�O��FF'��խ2Я}�v��c��kP<Q���Fp����PE�և���h�fd�h�8US=ꬅ4��W���r����",�T��%�Fm<k�'�$��O�Z"�&����;	k����M~
p����'9�t�;;ry�R�b��������5��K���0�n�D��A��)%�!����67�fuܿ�����F|�D
��EfR ú;)�Q	[��j��=��GŌ� _�[j7UF�3�9�����$B�[�� i�~�v	\� ���V�|�B�`�icyj-�xwQ��@����7�� ��s�W`����a�a\��~�#���#�}�g:�X�֐l"��;�'��*�10�IiV���I�_�^B����8Nm�2:�֟�QK'f�A��������mc�I$V�M��mZ��g��rC�B��x=���nK�[�:e*O����&��W�Ǣ��W���)0,c�&�+��&#Y�QZۼ��8��qfH�Ύa�C9B=<�BglQ_��G�j���u�GxM�8E�l�M�r�J��]�˘�uC��DO����ҩK��by�`7��r'��E;����c2lU�����q��D���$O�
���ۀ�f�t�j9$��Ƕ<B�Gl`�@�){� '��59Dx.�A{'cB��_�ė��B~&!t['Ã|�Г-����i��|���ػ�K�w��|�/ja<�o+z��u�s��fGi=9�.�nN��gH%�3e���Mb���$#�w�1�=f�+�0��0��>u�y?����A��I�?�'`�B������hI��]֨�<����uSK�LLJ�`R�ZǤ#�¼,�h��̨�+�\���2?������L��~��Q!�fٳTPu�}]��BQ�3Ĺ.7�JD��}��7S
�1�y�b\ޕ,)���w�f�Aʩ
�P6�(!���v�1�q�浌��<���5�]T��M��{)٧i[(K����&�
�(���
N�+�QNW�y7-�,���$�v����U�Y[��ScQ��(�j�3Q�~L{�-��m7?�u�����9��Q����1��oa�\T��؉aӄ@��l��	�vaq�3��N��{�SNOչ����M����R��m��cB6\�\�W*u�6M��@CBJ�\�&�'t{�٩^plC�����yԦ�ɟ7����k��a�K&�/�� �&�Ѹi[���o�:E;�p<eI%���'I���;�Y��C�׆Y�����r����ݾӄ �	S��y��#��\�0명/�z:�_�� �:D�=�R����Ț[����f���	�.;�$�a�E��+�w\�
X�	���N�P��Z����[T	�po
v븍C��ܵt��kGQ�UON<�?�p�&��WGf�R��o��K��䢕�_~,����8��39�)����z->@`ob:�5��-��T|4��T�Qmerb�"`�z�}&�C�|��f�_I�����5��������q-��8���+Z��eoCE�<zƺ����%����=�4O�}��+/0�� ��ѻ��K4>F�u��ֺ��	P�V��7^�K c���d��o���o���� 򓃺8��o}R. �<	��>W��C�t����n��"��^��O����T�f�#�].�>��/_`1E���-Gթ��+�{������Zx%Pi-ZE')�m�x߭LױB��ދ��~=9vZ�j=�h8s�i��0b�� P��"����kD�S�i[!~�1bU��0�Ͷn=N�A2_��LTR���)Gw�g�Vʈ��D������ĲL���6���x"�+'�ni���̓�x����~��&U�2�'�,���0�4��ݱM��dH�?O�?堪7s؈) �M5��u�J�Q~�+�Cp���:�%>\3!E��X�M���]E�b� �4!����ڴ�|�9j�A��@RP��E�����@N�!d����$�SOi�_R��$�<<=3��SrCQ
}Ԑ�Eh�'9kr9M�(~��T`��$ش��&���q�����X.ȰX�Y�dWg��gŊ�+Dr�Jެ�ܫ�K�4T�t�RzJ���s�Ǩ~��Z53�����b6�,4!O��t0 6Զ7�OP�m�W+D��� �7�{��jy��J(����c�m�
�F.Gf��塑��I���B.�SJ�f0
t����M��,��k�+y1#�F���nMqXg�oV��P���!̯�Z���G���?8�@I���"[3��ԝTf��J\C����=��0���=���Ә�����!�u����׈}F�M�͹c��>�y�x:`��S������l��m������珺s��Խ�K�]���j�=�e�	7����>�h��"�F�/�#X��.��ʲ�r0$�N������#����ԯqW��nb�0A�i{*���僶���UXN��R�K��F�w)�(j	-��d?!�/߰��q�rSP<�kȱ�h��<�zH���c 1��N
7��.��[y��
 ��OZ*Wf�ZWพ)_�������W1�]D�q��$R�=H���e3C7�So] ��h��!-̈́E������S�ԁ<nh߸����' }�����<��Ι��%F2�-G�7��������K�!�=�ϹfȜ�h�E�Qp��9X�n���� �K�m��ݳ��k��v��8��J���K-�FW �����'�;Ђz������.���c�c�۷��n���)�9���$�T�V`��x�B
R%�K{.ܼ=U�MP,��J�eG���4:Y�<��Y����\�MY'���ErE�R�f\��
��
���w֡��f�̌R27���#7�J��Y��>aٴ$��(6�>�6�I	��/����4	��-;��2�Z��Y�rs��_Y]��x�pg�褣�ט�n�Q�)?y��`�x�{���B���F�`����9oݲ0~4ɬ���|�����F ?�ph!�o���☥��D��b��6��Y�5-L�v�Bjs8��%ߨV�� ��"��v��6�g��[�z8@^�AL�ڨ����\%{
���-m�4�����c2)���:�:�����y���k9��݌���?2�S�#�쯖�n]O��}�����LH�t��(��/��,�R~40c:X�c�z8��z8�`�G&���._���f�=�27���l���7�p9�Rq��xK,�5!��6�8���3�j��7�`Z���&�w�qޢ3�ē���wE4��B`�R�3��Z�]�H��>54K����n@pɗ||Iv�dzh䮫�������1�]+�U���fr�>A>l������s�1���F�ai�z8�֞@�l�/{߻cf�N%�U�H1�#�"-�M�+?��d�D���y��僭r�X�Mh͌�3��a�&O�\L�y<5�dA��� ��A7Md�H������	rGa���X��h'vu\@Y�Bu�Ǩ�
�^����Vo관�������"����f��B�:x:M�z���o���g2&`���N=\"� ���:�J��P�:��<܃+��f���V���BHy�,��[���'+���9b�kj���ȲA������3*��H1�j��g�	�<Uk�R���n�m�v �#�SYK+�St��k.f�6���n��C��j�m��~�2�G���bГjkQL��t8[G��a��q����00�������"G����.�j��~�6;�$��Ąd_AIфP��d�1l�C�I@�l�ʤ⛶����(cu�g���L��tr�|��'�xW�XFD��-a�I#`��d1"؁��2�O��N���y�c���2�],�d[�:Vۧ���"ލ�'>K�,;�%��t�&���?�!��1�"vW/C5ҦL1D�r= ~�3z"�����I�n7�!e]ޤ�T@��,���Ǡ^MD$�I��?���z��N�����g�����˦�(�htZC{�C=�ήF���ͧ\V��VVy�ef����?񗓟���d���3D;���k�ɖmHӶ(�	�}]��l�3�l"V3  �k��	PI��'6�uux;DWAF�8� �4�꒻�t������7���W��*(�Z"��T.�pE���pS�H}Z�9�EF�{l��V]ϩLʏ��$��|_?ᕥ�x�l�V�����@�2�jd�����.��h�� ����w�`I�8j:���o�W�'X����W���ᆌ	N���;����:�ə� <�K���mbR�L�aۨWe�6�gJV��`��f�v8A�PR�z7��D�jfXV��*ʠ�`�w��45�d�5��܇>:��)��xyؘ��ν�Pcܶ��_Ҭ�8!)r�� h<>ѲS��m�Q�.&]53�ɺJE�Z�z7l��q��z�8&��RcfV+ݏ��!� ETZ2SR��,_���#z=�N�r`����Э���%L����J�H�w_���D��E�?�-R��0�̈m��WLyY�ަh�
o���� eS/��ao�XfB�Dgw�맕V݌PM�)��|z[}ǒ������&�����W;�E�	5�B�Bެ[�`�N�4�DN�(ֽ��B,��e�<n.~8�Bi�Ao6+Q��įI~�xwk%���&�����^xIk��P�[OfPޚp3g��t�;�̝�c��D�lC�BI*k·�����%\���]�^�>���\���J
�q`������'M�)j�|�ܺ�N�ox�6G��@B:S��+� ��ಣ���:��ݸI����`��M6 �2�}�����/^9�.�d�E�� �����w)a}^��0/B0�~h�IFˈ���I<���	)�� �oۻ�C�9f����鍀vS���o�n�Ծs�B	6>�^���?�S�g_�w�C-1ϋ�˨b��&�>�@����ْ�����,y#����Î�xҠ~�6<[G�7��؀C����p�K�O�8�{P��s�ޮU�7�c�dd�אކڜt�X�јT\�<�>�MJ"��������-��Zo@�bhO�%K���/��`�i)f�x�6�Mx��qs ��B�A�_��A`��+F�Pԣ�6(�I��ȩ��ho�I@�{����|�{,�Y��M�ҝ����-����fP���'gb���8`���yq[����(AP���2Q��@��z��WG��X��^�C�9P��0?����	�:?���ѻ}I�VԩjPŃZs��[*'��СC
�_*��@��u�dC�y��.LA��m`�%`=��K3Q�P�Bl���\J���H�`�;˼Ź�0ٸF_�[��% lxB�˞mչF�j�J.�ܨ���%�&^��M�ι8+�,UkDy�J�fD�#4aFf��K���5��y�b���A'MX�A��_;ke�$���E]͎ AH��oҼeҡmk�}t���i��>\�\�~~%l�������[@=��b��'���ȍG7a�8�J6bv����bud�h�B.����-�r�8��9k�My�1 p�~n ڶ�'*,�)^�K̋�'�5c��fo�NmcR�L����pk����D`Q��׶�}�.�~�.����\���D\x?�cR ��I�t���w��)e�����HD(�k8©�V=�ҠH��N ��*�R�C�ߐ&��ьP��×<��ڿ�zͳv.��KQ��2�b�K���詉7��S���RA�&p�-�y�J�����(�6~7`�I��"�-������ڹ��>����C�<[853��/%_u�^��K���Y~��A��Gj`T�0|��Y���Ry����{&��+����s�x�!=���a�é+�{�SW�/Y���c�C�������k��<�8�t���	�����2���e���T�`��ϑc���'��f:ŊS�5Zhܻ��9n���J��������OO�3ʿ�̇C:�x�l������{w���n"�M���6և�=L��'�>��,�v�gIQ[�N޻s�_�3����g���h]&&�<u� ��@��^a-���/C)��cj�p��8�����*G�����k,G����c��op�� �-mI��@����z�� b2��N�Ɋ}y�J�RA�j��K�~���ZV.�g�.D16��5{�>�;�&������M&�u'ʙ���V��p
��q���23Э� �����r[f�D#l�v�	��g�7	�$m�X{Xf$O�� d$_\�(�/tT]{�i�*f��]��HKB%��aTP���>k�Ļ�A��E�o�ȕ����bz��7r	��Ř;' Ti��B���*%!u���Z�>��B�Cʧ��&U��A\��4�����|.��"�a�5jV2[�+r��**9�t�OZ���N�DP5;4���ސ����7%�:�br�Ĩ���(	��(܎mf�ѳ�դ���B	������!���ml&�n�b�_�H#�$�m.k_n`qv��'�����uk2�cܡT"$���ex�~��	[w3�4�h���d/��@?�	5.+�<��y��L����0����f�Ly��Y���z	��ݺ&��LWR%�y;����J#F'qN������ގB$��ّ��F�S���nz���qV���V2��W4��%πߪ	I�'۫�Z��������*��N�[��;}B-��gɜ����L@v��0��{=OT���B~�Bb+�5���o{V��:��N�y����=�e��}�H��}UY�\�ě�����$�t7���u˒����/��19��ԓ,VǭȦ���4/Z���	��g*ғ�ېC�Ru�՘$���"X�Gw��2�!oA��\�~|�>��P!U4������h���@[.Z��%���� �M
��"��P�\@X1p�]tA�����OՀ�������J��`����ƻ�������lgs��V~|㏽Isь��a�}Z��(Xƴ��߿k͊��s�`�F/�
�h�m �hl��"|�'�OW>������:QX�7"��`^�;��#�se
�x�ԫ*�Z\����D���-�'�SБo	>o��ۺ����}�Kkl�4�4�#omK*��b���ׁVT5����y��q~t������e�xۗ��5# |��#{筸�	�����+�Kbw��ۭ׶#˼�"�q����U�ߓʳ�٧�
*�6�,*���&	���m��$"ɼ������=}���M�6kC�J�3Uu�.��j&��S�k�YE�e�f2�J� �
0!����C(��
���u�0
�1ӗV�iI}��;�����҆]�m��W@����� 	�#�5�2�@++=��B�!��a��.6
���d�G���a��)d�"�sT�	�_���o�Ks@�YgT����e��hx`:f6�������1Hxpm��-�\�4��t+]�-����i��<0:Wf�=��H]άO�<�l�6�A���#R��A����䥫�:Ͱ���T�d��b�Y���S�"it���F�j�[�|�-G�����h���Ⱦ�1������M�᳹g�����w�0�ZV�'F;��n��/�1I�Z#��Jg�I ��5�_�n���Lu�i7ĥI��R�d��؞CV7�9L��o��f*�Xr�TA�M.�R����",Brf�d��:�_��n�r��~�x��Z�����7q�q�Z ���ov��O�^+���Y�瞣̎����AOL,�$B6����[q6Ճ���CN��QY�V
�6��6�RS�> ��M��fI�iU�*����]�ʢ��	��f9]�H�k{��M����ɉa�`�b�g�w"'5w	��Q٥p{�D���#~���vJ���iR%��st�:7^;������ѐS�׬�����W��?*5��Yz�,��� �,������?2i�;jf_?!C��Q��To�����}�p�~T��P9���zj��g�f�[:�u�2���5�}�Yf�[*�x�Um`3}�����,i=�D(+5�m^�`��Ff��~��֖�Tnɨm��z�U�T~/[�=t�B��|����)�8c L��z^���B���9,�� ���v������
�7`U��e����6OM�p2Q��4�B+O��2hصrr��X4���N�Sa�{���^�?MM���v�u�U<�Uff�L�ɔΥ+����ٖ���)�G�'Q>���Mx�4�nuI&%�xy�-6.��b������m|���и��wz^�� ��*7N�d	���hq�����T�!#��p�� ��ַ�l�� ��U��_K�I�ɐ�C��!��Ij����<����/����d�����Xa�Q�=34�b�rb��}C	�������[o3j��>�@>�9�(~xԚ=������Q1�2�*���__��&�2����k����SKQ�8&*8r�7V8�`�	��+a���yo��l�E-x����*�1�����D�˄�6���B�7l9EUH74uO����>���U�r�DyO~���o���9L��ݶϧ�p@��Quu�� b/V4픞�k�f�[ZH},�s��_�����y��䚦�4��B�GQ7>�<�#Ѿlz�դy��.�`��ԅ�%^��Y_�ˉV.E��8��;������9Hu������qOQ�q۲Sx���!A�������!�7�PGA`�o��l ��Dl�+!
�M���cv@�����ޣ����s�7�)[N���s�ī9g{��#}(r���/;I�ɉBr��B4�LA���8��B�pk1'G�R���A����E�G�(DZ�z�F�:.�� �����a,��A}�9�`�RIDU��V�BS�鬙XB �hZ�@a�!+�_�'��ǰ�b�%M��l��l�}��S���W����1Q�SI���l}�hs/�o_ԱaL�����پ["��EG��ecC��Gy�L|KS^��i�v��`�:,6F�9����K���&�O�ML�O@��N�R58��������ySx
7]@S���?M���W~�l�^���L#,4��k��xO�w:����:��?5U�)�Ni�YQ�Ҳ9����-$�T�RX�t�!m�kW�4�l�?2=(���$��1`������e\CY�[�@�ş�(�`PuZ�j�C�H�h���a�~�g��f�nt�
��A���}���C�ڕt��NI_�Ӛ�;��tMi�i��t�e7���%���iS�����`4��-� �S!��1�����Z�����ǴP_<,ʞc	iA2��Z%y��L��V�ܨyZ��.o�B"�P���t]V:,)-(e��c��d��u�\d�}:x�F�u3ES���M0�0�ը���kS�3�\(ڂ��� ��̊f����ɂ#�;�i���c�?c��5P�9@�!� M�k�G���ٚP٨��
J�Y�]��G)�s�c���{�;���X�*K9|-J~��q咤:C�"a��>�R�z ���bX�"i��h���ih@	+m��V�XC�Ǳ�з�ޮ�6�*����L��z���ԀbeI��_�i/�M%���Ԣ���Z��r���\F��%��),�M!���A�E���9G���A�fm"B�a��6�����h�u�l�R��{W�>��gm\%�մ(�&A�)��/ݻ���FIꦗ�v�+�Eַa��6�r��� %�|���:y�(�m��{U_MAeg�]Gl��I�����0	妔���j�.�*���52�TAj�oþ�AofnJ���
��_�P_R�h�^J��L�o��a��4Uȩ��'~J��.����Ly�p,~�cT��\���T�g�M:8�&�ڵ!y���u�qƭ"�B@�6%A��~�"wa�������{=�g��׺0��H�~�OrW��N��1B�Z������C+f&_��9C_gF�9T�һ�9S����>�����Rf��@E��,lª7b ES�(�}��r���zw m��C��:^��5��Ίa�Rn.;�_����i�+2q�������֛�l)S[�V�`ʷ/�O�:m.���&��&1u�� W���Y�8i��@}���:>��8�3h�p�fڝ��xW����5��}�	J�Whj$8o7;��rl�J�3�Q���bWԳ0=���h�X%6��\��Ab;Uګ�"��?F�z�k;u��f���/U����zX��M>�p�4m�41�%�,clO���f��i�9C��V�v�)���'��H�?� d�bQY;�s�oPK�c!՘3ˊ=PD'(A�8�3���S��>kp��9t������/��hu�Y�y6_V8�o�;$	x�ZK)�^��O�0H���3���蠠�Ub�����Z]��H<��y�ȊH1H�ݣ*b__�?��d>֘���'�#͖�����2 ڨR^���f�i�4��;s��3^)Ub��z	ǎ��C3!���ֵx8Ṣ�xK�Vx�">v&�=c	2�f6�W�\��Z+Dw�U3��r���{KJ8���Tl�k ��)9p�َ�u_b��@�v������{��N=��a����o8v��c����R�e
�9��Gw{zj����\�|O�тՒ�k'�~~�?a(�@��no��췮�xN�`gd�2��8�ؑ�t������;��?��#��1�s�Jl_�ʛ�[�8�ݡ���=��(�6P�?&&$���8�Ԇ�&���g(|���^�\}PP:�1��t�h�%�uC�L�7�r�*�kؽ+ל�h��[�"ƨj��y����$R�js�o�Z�)�vxb!��l.�d�M2 ��d֣p�@{��
 ���b/r�qFei����פ�'��tC��������~��'����M|IL��÷�\jN��ID���Ƥ�.&ǀ|�0w��P����~4b���Q���'(`��*�b4���W	HK�}B��6I�~���RHS�g��!�(m�R�sUyQ��$I��}Cv��zz��/�lo,�/S�n?�t�� �ؔ���j���N�P��hU��l0?���q�N�t�tI��Z�q�/�8�w��XE�rkA��ݰ��e��%��p�=�.:d	W~u*����AUe��� ��?kH��`��, �Y��ڒ�>����
���^�8�����fh����p���@�!leE�E�
6�d�P���*Kv�q�_ia�x��%O����ʔ���	XLyf���=�޺:��� ��<M����U�֪������ٿP���~L�W���?���綖a;c�ڻ��?�i�&6ꐑ�'�G�j�O:�qѾX������c���lf���F|���'^��؉z�(�+
�[H��
A�QXsd��N��a���3���FA��X"�-�t��-��C!0��1��\�\�/V�v�Mw�A�g0DsHa�Č�Y�-�@qa[��;�>��9��d�1������_��3(�����f� �8Zf>���t�]~�޽�<YZ�I�R����ƦF�.�L��u�M�l\'?s��!�o�e��O��J��Դp�+��	�,7oc�����}���� ��@����<�|�C�d�i�4���'�Q�;o��ޏtෆ�~��ޑ� �P[��i�!W �Uz�y}���BZ�	�$I��+ޢ1��4J��B�	���xXh�4Щ�����#���-�������{Yk@D�H(�Vp1#�`�|/� ���Xۘj�3��Q=J��Ojt�d]H��{)gb���yɵ�;u�^�\ϕ,e��Fd�h���䩋��+e�͊VJ�-�9��N�H*���.��cӋ��n����^$4�ļ2��4��H=��yP_?qx��9�Q�U9��b�G��=���q�ڋ�u�EDr�Tn��K�X:�5
�l�hQ�\��P�����������'Y�/��*4-�f`�P'��#W��i��|JL	x�k����)@8�9�q���5�Ne�����|>��$A	�P(���6"0��NŶ1�ڤ�&�_�u]7]�����eH�8�����+�h�\���?��T*��j{=�O�j���紻����G�+�9�!Pk����Rq7�;�1w�W�XD�'ގ{T�@�<z�Y�O�!u��An>Y���8]�$|�kP��&v��\ņ�!�K� ,]���u� ���}S��U5N��1�����f���Vn�	x�ah��<�A!�Q�%/���ǥ�8W{�$�����B,-9c&!�Z%j��K��U�r[��辍�`UnO�7p�P��n4�D
��O��tNŢS�~x�C�e�Ct�Vi�q�L��)ޗ*��&���b왌�O����.M��1s�{����`>@e��d�2}x��6���gH������� ���rǱ6�2������`��j�	�h�X��6���+-�h���-,[�u��hNd�9�����6I��H�"ߵ-9���.2�X����v&�i�ة[��8��.�� ��ӫ��=r/�GT켂�g���I*���5�iR����^�pJP!��V�[g*u{b�5�4 ��v1�+]qu���A�/�}kd�GR���Y� &9����*�O�����c�EQ��0S�)�0`�<Z+3�y�m���O��u�)����f�#��o}��ؼ=�V��_2����l@t�j9wY=8S?�9
̌������{���x6�&��:�8��.�����S�0ˬ�B�Y�gB��s��#	j��cS�n��H!H��.���T�@���[Z���d,`�-YS�����LyM2�I_	nE����μSO�Wx�T���d av�;��ڍ)ZM'�Xy=��z#��������G��qW��n��^k�t�g���<���7�UHJd�h�y�9[OJ����և�[)��k��S<v-څ�_X���͇�x)&Ȃ9v\�,��+O�h��'�VS�|+I��r�F�n��ޚ�Y������7R'�&�Mo��� _�db�s{�wg�=T�X��WE�[�[�W����a�W��2��r�c���)D��ɓ��5c�:EU�h*���i��c��X�Ī�H���Q�	��������Ӧ`�SI:l�^n���X�s��Yߡ>��ia�f�G�k�O�E'W��]X�h���L*t{�9'#8C�G�������b�����a��/;[�?��� S��6����	�t�Ȧە���������bփg|��@̃�\ �-f�-E�a.K��l�.;Ɣ��>v�E(+�����C�Z���ȵ��XrÝ��W�x��;��G�Hpep*�*�������*f��3N�+c ���#f��D~�Uq�ETE��I�,tKpc�G;"�F_ i�hdn$e��B4���2`�禲
H�o6�3J�s���47�Pݒ�3���֩Q_�i��!e�RV9R���	��kH�/ڕ��a#R�WH���f��xh���gU�<�@��}��X���P�eIL�a�.�[f�����W!J� -^.��U�0e�[��=:�G�
;#��,:B��zo�h!��!ε�(����:�u>NL�5�UW� �Q���R�M�y\[h�j>�_��a�y����nU+��-�=�4�D��w�u@���T�0�����U���ڐ�'Qe%;�������6��=��|�8�l��̇yg��N��q�}g�ȉ��ԼP ޳ I;�5�>'�N�@��w�J� /F��|9w�,2����'�;+��-}�
��-�x�<��rE��K+���a�#8zI����O�4�w����;���-�l�YI�r�f^���N�<xjK�QOQY�̤P�Ld�
:� EQ<�=�3w��3�ruH��Y��������
��ITᒻר��/�9�-h�	�]{��u�Hpz����'�Ϸ�]n8/�}=Q|��AR�9ە���؞���y8��q�ކ��d)�`l0AOm��?���Rcxe���
��Ԑ�b�8O�}}� ��t��(��:�2:�!V���Z��J�p�- ��]|����v����O�2��X���0�Θ���k���XFK�`���3�S����Ǭ���\�ſamr�ay!i������w�<ń��k�q�V��\v����B�6͋��>"�"��,��_�@8��RY����RVSi���I{�Z�V��aՠ3�jh<Ȯ��ǴEp��K�0������%�ʲ���X���Л���%�÷蜐��,E��0A,���G'B� ʧ�SOڔ�;�g� ʁ�]V�2�c$��*���Ky5�� ���W�����Ӟ@�|d���hε�ѽ�f���g ���-�4_�5���C��B�k����\��J�0��E> uL|Rd��j�T/s�B|�\Q:I�<i�o�%#��DW�F�%
E��qw	>v��U��r��ME�K��4�P�z�ޏG05ܾ.�K�+Z�sw�eS�A�[�ާ\xAK��{��$�@�B�?� �=���I�j��Į���Ǩ�%�$���u���*l�dv;wI���������]|��vi�!y����2'3�%�ƥ�Wt9C�.p�h*��씥�w�F�^��s����%9��o1Vz�;�|#����\rp�-�?���n���V;Q��i��<t�i:����?��9�ˍ�Þś̅*�P`�T��>5ۋ?�q�4T��_�X�4�Q�ނi�3B�=sW����HuҘ���K��X`�ʵs�RNv����?H��IZ� �g\{������]�T�2L��#�zL�[�tf�r���ӓJ��@P��:��x~�m
��|W.��kB��;�m��s)3�#I�w�1�a�̘�yz�z�|��F�rq~�� �6�f��E�3с�mF��W��L?�g�������7xg�L�Bd����XF%�1o�y6�ה���vˠ��F���)�T��#�9$������UWa/H�6�Jc��B�U�^������`��9�#h*�7�p�J���8�Zd�[#b"s!�i8��(�L���ǲwY4k��"{�D����>�<S���C�[ǃ�q��n<0,���3�i�K2��ƞV�9|(Ɋ�%�u�̽���@����1���;����Յ�P�AND�Ǽ>��?�a]6j���s,mg�)�9��\Gִr\ƅE�,���p=��F
Z����`M�� y:�<�g��`�g�kmyn�L�ǜ^~ǈK`5��Th^o��`j�zұ�� 80S�G�7I(�.:�5g��R��i��\� ���3%˲C���9��w���s��=:�ʖg��4z.B��u@f���y�ʁt��r��b�]y�6��}|�ɦ�s�5�|~I��wB>�|��h�n��-qJ��;]�u�Ƽ�=�IVU����>�Y�7�A��͢g/=
���v~��չ7�i��z9��2~�V����ⶶ�Z��e�r��Ѡ�^��d�4�A#7x=^�Fm�,��.��3v�	����b����$�Ǆʠ���R(�oQvm0G�Vf�n �
��me-�����7l3�E�Kݣ������o��t�{�4=~�R1ܥb�i�����_�8M/*������R�̼JX�pw���}�Yu�;F�� y������L�ࣷ�ש��Z?�U��uٜM�B��}�,��~s��Н���J��hb��4�����-O��",\�u���h�띹!(��z���e�lʰ|��s�Z���^��Y��[��bw�O2|���E���C���2�3*{)����P:S�}�g��Ts���QN��gkz�$�r������;O�?�׋R|�S1�팼瞓�;,�����]���M!�5��U�J��Y
f�jOQ�j�Z7ǻ>#�N`�;�J�L�56��@�Ÿ?5'?0�=�!O1�N��W2{r�O��y;4':�%�V�G��8��;y��;�
Ĩ�K�Hi��O>��
G��������r�r��`���m|�C�L��"����0(Ĩ,K; &������ p�� wϫ�=U��D;�>��x�l$,���WF�5lO2�@=tbI<?x�tq�#d#L."�zcÌ��Լ}���	�(S��`k�	S^�3����8ئ����>ǎ�Xa�?â���ĭ�x,����xu��ܹY�_�j:����O|��ڑ����4���+LO�
0�Q�.\Й�HP�3?�F�0{e�/��F%���a�����O�g��k�d~׺�&���F�̗����Z[�l�(��P�F�V79D/�����<hk��4�1��9mL��X�/`�u�b�k\�f�xs�`Y�!w��BSW"٩��'#��ݛ(�����
����Y3��ӌJ������V��q�
���T!�=�	#�0Ҋ�W�����tw�L5�Ư�:�{�Մ�;�����}�"`Ǧ��	�?��Z��>�ƕ�~z�K:П ��c;����Ou�@�ؕ��(r�N��!aj��w[G���K����{iw46'l��S'���;�@�"^s=�w?U#�(^�b/�T�-sG�iD�x:�9��Zb)���h�$�4J�!^QغT�x���ˏ�ިw�/�R�N��8�}���2�[�D�#�Ѕ�N~'|�QT�B�w�w�=*n�u}T��}�˃��7���7���vКO��-3��aΐ�2�^J�*����Ľ��8:,��
��!�\׀��^�a{"CmfS�� +v����g���g���3�YɃ�tVv�腟n8߻�a10ߝ]xC���D�Q8����1�x�bgAC �T��p���O�t�֖ �>|9�I�>s(��K�����s��{�:VL��P�%����2�ld�D�dN�
�2�f���S�b��X+�2�1H�-�dl��'���r�-\��@kO��`��%K0�Ɋ͖���yx�Y˫e�mO=eB�����-%x0/r�]#w����S�O�qw�W��y�C�y����ՓO=���;۾؏��m�	�9���q��f쇗�V�f���U���A�p���\lm��V�Ic椽*����d����l��� ����V4'�/y'iQ.>w���u�
CIb�Bs��b"&D��)2�*��P0��������s`�Io�k�����K���VJ�}����y��W<��GD���ڳ��>�(��I�����!���\��
����֪{W����E®T��g�{�s�����U�.�:���+2>�vXM�o
w�E�� ��~���qK��V))��dt�$S�#���� @ޟ{��޽���z�1,�zzU���:�X����<�A[��ŚR���/��y�h��C{�i���� ��&:�p��������O�oҳw����z/�	Q:9��*�E�I��	�kbĠ��	�)����?�Q���P���O�?��Y%����/�t��v?i9:kr��b��&)�f���@��@>ܑײ��)��s�]'>�JQz����݄������Tt�.��(����hʉQ��]g�X-m'L�즄�k��]�D�{$"I�k��e��JE��e�i�����N���V͐T�wi�l��4f�?t!m����0�L��/���=M/��N����'�ꃳ�\j��XY
b7����wFg|�?6t�i3��+ӱtF�Y����������"���Vt��Da	g���Y$�t:1���}¬ŀy����p}�b�"��L�q�!�7�N.o���L-�i8Mnߡ-�!��)z�<Ye]r.?�5�FQ�v�{QH�fv?�'��Bw�1�:w�ч��a5���<K���R?#S�c����P�S܈}��f� ���u����r�w��_)-~�.$|�Ȕ�g;��pfJЫ����	u���B(Ӻ���M��0��=��`����I]z8Ҏ�I��b�C�,}z�) �ﾛ>�{ϣb��M�H~k7�i���FW:��F_��P���-aE�	��n�5M��~ł+�"�� �v�|0{��i^�
dŇ�߉ �7`9K=�������ܻp%bͧ�Z������?�l~�ϳ�����F}�h;A��Q�VX�`�1H��E��NY��H��n#��_l�[��ϼf�ܶ���f��}Ajb�]V/�߹�;Z(�E����e�@�*��z���.T.)LjL�rc$�v'gV���o1��^��E�+�GaEIxH<������M��SX���9�*
K�2ڰ�"nz�n[��V�aF�[Z�wl���'9��l�-�"y��>�#೵Aj�9���B�����$ut�(��I���{�2{ܴ �x��#T�n����ِ�f�a��+2�ܘ�/ S@�3�F�;�:�W_%&�`�o�e(�]���Ħ���b ?~1d �����L^��L���� 3<%��l��>�⧙j|�x�k�����S��^('Le��'� ��c�u�ٶ"�ӳ/ ��0��Ů�ٿ�B��Ɋ��1Vm3.�׳�i
��K������C���LH�Q_�c'~*�_㐅 _2�?A�kӾ�כ�64?�b�b4�~8���RF����X�7j�\L�ʴy-�QK�*ܑC�.3L�Z�&�z�;ms 7m�o�J���	"lc��L������=Ġ%���`"??cv�"倠�-�I�ݘ�(���XJW�ܘڧTSr��vX���s��E�q\O�_cp�%���$o\/n�Q\�[����Ų���d�g���.��u���9Tf�%փA�V�2-y�Q���:�n�Z�P��
�(H�e�1�o�����P;g�U��/�u�nZK��J��S9W<�ޞ�Ķc�+<m�%�|w
��U�R>a����mk+����1ZvZ�uw���uHHi^���Ŋ[������CV!|�v8S}�;����`�k&�3j7��\-��)Y�8Tg�<w�F��t�W� P�-H>�Ŏ�J��1�*���TV�j)�Q�����syVw-��)��)�t����;a���ǐ�
��f1��(	���-��S�(�y���R�S��<�R��Z.v\=|,�D�Y��&���Pń��iK_�����f҄1\��	,d���6���f��A�iY��[��D�ކ4}'�n��yt�M!�, v�V)�=e�}:Dq��mB?��������ڥ�?�W��6�Z}��M��A�����i6��e8M&�]��<��EG�_� m톰���[)���	���DKc�@Ȝz|�p�.��Z�t.5ٟja!�g�J"��~8�J�2k�PŤ�����	��7VgM��G��d� �v{<1�'���dy���.=H��T3Bd����ՠ-����Q'���8��.%��~����@%fU#g.x
��O]�G��<�4 ���[XN��S�1�L��{b�\��f�o'LC��8p����|=Ye��=M��	���Ưߵ���BY.�秄��"{��`�_5����^�&g$$AF����7ŝS�0Z�*6�fp��I����rD0V
�UJ��4�qC��⵳��Ӟ}$d<ܩ?ϖ6�]�+Uw��T���9��ձqӥ}+��.����ׁ/<bc'� Q3%�wԓx��/��&k7	�l��%�վ����D͐�KWÖ�f�����Qz9Ų�X%w}*�ذV�� \�l�1`���v�	1����ݗ#�L��b���i�s����S�+�g�m�o�'�i���=���A�(`��@qS\3�8}U��t���a�* �0��tJ5�*?��S��+�sq��Y/���4���4�P�y�3�#�nfY��*\�ȧ8������F�������-�6Y���I�V?f����R��ǧt�o��^�+k��ϞHجT�4[��iM���J6���أ�*u�-=t��|>��a�t?P}+}b`�Q���kpa �����um�sd亢}�Ej{��� ����?������O���'؂�&��9)a��	(��
֓� 3kG�.ϛ�����ߩ����ҙ."~r�&MUB�P�	S�S,0Kp�%@$Dd�=2=��#eJ�t�F4�q�5�u�"/~�����yt%�����-����xQ�ȱu�B�$�a�p����I��į�+~�k��K◻A�J��<���c/d S�ɔU���N�Y�q����Qm7�w[��B��p��4�� "J�=f�U�8�yQXAJE��i�)��IS�:SI'Z���abT�j �J�kK�},;���kw(6�2�t���z$\�5+�����텮����$�x���3�����>�{�h'p��)<a��b^�AV�P)�hg?'�L��B��n1����O3κ�3�݄�J��ar�q���_�$"=���[��=�mm�+u�P#���tM� Ĺ&cV�A^vHҽ�7;|1�f��}޿���w��s�<0j���Bc��Z���>��e&���Bu#��౲������. {Z]�ѳ�~xuT�'�|�y�M���HF�/!���u�N=�����l����q.|o�<��E��ୈ�rB�� 5��Fr�62��i|��TD%91�,��I{zP�w��eڞ����3�ƶc5M��GfQף�o��v��Q�6�nb���ၿ�o-L�m��?Cpa���rhF�sx��b�x�ef�`�d
:�<�n
��Y'��=��#��l���[�xχ��h�z�K9�*�U�*����I����Z�?˫Q�Iĳ4x|X��_����b��f�Q�NeE�l��&�\���L��G+)V|NhF�R.Y(��$�N\�Mo�x�̙��ClE�A<�� � 9l$�q�d	��|�@�������g�B�:"��a`�Ѳ�u�oX)x��\�n$���(^���O��2�e�>�����]epH�4X����ώ��Rsx1�m�"b�E�gr͟&耎�W�rM��:a}�*��8��5�X�G9��*��ڸy��RW��,L�^<+��p
���kR�h2Ҍ^�	�ܜO�	.�$�ᛐ����4xS{qU��a�[l�xz��*�].�]���-#6������P�½�-�R����ɻG�b�@���5Lg�7�g������5U��Ȃ��/��`�{e����{������ћGq� ���`6aR��P'��<?
5dW��j��C��8P[6�����~/�%�8p�$3{�w��p0&��X��QaE���r������r�40��P^,Fٚ��_��Tz ^d��X�V�M`�3a_�^�$V�H��o?�XZS��$( HЍ���Z��'���k�$.���i;�����x�iF�Ꭰ�d>h� ��?��v�1�udH~��"���dO(]R�#î"FѰozt�.2��\Q[�wg\����u���M��NN���#ԩv7؛;C�����&��p�� Ľ��^�ʧ�tDc�~����#h�K�һ���Q-˺�jY����f.yc�pj72}����Ed��O�)raU0P��(l�?�f|鮭��|�,?� 40m�1�t��x��i���Җ9�����ś��rXl���vciR'����&�ǹ��<O��l�[��=iZ��ؓM�XQ���L���ۑ_�xk:s�|�k�R�o���`	i����&�\r��T;���1}��p�n(��]�ao�|�h'w�h�S�.��H�"1F�v7���8��	ֽᖲ�E~u�֪
�`��tE��G�0�t"|�#^@�὚H�ܣP�mK�w�&�v5�^����� ��R��r+[�32Gk4Ǜ|~���s�`�j�� ��()��P<q7)n���6]e�zYY�r@��*j�����k/ܲ]�c��<gC/�V?�Վ4������M)�AC�TX~��I�w��A�%E�����.���ov}�!���V��6���?�<گ���=u�Oa�����[y:�6�Qٛ~p�`��g�w�0o�%�ܼ���l��%m1K��p���M���f�����e7���|��x������oF׈�����rBjxr����5��[� G��u�%Y�u$�"��ѿG%7g�g�;ȴ�w7\�S#`	���<2����ڈD���[�ÔMzQ�K�A�l2���)�����>W;PP%�Q��E
`	�{�?��iI�fV�H �:qXm����>s��iIIuZڸ��,`�=��%>t�4��`�@����(x}4r��7���T�<�n69?�v-B�>�]��S4��ӵ��z��93�� �'��C�����Ȍ��<�/_8�����@��62��Le�Df�N�I��ʎ��H6�,��4���A�m��H���:�rYڋSNw7���ˍG��-��N�0d�<���z�f�y�I�����!���<��XS�!��H�_���/�V��<t�_��վW��ݻ��B����l�֑'T7nȿ�s�N�d���f�[q呝E�=&��~�T�8bz��z���b���m=�l^R#p�����!�J�#얔�M�
���1��s�|�U2gX �Z��zm!y����@�N�p�O��pB�_U�q�f�:�|�C��"��djw��
 �:��&�+����I�T���N�d��N z�+�M�@����%��`]f }�������8�va�+˹sz�@�u ��gɴ#�Qk�Cy��^1��IEPǪ����yM��q�i�7}44���r�����;��h#P_�*b����H��cӥҷ,(�T�볓�o�W�p����I�h�bD�`~e�h�׵����!L4+���f�����;b_۞?���;�C�47�ΩF�\�p�M7lt>N����z�7]��mR]X%���_�hG'��ݱY��&�Q�4�HTU[���ރ�t�x���;o9=��_X��%�P����I�SkJ�)����[j�+;>�.��5_���ސe��DH����bL����P[*��+Fjk �%P�JC�/0��~�EIyi��j�Yt���S�;�k#%5m���tʮ�'��bz=lօ�n7��K^�
N�k�� O_i�2�u�CY҃�_�t?�|��I3T�����ׄ��po�yE�i��<��^��������o������{6J���/d(����2!RKr���!��2H��U�,E�E��^�?�O[�<@̢g�Da3 y�ʖ�a6�F��&�ʗ_J�+��-�Il/C��oM�~*�B������ T�L���
���QGe�3`C����	Q��B��E�t���3�Bתhr$���=_K?�l�3T1��|�-?n�|y��<�:c�~�ep�����ؙ�\V�@Y��y���L�S?z�������&���i,������i4���X8�52��q��m�j�K�01���)���Y[6ϤbP�y���7��D4�7"��D�Fl���hާ��J�
K�ę�S\��1g�����R�>ۋ!y�%c��b���[s�=3���泰Sa�/�Ƶ�z%������9���1FިL���q/���i�Ā�q&�[?��6d'r�{D����.
 ��&"_q�ɯ�|l������ <�)�)8�����u���������	�Tk��Q]|f,�,X ���~��r���o*��G{.I�/M)z<�Lۧٕԯ6[B޲<����qaՅRCz-�������8�H۞q��%��MgufT�-h�#J�VUYI	��2@K���� @��N�{�	��9J�[���D�5��B�?�R�m'�kpᲠ2@I������c���F��+�?N�J�v��b���.SF���1�8S���Y�A��w����]��_�C�}���T�a�
��"�F˱�\h>�!�Z�Հ>S�a �Έ�?C��Q�f_��D��ًiw��A��gޝ��ݫuSOqB�Ƀ�~0���0���INp�� /h�f���;�Ҹ@���%3���Ӷ7���4��K,\^n�,+�Gdm���gxѰ�}^�q�ֺܺ/���\�P�2�8֍����m����'b�M�1�5OO�fF�N�3֔Ϫc��{R��98�X�K�K�bz��Z��O�9sy�ݳi���ƏǬ<D/d����!+�H�S���W�u�m��TJH�����ٟ��T'�}l�nl�x��wg7��6�}K���������&�A��}����O��j�0X���iT�3���p�`���`)����b%�k�}�D����}[�X2K����)��6��^��?��"`�:�:��[�r�I�N�ӗ���}˹���I2��o���"SJi]c��0�i�tLj��삠����U�����_=�k�i��/��V�[�LmϜ�ez�-�P:����i��F��%�����<^@s�<����~Ta7����Q�F�s� ����4��)�<��tpi����v�Ȝ����N&CG�|_	�,�:���鍾<]�e 2��g�7�A��_"#OZ�g�=�\M{x���8S�7��ƓF���H�-jpU&�µ ��;xvJ�F�����Sq'�7�����/M̴OI@��p�JE����8�Qj�Up]!����D9�Ϣ�[��
/��s3@ ~Y<����2�(>Mi�5Ez̛%DS���5uʇ�D�؁߹���GkVn�T��Ǉ_4�}�`�? l��D�.4�L�r����	��cR�-�����K�&Z��^�RPA���n<�@#>,ݬ���j��ኔ�iҘ/u�bM�S��8t.�0�Uv�d���2~�&�x�ހ�>wӺV%0�&osr�W`�3iev�U�E �M��	+���t�b���ˀ�D�-�IK[�E1���Z��F����CK��w �G�0�ȍ�e�S�`ޟH�@�H� =-�B-V&��GB*�s��)X �f�L� {�������'iK��zZZ�hS~�<8�yo��-h��C#`������lh5a�C1c�Յ
Bz7;��x�!n�o��>�!B �1��GF�'�kQ���/����zT��	0?��s��p_?]����j����N6лI/>�M
�����|t��Od&sd sYzdy�!gm��7	+/q��n�����5��( ��>���#l�[qI�w�|�@��
�8bA����|��}�a���ȴ'�R���PtD�����$s,��?�0
{�&_5�����d)ɺWcҟ�㌕���ך����2�E��l@�4Pl�<�綟���8�������~֝�8S�^|W��m?P��d�|��&F�
�y�?�m��H�|�=��c��ԡ/��[��~��;��:rU�p�Ȁ�]�$�+�w�j��˸D�9�?� ��ϴ{��P����\z}�|�P��F�D��P6�����S4�i�=���Shfޢ�/�6�I*��YN+ �9��"�����?�6q��ە�S#�Ғ�^L�X���7�(�2�[C�I�C�S���s|Vq��N>_}Fm�K�{���B�Ҍ{��j��e�����)z���26*2������8ǨZ6��G��n�N�IJ�Ƹ����(zSB�i.��+��e��uQ���C�w����Y�1��0�؆X��H �6�FY57�e-W9�gݒ�І�h��G�	ڹ����eIs�-�i b8�+���%O�>8V+�`�B\�gF~��o-���J�I9P��M��if�w��et-�D�`!"�b�V�S��=�c��ϗ�{��/lKk�\�}#�ɻ��0{���p!�� v��E�������l����@ʲq�&u��s�Y���#�{p��C�\Hf�/����i��lyq������u�w~D�nϴU���Y͒�mу�� ����)�tҎ������2igE\��.�*|�k=���4`
y��d���6qD���*S�K�q�N�^69���?
:�����$ܻX��_� �� L"�)/��@ �b��,������c���)e�g��X�u�g�6����r�����2��M5����&�N���Y����Cx�f�B5Rn�v�wnnMamWY��GA�s�09QY�!�|�KX��kOo�{-֌����b�9�D�����=Y�p�DH�O7�kuɀ>)����k� ���� �Q �&]#��gQ��ICzx�+˳�?�{-9X�)���Œ)�H]i�('y�@Yb��U���ދ���B9V�p៭ �	7j�G�jm/�ûҬq��A|�|ص@A=BK�%�œR�TanN�߫����%�E������I��u�Q�UK
�]�%LO�^BC����z�;�����e�f[20��#���K�� �Ms���41CtԐv1�u$��.t�؆�<[�6'xr�G�1�S�.^�h�`����S1�D&�� � <�XP��&��q�ø�$�zRُC�=�w�����9:�r��Z�C�šD�B~�����
b��ɚ�j��&�m�@��C�z�ɼ����x;@*?�}Z�dZ��p���>0=��Q�=�|����Wi45�xP��|�SJ$xj��s5j��:�qD�`$e�����0�V�N:,�	�)|3��Q~5w��Z��9�n�<YE����� Ў�n+���wT�jQ)iۑ�O���$l�-��\�c���gD��'��%c����`���(�>\��݌�F+W�gu�$�N2�2��v�7��m����W��r�Xz�NR
I�W���78?PG�&����/�	[�(�f� ]rT;;�Kd�u������z���O�]�]uE�e�ab4��H�e�����ŷY����O�1q��͒����~!������ޭ_��$OMO�?�{H�F�G_��i��Ik���;.��Ȁ3�Q�5E�h��8��rG��<��VϩRt;'|wUh�7��y�=��Mg��-�++��ט}��F���;ا��<h�^�H@����ӐG�Af������3�:Y����u�Ӌ�L���C;�p���ҫ��)���
t���0ת,��(6��;z��$6��.R-~4��[+���p�Z��|��zn�|���Y�h>���ۃ�I����8�,��̅1)�-6v��b���V�\��_f�+�ۯ`�uaK���ln��R{�3��y_ả�Fq �������`��Me ��%��|�֐6��r��ā��k�ŭ��PML��m⟮׊/m�ԅ	��O��B�
"5���g%'0a�b��hel',K��SB�����q��Ջ�Gz�
�3ߨ�j:4(É£�U��Գf?c���*E`��ۙ&�=t1B{ǡ Q�o�\J��H2����Ϧ�������'OTq[�ɬؙ����sZ�m�Nʻ����uV�mh�����ޭ;8=��&�� P���O����0�<،�t@��h.���yz٪+�F\����w����y���VEj5nga̴B�S~�m��H�"P��ʵ��5���C��
�m�"��������ɈM�'��~��[vD��T�s~�@���x_�}Σ��忊�'�����(�l�ˢ5՜�"țG怓M�M)Z�1�_~hPG� �·ԉ��ɬ�%!��H�j�һ,�g��g�4��S�9 ��bQ��8v��9`��#�n(��L��Rz�ta�{�q��&A).�M�E.g�N�r�]���짝�x�ӟ.����P�{�����3����C�Z�$��Zd�2#��r�&qK�)%�<7�`��U����q�3H�m�
j���P�o��AЗ� �-?�.�t)�R��rr��͝��et���`���R��8���	��R��o��� M��6"T���Ar�{I�T@�h�S���@����O�� ��ma�L:}ԫQɞ��=��(�9����8���6L�y�b�1$G�lF�B=�eC�+FyhRv��>�b(>`�׍�*��pZ_��� s�bg#��@��~5:�K�P���А=��R�%"�(����i
�z8���ŻC$Kq��������Cg�����̉/�����_��RC�"x䕗x	o{	X��k4�>�%�X)wx=�7sn��86%]��iխ^8�`�b�y��G�9�1�։l��˺�F����E�ئ���9�%tX龃���hQO�o���H��xBC��gI�Z�-�~:z݈�d6���!��,�~)k]Q�* jH$�����J�5��[�鄾ӽ5W:D�5��;�T~��ZZq w�.���@`�����^l��<4_��bD�A	���n_���*�$Q5QH���KX�j��1�����rj/�\��W��9�e��E����c�*:8��`�Ѯ�	����tf��+$G�_ZG�����^+��R\����FG�"w���9N�g-л�Q�ݔ[����8��*l����֠{�@�怗��W��GT�)G"'E�(Z�~@m7Z4�Y1Uc�6F���6�qՆ�n�\���s3^|lCq��u�-�K+r�p��Ç�l�vQxQ��9��3J��HqK��E&�z�ZRC����j�ْ���g��u���E��i8�*�5����H����W*p ��]'i]=N���h�
���BTU�&�)�h�Ցr<�"Nl�H�pG����J���D5�L��n���N�a�?�L,���LpFo��@�K�����ё	��#�
�^����au����d��XA!�	~���<��T�P�J����"����"�DV	ׂ	m�A�~<�h�&^;�a�g	
�G3d$��6d�;��be����\��|7r��W�Y��]�Cwڛ����PD��:]��cL���d�	�p���3o�,�uv��;5�M�T�:���~Rz��v��:��h�յ��p�[�^ۋ�e�i4��JBU2'����g�	"_Æy�t��V/���c`!6�$i nE1�'r=�~<עk K2��dWY�n��1��)�^_������]��[-j'�������{C/�ugQ O'�����j�	� g�G�o\�/��!�j�̊4�w����7O��
#[a7�&�,xtT[�_�L����$)p����h@���V�7HB]fUs�,�Y���"�v�s 㵉-;��aN����[��,]��1>�g��.ꝲcݷ�g����V6��j{�{@����j�"�x��L��L��h��J��`9�/�D�g�b�`es1N�+�u|�W��3��>^wx�R�3��y.���.��dUN%��U�57<�,�u�>弩T!;Z�=3$�9��͒��8�*ͺ�A^|��������L�a2?�� ���2�޹�!�SCW���&	- ��	M��L"^�M�Gθ�̷�DDVC���M_/*�s����"�{{R��Lee�`���b��I���M�P��Өa��>����O2��O	�|�?c�
��A����!pg[^�V�s�Q�����%5��l�e�����]E����E���y��Qb@��~�y*�p�_�@�`9G$���~U/`&)���^���u� ;Q[#����}�J���F���LE#j��,G5q�O&�3a.q���x��hI/߸�!�%-<#��W�J@�C��Zz�p���i��,��Lh��M����F����Q!N�D-��_����d҆��J��B��@,�-$� *��h3�¨C�&�2߀$n��]4a�o\ش�>��[9��z�@���H��z� �Q�<^�h~��K<�E�n���?���l{6�fP��w{����;L�m�,\�V�a�g���cҎW�nⲒ\���8����A���c�G�-��*p��I���tr�q���ϽC�HUq*��Ì2�G�$_t�c�J���ӏQ��8���ڸ�g*��2cFB,=_ZU����[�>��5S�E{ӛ���dUKp���fe��4/ �B"T"��8*󮽝�U�Q�M��i_=04���t�Y��(=׼`��cn��y��wuYp��Q�2Y���a��v,YeČ_�cO�K�#�ޔT*��}?y4��$E:|9 !H;Y�.��J�Pqs�7�����Mԯ�tZn��-�-�Ӥ��f��k�~��ٲ�d������C��wZ��U��U\[�$�?А���8�˃�|2UЯj7%ȵG���@�)v�������� 0f����5ݟ�Mv��/4)/7ka#O)��?��-��V&���>��*r[v���;����L�'6�������W�v��gp��=ҡ?�}e����GD�r�i�7�`�/8�����5�h``��1�T�ߦol��֙�i%k�h\�x�"��K�=��%M4���>�~i��������z��¾o��E.4��݀f���`����s�ܐ �I���O�
�Y[uW�N�|�7�x4���x�I6*|�U��!�W��jCۿH����&gnp��o�D:7ƼGT�]ǀ$��g��$��؏��P�U��Fy�I�w9~-��#�ְ3�%^ֈ�ip�	�~�7����w�E�R�_2p��<`	�P����0��D�M������#e+�D
��L|�ct����?���g~�U|�ʖd�J��̞j��8ćt���)�:���F�O�����w� ��~�v�܂��k�c�$p�u��V�f4+���7EC�_ L���l������>�d���c��D�ϝh�к��8���ur-��L!7+��q�����nb�k��{�L�i�ɽ�n��3L}�V�	 �o��}��j�[�Н�e�B��F�iJZw���#-���BԌKc�����+�W^�C���}o��[�L���#�	�~�]u}Xh���h5�������~;2H�8:�4I-=�" '�ƻz�#��E%U��N8s�M�Vq��5��M���v�z�WX�̂��$��h2������]����2%_�N��q�Aa�K���Eb�e�fr�Mvu�F�(�N=�)p�k�"O�%B�u�,�D�qɃ��]�#Œ��{a+����T�%���wU9�<\�����5M���+ز�P\Ǩt��-l�h��r7)�d8*�2^�i��0��UWL$k��-8>�*H_0���D#��@󳫌��H'2$��2�b�8�jƯ6��N�oL��լ��xI��8H@V��B:����G�[:���ƾ�Sl�����'�G"�nj�Kh�#GJ>����l`�+>Ǟ�B@����2�m�'���iEG��A�Hu��ƻ�?�]�Ŵg���o�-w�[�+yva��d�1vj��Y�V��)s,N4��j���F�;I��p�<���t��X�׮?��;���E��W�b�Z1���iy#|+DCC%Wug�Z��5��39��EF�T��/��ZY�զ,嫪OB�#D�̢�5!=N��V�(m'ǵG����!��Ͱ�!�#�2�R�Rjh�$(D-WWGF�N+�M.%�����"{?ع�����ſ3�6v*�� @�X�� U�#?��o�Fv��gV��~���Ҙr��"�?^�>���*n�}�!�	��H�İ�b�U��A}$����sz{�F��Mx�tߑ�,��;�� CХ83h��`c��n�ͬQ;�=���q����6�kv\hmPj��%��S������5�!e�,�u�/78���4c����!��PM���y�
M]DkЂ�W�-��,�Z��I���ɘ�����Nd���m�-�d;9�L^
Uö�8�VY�t}j]U�e;�ڒ������]D5�@j�?�Er���- ��v���E`�@"Cn��G~��J�XK=3�]Mf�3��OET����ꢊ�jm7%R�1�i�Ónz2-��m�F朆��?��D��םVi�2\�k=��kvIu��ճ_x�|.�W��A��llv��O�r���0��
	)3T�j���AKg1��ņ[	��6�Q�H�����UMlB���5�7�8t��R���{K��R���ay�?�]���� 	3ŌQ�r^�Y���n�
L�8��|�W%B9��8�IȀ����b�U��&EW/����}oYAL:8�����5&�L