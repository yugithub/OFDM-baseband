��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6O���b�;��nͦ��2k;�O�n�@�m�r�<[�UZ��Q�Qz���96�$�����J�L?��;��iܺD�Wg���Q+FVU�2<2"JA��JQ����h����b�B0y3j�2i���l{�4w�2t�3Q	<���z!	!:��-a�dB_���ȿ�"R �̛X�uf5�U�d'���8��y���;� 8������ͽ�xl��lO�zlt<G~*ްJ�x��c&:��O��#ŝYv+����?�D
��8 u\|�E)����E��E_� �?�i7���SG	�=�d4U����4���<#P�o�5�Ng2X��X�
�/����Lh�$�ۮq�!����
{�{O�Le	rZ+7R�����ⵣ��|:K�Ȱu<i���n#���ڄ�~���j��DX�����-,��@���ޞ{R1�Xv��Ώ(]}�U�,�b��܋��֛�C�I��u)*R~����qE�"�x������Z�we�&���?J����o�c�6��m��U ׆k�WLi�O_F��Tؾ�)\�����Ϋ�\����V��zS��K�71��w�L{��UӾRj���cm]*d�t�N)Ӫ@�����f��?C?�A�b>Z{��>o�q��jV1'���|�a�\_��Y�d��`�&��3��k3B���+��z�S���w�U���}��i�w!��s���}�V�fn+8[�c��u���!t�L�X*�}_����ZH�9����H�4�}�{
^��h=/4���mFz�Y�s�}5L��si�:4%{{��6�|�f�{$��mn%�+�uR��;���M;�+ %�~� 0 ۡ�v`�- z+�s+�P�Fhj*K!XA���-BǞ{�-S�)eYv�7���]R�&��mv*v)q���7Ras`9f?��w�_����(�wq���XVPx��@�Vg����w�  ����0�
UB���^�z��y�/8��ԌC�㧖q��w���Kז4:"$��T�z�[>gc����$F�y�O�-ε1+6XkQ��~�#<h �J^�M��1��NgN��K�}��3j̔�{t�}Fy��H��s*|D^: [w�M!��F	�V�o�x�v i );]��\��'c+J����@��ֈ���n�����+��Ľs�Nn>�|�b;��Yi+�S~Ť�	��Q-F�}���R����-߆	��H�A�l���������q
������5~Z*ba.�X��Ny\����im;s�pb��#��~C#��X7V F~�I�
����K�GB���1��=���7b�C[]�=Yz�Ę���9'�ў��BO�1/M@��R�5�T��@���J�3� MƊ�#�`:�⫫[��d�β��w �l��7Fkl,�esW��y����zƮt��dٛ�~�u�5Q����n�?`mI�t.B
l����d�L���6���ƴ��ՔK��^طi����:.Qc��նc��]h� �l?��8WmB��	⺗c��'J�/[�E�^��.��澞䜛s���KF�F�&��J�"��?�E�5e!8*��B뫆_���t�g4���<?���N�;T�/��q;=%��{r8 kJ��[p%(&��X��>cmQP����M��������h^Ղ�,�i����5�<�����JoyO�9/�`k܄�7#�g	ȫ[���?���C��*�W�[�ɨ�����*��6l�F^ h^�ͭ���;��w�N[��H~�[�p7�Q��;�"z77&Y���$E�bD#���ND�Yq84�,�]k(�.��(���P��v]]^~E7ο���r��`�3!�i��	Fm�W)
j��Za�yc�ߏ�/�a���CB�nٲ����%�d`�*!S��t&ߺ���x�H`��4C6�-L��>�������Cv�:D��v!�h=G�e#���mU���SsA��޽v�}��(�R�mM� J 1.����Ka��I��
�R�N�v��x�����Wm�.�^�y ���g		�t�r���,eHB���ʋ$h�M<P�M���Ub��΅A�p�E_���g������_s�O�6ĕ��c�����j��=r�/���]��@�Ӑ�ﳎ������i^���S�ghZ��QN#�.��!.Ę9yc�0C;�W�-�~N6	���0@&b�9�A�ڼ(Ԛ�C%�M���m���cg�<�V�1�8V
�Mٱݠf_��0a�~p~th2ޙ����m�?�8_&�^u�r�<ol��'��+� 4�V�Bo��@b6��q�L]^��񽝎Zd�"#-o�x�����ޖ����Ԕv�h-����=�YX\2���U��
ٌ��1�Q2��c�}^��<�K?[݃��@l�㲾�tԷ�L�D�$Llw�Pox-�\���t�G`��?���3,|r񣼆f
bΰ(Md���>�l
�&�����	�G0"�.pQ�NO<���6�gMq̬\ �}���hE=��(�7���
����<�vC�@+X�T_���z9���]�& ��5��]6x)���*����n�}F�&��n'�衎�g�Qpc����٪���N�ck>ܟ�=!"u��!��{XҞ憔Sʰq��;�������f��������!R�Xx6�S��g%�=)���X}���I�� \I��ڻ��}���CE[����(�gZ/��H�gZ!�
��ՒUYK��< ��~f�U�I�����.�>[;蒁@\�gB+:��] �nA�D��_DE��>��I�?I[�]��z�x�)*1�]��0�Ҷ㟔�3ѣ��_Ѻj�L�D7�nd�0/?d�N��,ZȣNU|��!��O
T���M����c`[�s�/�{3�M��|�X�?�Pi�eP	{A�ޚb�g����Q-��p�^Q��i���+2��IY��rf����k��?�i�������B2��r��0Ї�K��Z����i�xc��	�-�� �'����m��^�"#g*��+i�s�~��hds�Y��O������5���D	Tc���|M��?�B.qL5Ƒ�����|��>}2���0���MufF��Nݶ�#vtd��� �ƨ�\���2�m�b9��}�d�y~���5i<�x%l�fI߷�t�MV����&����,�(�� 7a �.ђ��q[ō���ĩ�k��6�N���J���M�V2�w<n���i���D)#�9��5�X�٥!NM��T�@�)�pŮ�w]�͂�R����	^���zw�c��:N7����*��{6/@<rJ<����g`"��mܓ��];���G�	/�ـ�ba�G$���#'T��w���,r�T$�a��@���~�]���ƨ=�O��;���\���VY�C_T���C1�:ĸ���#��ZX��gC/R��X[H����X\��sZ@� �����|�K�fK{A��蛃Q���6q�O�|S�ۨQ��� [���c��?T���6���s}��A�"�i%Ya�n�o�M�1\�I�����~�P���Z�Nd'��R6�i���JN�#�#��8^��q���:�=푎���5��Fɘ~��̫���j�*EoA�pQ��"�9#��X��<��0�k���ґ]��.5�K��h�:4
j��lxTྰF��? �p
ƈ��ꑤ�|��ȱ��,*v���/>ĆZ�#`w�񶡳T�BG�]�i�ug����Ëgs�&;U�lp�AHTǮW�(���G�">���{�t�����7ҠH��똭����.x�c�bMg���[�55h2p�>K|��j9_Z�@��U'MĉX�V
��C,>ų�A!f�pr!pzG3�����Q	��K�Q����ٕFP'
zw%X�]��d��8]��N�c�y�\�=z��\�o�t�+�84q|puY@z�?dk.�;��anU�+Mܬ��)��FD6[�h�],��2�SɝQd%Eq������a���m��6�;%�Qs(�Q���,�߈��-NY����^��[Ml��V���4]5��u��\�Apdċ�̾H�?�u~�&�x�t$W���-�i,a���"Q�ghL��g�/H"��c��/��n�:��S�Jp�V鞬�J��Y��^?"Y�RR����i^��TZ��<�B��*]�v��ޑ!�{9�H]���,0F��8F�B�ʲVx!�k��[b�M�	����D�Py��4I�e�2�m���)Ga���m`������۱@~%jȂ��@g���
����A�]1 ��	Q��Eݡ��W'�� ��B*��F�N�8F�a���n��|���K�@�ko�b�Aয�B35�/�����eȥ��P��ޜ���˝�s�P�&�u�I���;����b׭�5 �G�rv;�+�h	%%�ۊI5<���;Ο�4^��Z��U����Ǉ/�����d<@5��&v�2L��U���I$�xdtZ��+M��ͅ��8Qi�+Z?��?�q����������AC���0�je2��+Ʃ�m}���ȵ�Q�Lc���	"3Ӷ\�����"�MV�KY^���ʐ<7���G�S��ʉ�m���]�gNP�*�/zԓ��s��V�]�Q��r�dn &ߨcn�c9}�B��O�q��L<��J5��[Ӵ,��s��Q��Y&,պe��oʲ�2����v�6�+�X��af��HE_D~��ͯo�������S�SӺ��J�H��05/B�����!Z�a�ں~�5��p��_M?�_6���>%��u����w��Ju��Cn9XY2@{�2��*:�Zw�Q�a�͎��0��l�<ڢK���
;������.�j,���3�� +0��
�e���Y�h���A�$�|�B��5*��t�����E�?����4��|?.�4'���@��-�
�����p2�?�D��S3`S�l��}t����wj[[�rk���\�]q�fn�V����%��I�:���T���|��7��G��rUH��keK1?��Gw�k�zU�m�1���r r�y�SK�����.���<����zހ9ͱS���)0r�O9yPڐ�o�BnL��s�ȋ��3>��a� ]YsOS�itW���%!8��3_��4QysA-u�5��}-���_@7:<�:/e{7;\�9��F5a����A��n�X>\ꋘ�	��QI�3OƉs��2������P�`c�8����S��)�h*f��*N5� 
ݽ���U��{��]Q��� ��N�0��3��m�7��wm��s�i�^� ����.ΐ���;z���	?�n:�c?j�M-�v>�sP[9Q�衟Za�H2��u�x@k8�ţ(M'���YR��i{�m٦ڻ-�J��{�X��R��4�����wŎ<s�
�^��xlIY����i}�yQZ��dYf�Į�:QoqPǪ0�"���H���̗��sW[�ى��I�fH����qT���3�b���B�@��[uE����w����]zl>S��Y�K2PJ�l÷�&a�i��#;��qC��
����D������$��_�6A��c�O[��sH�	�	�~?�C�"X��}�W�]3���-f8?���i?�������21���&��x͡��H��\/|��5��vX��=���6#V\�o+r$r�܉�CG)��6����P�B��?�Kp#f��s�t:���Gg����90Y2�Z�D�.���^ERę��#�җ�*+g.c����c�
� +�N��a�y���1'�F��a:�P��������B+�(���L��t����������	# �%Q
2�����g��i�r�7K�c9y%{lv�{_�)�;���B�\l�������͋��IJ���Q'@�x����&�Η[�E��'9!��f�~����A6RO�ޭY�@���PÀ�L�X�R ���ś��0S4�1�SX�&?֎�CĴh��E ̴��rN�M�:��~���1@IRϞ* � ��$���w�Bq�y~�tQ��5<��Ea��[+�Eh���Z� �FA��A��TN��1t���d^K6�&�w�����J����^�i=π��q���J���Md�n��[��_�.
�+š��'�jr4jj�D*�Im���&�ӭ�ͩ�v=��Ƃ�dh�ِovI�"FOq�WcDr@����[r���8�	�%F�SL�� �w��x������?��g���F
���L����p��S`Kr��\K��GE��7�7Ң7Lw-ϼ��7�RrwFP���Q�@a%���~+��G���!Z*���(U��U
6��l�����h2]s�K�V�9��=�s����Y���?��:�� ����rGd(��b�ʋ�pr�ϯ���J0^ 0�)�C�摊��K�4O��?o��,�̍��	�l�s��Dw(�2܋~5���7���w�3녹��:;��i���ca9��u���\��Y`�����	�+~f�����kzvU*�Z��D����!c�H�
�`�m5��-���9:�8��Ou~UR�E�A��e�)�G�c�A�ww,�`���;�տ͎Ax��5V6'���KSV�Wp�"e�˕։��gw�����ls�Ř��*��S��Y0�/��)�}���@�@ug�H'K6�
s�\G;d:RgKt5����NBy���s�X�,�r�Do��<��J�0ݾiM9��|�gsӢ�! 8q�$��Q=����Z��_���F��T��b��>x�gy�]��\a?]�ͮ*p�<�;�W���Ơ�cZi{s�����1��� 3���*����[�L�vN�D&G�Vc&���æ����^���l�,.�����3�!��,��+y�q��j�L�Ѧ��(��;�U4΀�#�%��>�'�b .^�|�Ϭ��k��B]C�� ��[��(���9[������0y������9�q�h�4V[]���˹e'e����އ6��.������$ Ȇ��Tua�c;�R��$�؀m�c T���3pF$�J�T�,*�Ć4�F��k�h��������(=���k���B����,L�<�?��q��i�{�Fh��SSW�]w��桺��8 �� `D�:Rb�+�2�TTj�V�F�D'?KG����B2�{3I�ko����(&B�ș�=�`���r���T�� �Ɯ��y]SkDJ�J�S���	y�woW[��D���P,Z��t$��r��!NJx@�$}��x5���4>Z˩,�	���)29��,�5�=<d�����Vw�#�o�8ϵ�XB��'x�Z�����k�k�	�;ۼ��d��Q4b���=b��B4�V$�Xum|T�v�j�3��%�>����T��_ �	H�����k1,���}�!�Hh7󉹰�����x�ou�(�͒#�t����I$���A�g޺���-���,C,4�S�����r�����������+��U�u�C;�X�+�d�6Q���V]�G���Oz�>b���r�%���㾢�R*LB������2� t��Q?�te��Jv:��#������?��y� 6�sr���	�ڼ1����˅�%n:��to���Q��|6���.�u�H�����r79
F���i2Q��" �)~��
ʍț�H���s��팒����Mo$z�_W���̙A��U yӺ�F�$����$��eL�����������������G[��"hQ������/4�do����́	������<cB�v�d`
�'ax �ۦ%�`R>>�e������eFPI�;f�h0��ŞC>d�P� ��ʱ��r*(�8}��P��͟������Ð+���8�%���ɉy��8�<iKz��8�=;)Y�R�P����`�����	�`Q�i�a¹��o�t�d��}��͆�8�_�"D�3n�-�P�C�J2�z�vޔsQ�v$���o�����>6�k�	�c�o�h�G��W��#�z(�U���gR�n��� �]"�$�r9�l9�;���᭚�%�Ϝ��C���㕏�4�W�RY�O?�k�J+d\%��'�wY_;���Q�����ĉ�U�?����K�`���kB����28�BԻ��W�ё���c���	g=���#`Wa���=��L�P�h
6F��5{Ng�&����X���9�R��D�L*�6��.�^�I�R=��H�.�>�^���፮�Yg���ڻ
�*�%�]��0+�ʶҽlu�'���������.����DOI.b6L�y�R'��.B�,�1=���)+�A�-0��e��j=`9���4��TLk$1�9�aA[�[AYxzq@颋n�4򔾅!��P 3ݮ���M�C��ق�����5E���WrX/��.�ӣ|�We�|K�L�#g�k>e�<�G q�|��^u�^�8��Ж2��#�N�u�W(�ɺ[Sp��Q��?ġЪXo��+ m����'�$�yW��(b,vuo`\�r����h;jO�%u�v��J��C٭.��h]z?#(��&��WZ�����ˆ�dq�rV �c�`+������ :�nv�Nw~ۯЁ��פ~ V�1�7?-
������g!CrQ����¦Lн�QL$�/��}�"�Ԭ�Ʒ	>���
V|ڱ7����PX6��&�pyV ���3~��u��
�Gڔ���7;�����kA��%��`��e���8ĒG5h��Z>��~�i�r���Q���^n
�'o�<�ݓt��F^�\�H.�I��6*z�mOW���0�O|Ӆ��n!�F�G3{qFS>M�ǅ��Ԛ��\*^�g��V��k���i	��'$s��$rl���,��u�_6	l��OMt]=��ԯ�W���"��I���[LX����$�����$;_A)*��3<ʇ�0R���-d����꒤E ����Ԗ1!���{��(֦�\q	A�l���b���:ĕ���,��u�P����T���X�=$Sa��4�YCdJ�)�[ǟ�t$�lf�"�B{�r��1%�TĊ��&fJƬ_%�F��������ih׀o����>�%ۊ�H�ݯ-M46S`�1-�OV�:q���׈Ή�6�E�"$Z맳�z��,��8�,�3vϐM���$�Y�5	�q�ߟ�6�ɏ [0��$����A�YG3UHO����z�� ���q�C��	�k$�o%&'X��%x���nB��ߞ���v 4M�oN��h��2� @5d��`�&Z^�u�z���@1�C��%l������f�����bZ@
G=��.�kTD���g�0�ICX��ؒ�C��G���=����TM��\���Vv����W��`����63�y)�>�m����GO���=��� J�g��v܉���<�Y�l�]Yl���\#k1�BH�a�tz<<�R}�<e�m�֢f�t<pX:���NDV��]���*C$?��ȽfR̶�4?�H������b�MbE�=�;?~�(Վ�l���H�����`�?]2���������{���++߸�v��G 2�kGRΐǘ�X閆U��s����7wWC�]ͭNHdkE�s$�Fu�q-�)���$��~� �e�<<���W����hh�6K�B�U�AC���P}b�Lw^�5
�|�02-��mڠ&Ǿ.~^o�#|�%�����*z��yJ�\����H4���5�0�����>/l�E�:صP"�$ɛ;$>@ֶBP(rB��:�U�Oh���f��Y������.�B �����v�j�̌�jn����&U%`ޭ���H%�qU�c����ڤ�K���B�(��A��n��� �
�k�E�4�����mZ�����UF �~'M�Z?�O)��j�-��.��
a ]�^��$'��bF._x��be�����;�"�̟��}�7�7� )Ã�Xc�j~4��=���`k���k%��V�k��׿f�A�|�Lu�+�I��0��h@����O
�꥙k.�]{:�y����)��e���5��!�UTɎ3�<d�Ε��G���c��6���4�+i���"����6���7����o+0�a���癩�J
�԰�s�}S�d���ئ�2Hgw=��(��yӰC߄�_TF�a��j��#Nt�����j��5RCD�����0���1��;m��W�],��" $�A�S�
���
q�!�� [V1�#�ʌ�a�Z����`%<�
)8� .J)z�?W�5@���ܣu4����I��&u�y9:�p�(H���Rw��޷��|�y���$߇Cw=	�k'����yΘ������a=?�}���X�=�k_�,��٭yI���ɳ8יִ5�^]Dx��C^�xZ��X��ݑ�fT�(�]b0$*��,Lu�X�س�!b��=����!��"]���> ��q�:���Ĵ:�VQ��Z�ک���!��!З��� ��&'�˯�/J�Y�Z �W+�L��u���/�g1�����=��|�a5nn�fPxŊ��������)��Z0�/9��[�),�C��L/�]�=|��2UZ�~l��E�����uN*�j�5t1� ���qXr���]��E����M��5�:˯K*��F�V�\*m���Y^���P<8C�)n���v����)� z\s�YIzt����J;�cz�E;�]�=ڪ
T�J��3��P�t�9����#��`�0*кIk9�R��S��Y1�%��r�[� !, ��J������w��y�aA�V'���8�Kͨt��}�YHŘ"Q�̚��l�0	O&[/�m�QUFD8\���_�������G֮�>�� n��Wg	�`J��SH7/⭪
jg��m��ca���7�u�}�]��!SO���Q� !��3$>&�k�Ӻ�<�+2B��HY�Qo�o���IݯHÆ�j�m-�Qגp\�yc��@������̗�9�u�qM�6*�-XU���2)8#�]��zKX�y���/�⡵c:Q��?*v��rm�g�[x����i7��V�$(&&},:��ճ�N$_��0[á��=H/,oE6G�c����"0^B7,���gf�2�x[_:�;�EY]C�BAJ�8�}[=�Ⱥi��z?��`����~�z��	���ǣ�DA/[�nZ5�}U�m��c�q��c�l���؍Eښ����I�f���C���ǩKg�R���	��$l����!����#���%�ekM1Q�3]e=y'խ�M͆�x�W��d�+tϚ���֕�;ŭF������V�B�Mǵ�e�v��4�O2�4�8�Ӊԅ�~d�H��6�Wr�l�c0�DE��F�"JX�Bۡ5J�Z�(=@%Q�,!�9����Y� k�5�k�����ͺUO�����c/�e�3�Lt?f:Gg:� �ƹ�-�כ��;1a�ذklb�>�S����q�g�6����ə=_���ԯe甁�����F_��񷳫�N��Y���ƅ��oOr��]�eP�4�6&��#�J���f�9�_��<�4IZ�����H�SA�YSȬS��G���h�h�-���:E$p:dě��d�Q��~�,�'�1'Ѻ|�+�㱗|�'"Q(��ޏg�o�&�#vA���V�S�SR;:�|�LC���ض
�k�a���E�B�����$Ɨ���FM��i��ā8�3�Q�uo��VJ���5��_��B���5�6��&�X �,�-Oҷ�W>C�$#�0K�z�Nv/8*-�B���nF5�.��;Ki�x�h=AB��ׇ)����?�F���U�E�����l(�1<5?�����O�M�DY"q+9�(]�ǹ�F?�D\g�`v��,�bBq��͏�o�	*��a���(��E2@��J�If�h&gD��}��Q����xR��2����{���.x��#��@F�=�n�wAF$�K�0_(��~��a�/V$�;l&'��= �>�<v��s��Gf��z_���eT�^��6�/��QtW��g��{�m�ᅜ>�o�r���j�
G��?C��%�H�t������PUz"�'<�iʝԱ�A��e^�����mʃ[�*tZ������[���t3���S�,`~�=�L=g&�6�Z������ˣB!#�"]�]�����eLj���jY��&"v��I�e�/���͵��3#��b���[�w{kb���$]Q�+�Uv��������k�5�B�]U)斌8&{��A\J$�7���'!����}���\�Q'�����%Ш�4��S�M��hO_�Tw��<�����#�a�$��VN ���&���S�>��{�x`�[��&rv^(��}���#pX�ʲ�)>���T��\24X�e��I��24�8�p��`�NR�Nv�UÈ�P����w��D�܍���a�p[E����1On:��}L\��v�>�Iq	JY��\<~-������ڦm���+M4e)6~4d���;@~�H�(���1��v�U��cv�i�T$9�?μd��І�A�5�j�$�1�=�x3�b���������1�����zl�W%���WGa�[|'�(��B� ���U��-��gŊ�`�z��b.0�,��>�8wJFf��U�I�P���ok�+ľ�)Rm�]y�bj��J2Ex����ghz�3�s�u�a��'��=��f9^�zT�����6��c��1�)�"L�8�*|��}�W+��E�7���#�1K��ۛP|�����T��Φ�<Ls�i�>m�Z�WA��-�V���u6�8H�19�1	��Q�\}7̂ LY���$�"��Pqة+L'��I)�T6f�;��������}s�p��4�<��i��sў���R:yr֔�0���+7�;/ċ�f�A� K���*�I�M��u^��3���Y�BA{yt��?D�z�"��8���>=��w9*�|��`c+?��	u�������W ��qs��~!���=X���Bw��ii��,�@��Y�v�a�hv3�������P�[ݭ[�D0��5��HyT^���{�p�U���-�ȃ�{]O(��������4�Z��4��v�ӧ8.3>��mnH�稠�{�;}aU�$�� {����H���y��/�'|I����9�y�#5�J���#nKBI��pܩ���Xc)��T�#�)���z�{��g�3�C.�&/Q`���$�� ;���T�E��{�@{'O3���K�A$j����}�Tb�	�R�}���x�Y�s���+�e�@��\U�_�#a 7��	��ގ��R6�;A�d��<_v+�Y�n�Q�� ���R�3CK���W�e�.l�p�)�$��jE�^����tK�$�6�Y�	��ܰ�ϝ�1w�`UH·=F8P�����|bԇe�z�@W��AA=f���x6>BU�<��v��B.:5S���p��Ӟn��B�C�P8X(���Yw��<���E��ٟ�H���m�Q��i0�),�nWU��%�o3,�!���N�nN�P1�T�%嘂�N��>yH2A��vR��������,�Rx]����x6�4��E5tSq�f��dE5.�o��sho�WG-��t0[�y�dF�����ڭ	��(�T�it��L{�����,��q�6�_)��b"jg}ќ+���#�e��m����͜�c��%놣�~��P�q����}i�P��V�~�D���ڱ����������*,g�������Ѫ��|�诣G�Ҹ�8t��=��0�4�����Q��T��-BF0\�{�H��<$}��b�qS�5�'¡˧�/QD�sTh�.�!��
?��������F� �|�4U��O 29�|�]M��mT�	��A�E��2x���D|�Eǖ'���%`(���|L\��F"t�l$����B�T'[�A��RD~�vt�jD��N	���v+�nP5Y��� H�4����X���������#a���p��;s�Q���8v�v�X%���q���-"�;>(�8S�+�>e�炥����B@dGk��|P+�.9�R��AB�	�߄1�Rӕ2�ypF!�R����IAi�F���n�h��E[��Iy a4=i�(f�^�a��	DA@oz.��� �6=��b;�̦���-��;"o���fž��)L��"��� Y���qv�`ӊ�����J���<�DQ�O��Ԁ�R,h: ��p���Ō�jw߾L�PL-�:wS�E��Y�w�_���zG���n��P&$�{gw�8�1��[s�á�w/��댝ut��r��ےH���L=�K9
����;�( \*�Ű�^T6Q��o��D�6զ>�s�+�r���Mӕ(�@e	�RCE\�.��[������}�_ToK:��Gwq�t��Y�~c6!N���W�7t���љ�_+�mp��S�Pu����Ə`i�I�\O=���вQ"�cߋ���|�!��_���`�H���?�j=ي�� ��1��梜���>���upb�Z�g�E�:�TԳ���[��e�k" �ُyP�Ou���c�&��3}ڌ�ޫv
���T�?�N�[6���zx���s��w<c��,�# �<���v`K�e���c�J ��`��E��$���E�0xbv�Gs�_���*)mÃM��`7�b[I1���*��167��_&v3�i���(XGb���c&g���U4�K��VR飱�H\ ��������2N�z��b�(u+���@+�.D_Y�s͂�?�@�x�5V�1�9U�$�%�=
���|���n����2QΎ1�������iɱ���N���1��bh�Uܒq>Y�:o���� T�ֺ�&�����o�D��̶��y�P�spWa?
��	��7�KI�0�Q#0�S��i�@t�y�~��DKU�{v�ꊦ����>N����K�����)y�M�S�%6[�6;Ki(�;z�Lg�|é��s��p`����6�u?��.��/r8�q1ii�P�&(p�n}+L�끈�a$(^M)TV��I���]��i�kz�+\���)��~�o"��~����=�{}���w}�xf�F��Ip��|+f�*_N-D��8���7ˤj����|�֢򄚐��3p������3tF�lï�w�/#��Û�O��~y��5W饉�����5�9�=�l��㝝QAK�m�:�8!�L�lMꚕ{�PW�&g�̭֛�g���O�����_��gi[�9�2��I���U�J���=���5��~�#md!�A���� �7���8��$x^�+���ib"p�:ne1���*����=��nu��N���s�,܃9��#�����mv�|�8��1Wh��#��74���I@��w�u���B\R�]�t=^�W��t&��>�������T ������u�[�#�D3�~�c��E9�/m�ȡ�z�vm4Pߗ�����x�;?����y̯��e7.ƭ��l�&W5�=�b�"���/�Ѻ�����p����٩L�i�Y��䳇����ge1^���I�����e���ϱ%3o��W�Y��u�7��}��C��[�Q��mB(C�^�H8���3R&Lj{�f��_Ϣ�M�V-�ѳ�Z�
j�)S�z�#;ɢ����ǌe8]�d>�-�]�O�Q����qֈpDI�
놥�@vq���6�DL��o񡪴U�r�S8�
|��#�q�Pɶ����?��&un*H�Ǌ)ԧ��c�i)77�C�Z(	��y��4�p�:�;#\*
���KSb������˳��*��̰���
�Y��3������P!׺�<E��Upw�;9�P2�
�01�T6�f%޴9y^A�y��/�����7�;oF�
���Q��5y���]�V�X���"��n	�M�׫�_\�'c���,�]���O��r>g� 4]#1����"P{����D��ư}�Pk%V��8�O3DM����`���yHvֶ��@�@kX�,)ۦW4��
7�=_ԋ.���%�q�:I��9�	��~�숻d ^ӛ��n�����u̿���
���f�Lyz�v�7$\
�]���E/:r�̼��d�!A�ӊw��?e*oǧ{�G���\�d�b<O:�Sgs_:'6�å���#^po�D탛�'�u@[CX9!��z�����%u��m4`���ExV��;;ݺ��u�w�\7���3����������i�q�2�+�13����A��"��;�1'�ȶ�%����'����^�	��vף=�eG.��}rd��[tM�g�n��!u�y��R�V���d)�{��Hm�M��vZ;�`$ع���2��\�s#�m!��O3R:lV2C���=JP���h:��/��~h^���&6F�u	��Z���T߀/~X{�&sQ� Nj���jQ6o�er����5���ȝ���9��u��D�M8r��@����!b��Rj�o�ĶS�1���̮� ������	Q��h�X�r^�A��s�h`;��A�P����:�����G��Ǣ~�&�m`�~ǥ���[�fڛ�g��M���o$Ƭ�^h���@��)�^s���}� @���=\��c�fp-K~t�:7l�|*���L���Pu��������$$��p�U'��;Ͼ�/h�0����p|c���fT�CZ"O��� n\F�eR7�cܝ��_�}�A��J������M�ob�N
�E}�+�^ژg����URՔ,7���UY/5�mf��������.�-2�`�<�'V>�R����^
]c�v����F-�ܟ2}#@�������a��d˪F ��������^�Q� ��TH��@'�cR����9_�t�%�a��/�!��Llg��D�toք�g�axOX�~��*���� �S�e�#�$���L,�xf�42�ҟ;g�{lk\�g�/s"�U�*<#h�N�	�u��m6[�升�����zDO���MS7�0�t���[��T�7o}e��1-��3�<�"2�����4�J!��J�[5��_�^rt~!զ�I^[sq\�3~u��l�{�B%�X5V�>5og��q�2�3<��t�u�,�9=	ҫ�l�<\?@!6���9~9�� G�KGj���>JW�7q�OɅ{����8֤kt؏?�7˼晾2�ˤЅ�3Ts��k]O�9	Y�O���A$t���a����Y�~%���_���105�uh$�ÛPM�ӹz�� ƾ�!P���oV��M�w'�J4JR�m̯��2�t�WTYd�a�r��qp�R�aG�H���% [�\���.W)��Y�6x�&�p�;!��?P����~��������_��(��5�����+���<�7%���"q(�P�tQܦO���A(-g�$�7��$�r���|b5�t�����Y:���K���>�������}�"Zݩ�5kEi�s��q�ֵz�1��\jR���ݢ$�<�	�����@Ju��K$,G�\�r7���Җ._�S�o���k�)C��m��~�I�`����#f�f,��w~7�kfe��X��;�?Ϲ�ǿ��H�K��o����q�U�g�.���]p}�ZI�*DIg�SI2���;�.�|�9d����� E��`�9��QK����n�����5ڦ)�O����˒��ڸ;�}���gE�[�0:/̮A@$�iM��v�~�Kݴ�!����e�0��K�@s� ��g=��ٍ�N�h�EV&HTB�w��E�uM��9���9���Pq.�Af����&��p���s��e��&�6�X�j�"QF4���Z����-i��H�����'��^����5Ƶ#��Û�;� �<�N�u�����pa�k�n�ٽ:T��N��� P�y����N�2���ӧ��h��m|��zb�f��Q�j�Oŉ?o��-c��+�"��dCSu0��H���v��ޫ�����ꑝ�����)J��h?W��P;�$-qo�F�;��a�h�_�8 <ޫ�2g/�%B
�M�rSǰ��;�6��%����M)��;V]akM�9�`�d�r�w���%�,�lyjb��p��oI����s�dB��	F�b�t.����[[,hu/xp�/�*���Q�s�aSR��f�a�5���z��p*����ڵ#�N��p��N���vL���3�V�+���?c4��}b�:�������LtMм��\��'���(�@h�1�c�z	��CR���	��rb�X�O%7�w��U�Y�ch���4|{և]�|ŏ�0g�]�7�n�B���Z�ߝ�;��N��6Ud�ع�GH΀=6��ЎPY��zl5*vP����2$׸��%������U���c�^���DE�rP�qp��a������Y��}H�¾�x���{��ŏs������E����@0�����O&�ve�S�
��l�Ъ��45o�Q{띍�+�D	C���4���Wz�[��ҳ/�j^TW n�	��2�{NCO2L�be����������8W
�?��h	��D�����;���t��,nt�/{{<�XLuz�˫vn~*�{hr>��D�~1��������8��!�<i��}A�|XwGCɬ���a�M� Q�6=O��d�VL��M�F�*�� 2�<��^K�������ub��j�_YAo����R��N��WnՐo�x���cW�&��%����m�XeA���Fk>�s�u���Wx\��:ͳ1�K��|��"Q�ǟ
l����Q�m�ΗL��ڌ�e��9��Cs��$�Q[/��-לJ��%�E�Zn?E�3�u_E�T�.���)�Y>| �]��`���<m�j&#�@�S�ݸ���X�z!v>�������60���T��a�����
�.��d	��7R�$��=��3�{E��}�>�{�	#�1T~�ٺlB���9���wc���`n�f��d�FeM��+��$����:��F\�"rЦ��.�.��o$~*@9t��&qr��k
.5y ƅn���O?+�#�ھ\j�U�C9�����ě-��{��ߑ�T�O��k�(	uh��*6�b0Y�W��v��t} wʪ��<���m*p��:E�K��7�](-�y�/�RI�#��/n���.9�X]�������O�YВZw�CX��gpn�6g!�h~"(������]o����5��>�|�\��`byՖ�����/Y':FP��]�WDՄ63FYEF�dГk�	��3
�ۻ�P�!͚=VDqx�?���;���G%MҦXc��@��&�����7��v�t����>��c��������c�r}�d�����]r��t/t"�?��#	!/��/�
���%��d�]����d�L�>b�ߐ�������[�㒀�o*Ω�R{�^�˞������D�Z	��zU����-����f)�#{��I�10߃���)�@�o]�2Ѐ��޿O��	�K���`7dn�B5��&�~ehfa��Kd�n��0q�����Պ���HW��#k�j�ԖL"Q4��
�;�#/�Fd��O�y�'Ӆ}F��@��X����@������f���#6 �Jt�i@��4�n�a�v��^��,I�y�����I}$~T6kx���Kᑛb�~C��QiU����U���� K�yqW��=�(M�s����KG�/��ڣ��G��!�Q�6@#�ʃ�Q,�1�
�9�p��i�[I�)�-,�W]�_��d�Q���F݂8���T6s�6�C����� 9/��6n�h�G�r���g:\�s����1Nw�b�&��'��w�\uءQZ��t��q^��0�{,1	H����f��݅%�I|.f�n4��m&����Tc�?��Tj6�Ё�z�e������A��_"l���ѧ�/��إ�c<?���Xr{�)q&�ˏ�A����H �;����곽eR�}8������dLhS��\ug�s�؍��\�7�.Xޠ��
J�'?�߂
�|]΀��ĄO�_�Lú�>�C��IG��`G�J��"e�1��I�; V~��~B��)P:Lwz8�+���/�f*�9���kG����"���}���̲"��ahm<�c[���$NRDKì��3t��Q�A7�P�1�]])D);��
�͵ẁH>�|e����~K��'�躑��-jo%̓2�EJ&-q ́Y ��sGlJT�	��,���hH�,�,��J��B�am;�A�K[������Gw�g�~�h����i���R�O��H���J$ދ~ �Y����ݥ`�T���8V�>|%gs,M���y���{��
��$'������usE���=�y^�)팰wB��b��T�)�G6�#�z{���)��N�#�!8y�亙&*���4���0�$~��8п��z�k�/0L�ȭ�^��z䁫я���������՘������Z��‒y��(Ff�D(���(F�8���j��������^�9��8��'�@�ܻ�ݻ�G��\�7C��W��(����� ��?�v�1
O� �Phw2S2P�����H�`�w�p���Ӽ���ڥF���V��ТU	�X��q�����n�7�^��{��.�5G:�Bw�,#��x���������?5.�j=u��&pg�~M��RFz�S�V���u	GV gP;kD�=C����5�|�p����PM)P���$c��n>£�����?�=e�W���K*NM��Nv���^��a� D[�YZo�Gw��և1a���wڛͩ����y�[b*��W��W�	��af�/�[��-4�RзC$��(qb�iu7�����B	ޚe��N ��w���C;����2?L0n�'�v�_�>AX>mu?r����X�#���]��ץ��yj(�QH����ڷ�gJY�"֜�2|P�9<����x�N���@5���1_�5mֆ�H�<.N#�9�=���� 0��f�9����o�D���X�����g �"�.v�~ږu=R�OR�5�C����}I��[��-��"<t��w.�IJ���t��/��lc��~�3�^����@�z�D����'@s��ȶ�N{f�&'�fA���`�!	>��_6�?G��Ϛ4i|&1��4���`Ζ;���"|���?,�e�=���2��7xz��+n!���aѷ��u[��ƪb��������<)�lBK�YƏ0�LPg'�8 ��w�4gE����s���E
�)��t�Np��jڵ�5v%�j��a� 6����Ɉ���<��+ktٵmF�D�$�.j��.j�J���<�q��6^<O���L�
m'�r��/��//=��c�I�?���.W��� E�M>�v�L��vwږ�[(����du�0NA䛐��9�G���'��Mu�hۃ�nȇ�
�z%[�����{�Zo'��/ZD�?�+�IX�ye~��J�:b��;_)��:�,�&��ʘ��.ND�P���R���	6ڢ�hA#AD2�o�nɈ�4]~��Sq���a���-(ׇ�{�8�]��%�Ko8���bp83��%cp[k-�6k�k؋�����WK�dr26,�i{\A����x�M�|�N�@���������zx2!���4O~��U��bc�{��P8�|P��3�b�����J�� )�&)��s���nT�
��e^�+��489��\2 ��'����ͨ�+2vn��I�9��{�J��p���?&�{	�tP��	�st�-�50�>4���`r�����rX�]���Y;YN�����~&�\�^����2C�f��/l���|���-��g��|#�G׵��(���5�0�V>:</�RmTҶ�e���;w~3KX�YGFr]�[]�lQ�3�]�?�#G�W���r��
�sh4�?N��(�+�<�#onEM�6Z|Ck$A�~����4�	V��y��Q��˕|:���-�a�BWdF��D۞/��)�U�\OT�N����Z��=�9e5��c����K �սÒ��!X���N<�Ҿ��*����s��n�J���n#�qG�b�>\5+08)���O�����>y��O���)d�"����%��]"t���pu��	1�7���ȗn�'kch��_GM��A�y�� i�tu/�?�����NYH�࣬�����n�Zak�2�������>�%�� ��`��Γi8/��h��2�Vʫ�;y�	5��Ԯ����)��J�J"�?���Q�;�Jb�넙*�P*�Ȥ��y�𻧣,��C��Ω���,ڞ�bq7I�	�I�ǅ��?W��,QmC8��	|�zǋ��M�R�=��r��H.�ٺ��WB>�D/� _�F7�`a,������xQ�_�h^�hVM�cBT���T0>V�
%^���l����T8�Pڶ��>vĲT᪳�����;A	0O;ޏ�Y�'�3o�NHa���I�K�0dd;�|lp]VB`��ҖwL��U�����x����y-�.��׃K�}�L f�.f�z
 ;Ǖ�ݴ�X"R��&Vt>B����U�?��`���2	v0�J�ȍDSwⅡ�
F,P�_n�LTX$]��AD�-x�#�W$�,��ݪ�ܼ�>���6�<W���ˢn��2}�|����gB�X�.�$���$�ǬBc��V�G>����28u��Ux�M]�e
\�T��$͙8#�1��׽�-�wsU�Ə^�!�r�'S�ɫ�!N����,1�&!���g���Bʦ�qa0nm_�l��x��~��=�qn�4̐C���n&��=`��+�ѐZ���n[�@�s�r8��ث�J[^˙�o]��`!��=
��4����iQ=�d���e(��"�@#��m$:�XG7�������|]h�e�J~�Ƴ�53��ˀ�ߌ���z�o﷈���T���i���pY1�rz�/a��'� �KV��8&2Z�b#J���uϾȭ�j"Z����H�z����-R����S,�?��IlP*�05B��c�Պ�Ү�d�/䱔��]A���|�¹�1���sqM9���_u�E���c#�1�,��ڎ���o�� ���{{q2�������:��:l26~X8QM�>�/�j;v�/)�ԣž]�Y��
��J�a]�����g$�~�c��/����
��[��n펫�"�A�����&Ph���~��\��WB��� W��8x���Ʌ�<�ʐ\�P��K�� %Kެ��Y�$��{S�E,��1��X!s5-����[�/�Y��� 
1�gUt������ �RG��9�T���o�ӛ"؇'�/U/��|.�ܦ��x~�d�b��������;�=Y�X�%	y�fq���*�h~�)�S��,:���-���������9����S�� ��-��e�PrFg����y�"��܄�$��Y����ވ��s������vH���ě��oK��38��́U�H�Ⓛ`G�|K��~�@ �[[���S�l���m��m�Ʈkd߽6�U	������3�����_u����X�Xc�iYg�ʺ�+	'����j����ԡ�H�`Ç*۰�DE�\��cO�7�w1dFe"����4 L�U2�������QWPF�Kp�r���#J�ʄA�sR�c3q� ��L� �Hp���K��?�����0���]+�Mmsƺ��h��_�~y*�+Ł�E����J�Z��)}�u���B�.~�X�#F��{�{����E�vy���}��]����?? �I�#0���G#�]WF��=ƺ9��gf"Ik�P賾�J�ӿ�R�5���������<2��������.te��{�~�eP���T>�[5�
��,�g5��μ�T�ń4�ֈxG�U�.��x�ln���/}���� ��P�����{gT��n��'V;�f�C9��FN;���b8�ӈ��D #`(��)���K�9����}�6L�R��0�N�n�X����b�P9R;����؀6��Z���6��^���0s-sXQRt�?X�4+�����L�Q�gx��DuC��'J�̳=�E��3�L=���]j��q�9�r@�BB�N�?��W��L�
Y�jW�"ȋ�Ӆtd�0Q/HѦ��H�t�3^�r��^�?\h�E�uy5�s�� ��kɒ̦��}=���W��W��?��3l�<�`>~g=������7s�{`�L���KT��֕����k[}$�� �V ���R���]�����q+F����
�����3l��5��֐6���k��9����nUѽ:�E����(����&

z��Xq�Q��2�m����V��_Ԡ}������7Ϗ�&%˹M�� �o����a��ū�Ϫ,�z�}焑��V��Vq5n��J@�Zhqݨp�3�iK�{4�'woi6�]K�Y�	�ײ	w4�$n��3��]���\d#}��!2@n���KLw(HCR��G�3_>���t�$��h����o|D�y��"B}A�!���Y	�
�Y0;��W\!��L��P��|sy�EFFc#�Wa�!9 �{ðt m�IF���	��P��(�O�}���$�� ��ȪX&�6�c�y�g�M��-V|�	��,F�rL��똩&�/�c����u�UǮ���h`Tg)a�� �pAwx6D�J}�H�z���h>�����`�,�����m����Rf��pL����q=�����R���;� j���Ft�OD!̌���E�'q�aR�[U�L��x� ��fiж�$KS5����q+���I=���R���٪ַ�h��%u!Z��,�&X��`bC�'o/�8;�Ȋ�9�Uz�T�S��[���ݡs_M�n͙m��T�`��q�1/�+7a��%h]��iէ��N��S�� @N`�Q$nc�O麋�kMm;a�"�tk���)�p��wB	�R n���XnvJ�Z�"�¹�o��,g����jv�@x��گ���V@��5�&:L)Hp�s;����"0��#�&A'�kg!���A�6�Nt�w�#��ET����!C�<�������*����1���<�+�`$ߋQ�݌-� �\�H�t�f}S'�b�o���"N߰1�n<ÜΠ��3�-/���6�R^!g��hy*�{YdtAA����2�����#K�s/�J�*)_[�5�XcLӹz�zҗܢhҾRق��p�����;I�Z�;&��:=ùX�I3�xG��x<:4�+XlX���I�X��+e��le���~��9��@�Gy�@O��Ӓҋ�k��Ұ4j5���m�Uv��t�^�q0�����ˀ��!+[�5Es�D8���f݉������j�\�^L����}!}�61��8��(�[*N<c����:�u+�8�H��wa�f@�tvp
QC��a"S�~�lf�a�v�O��W��2@����=Q
�^ΒJ(��v�ވ�);��v�a����8:>�G�nCž�da�!,���ֆYE���%V�u�Tu�m��6�<�vt���O�a�ʪy]̈́��0>�q�������7��	.!�(�=�S�v�g�H��1Ж�IO�S2�
)	G��-O6�ͷ3vd��,y��D����G���q��|��y�W5�aip�E-*��A��sx���h��uI6r��o1ڮ8�o֞��[�N��*-rnZQ��^n�e���2~Ji��K���'����rjF�r�I!}e�=x���Fa��^����J<`�����v�F��94�,\B��zX��^CN����zi��xQ{�(�m��� �^j��%#�;1H���=_FsfR�иN�xu���r�s�Gh)�u�$s�pdb�x��~�-Uw�6l"�֌ۚ�0PUXȿ-!�>�E���X7�X��[�U��`FCPT�	�U�_y�TE��V+�"N�>�xmn!����O9*;�'j�[]C�Է_�u[�ӝ;fK�Fz���"���m�*>���Ɣ���눼��l��������P�F�a�~[��S�t�I����Z��>��/?\U�1���������D�B3���B
�{Y0�
L���B�{R�(S#��4���=�'���]��S����E��bT�����>�ba��4HI�@�I��e��:v�K����V��;X��& �ҩ7J�O��Ft���ML�^$�
�6g������$��Z�6WYS2�dx�8l!=��i�o ��#�P�����J�J�{e�2br�?��L�y%�x4��V����߼'�7pϯ�E¦��4a�Q�վ�qk@2��!������䇥,��UW��cs�i�_����,u�PJD�+��6�)}�M>[*�L,�D�Eq�}��]�~��)����zNМ6�@���a��(���_b���F�Hu8�Yp�����	�)��p�Y��OJ�:��5(P�c_�c98�C�V(?c��Ï=>�	\o��AACG��F�/®Ma*,%x^�f`Q�̽>)`���L0 �.x�F��"q�U�!MY�[l#��($]@�%o|?�Ab��x�W+�0��~xJQl䕾�~Cv�_}. H-���ݯ�F���P`��A��!�H�֌C��-��t
3�+}R.#�H�����qPئW�� �AG(���]����jbb��s�%�U
�\��"f��Vߐ��loi�����o6�m�Z��l�9�-��`\�t6�0�ZBq3�¹�T��=��p�������k�iũ*���i�+�\���ސ�o�wf��wVz�Q�u�RgS�_���7��wl�hKSC�e������O<I$�'�&L�w�]Y����ƪ$�� ̌oIor9����i0�6�Ǵ54�e�c�Z��~��a%ݔv� �ǖ�J�K�4���ƶ���>@�U��Y��1n�FV�:&���	����~7U�V� �  ���
!�DL�j�R����f����Ԟfr�*�U�l.����.�����?�sXyb�{͸�mkD)�#C{�Y���O&�ߞ�]���d�ҝϩkX)����V�&��{�z�>'��&�{�t�
��Ь���DL}G勹�02:vb����fr"N��/x�x��ɖ������㰒r������x(�����K<���cq;e'2ʎRFC����L��=]����;��A��)���s�U��ԓ>6��VQ������5�9� Ϩ��|Dx�U�읫ᦡ9^�y��t��>3i|��Y�d����P	���1�	��E��GI�e!��ߣ&�ש)��C����$'��i@�]J!������ꤥB��+��t}�~���ғ;�q�%o����<�C��3m��8�޸��~ޘߔc�X[��ۣy��L5s�J�_�:
�5��Cf�g�7�)����ү�v�#��̈́L���r���ts���t����s%u�����/�e·W�=�7���*��x-�.��x���}�����-M��N&:`s{��)�]9h�>��O�@T�	ةW��LPo�H���8�Y>�E�ù�Z��(��݄�MX@�����A����]��'��%<��"Vx���+����Ğ�^���ݫ�e)Cq��+�fL�Α���b0~~�<KsCa��^���5MM��gU'c��f-p�����<W�T�t�v�-��P�Pq��1N��_�_i4
�3���(�w)5:���ބ��������F��H��=�́� ϥ6���*vn��H��;s�l(��W�$iS;v��r�[8>&������E aqW�io�'��5�aO�j��G��[�����=l�n�&�����d,!Dݝ�2$�!�`�<��(���s!*~N@��FI�|j� �E&=9�t(�w�|6wo;���uSv�E�nTg���8J��ġ���Qh�{�<,N����j���IN�Y�Q��nS(�`??wc Gt���
��Ӂi�V�$�k�;��-�~�"q���	��rM�[��J�,�ǒ����CT���HR��Y��M���I1��OT�p�$c����^2Bt�mD�Dt:�	|g�I���W��#��%5��\� dKإ1�����8R�g�:�"қb6I�����s�FQk��]������W95NK��Z����)IvRˎ���8�>�I׵�ev�P�
�k�Ŗb.�k�(�B�ɲ�x�Fm7Fm׾lM8'(����C����5}����9x�����k�0�<
�W�%���B�J����h$j�35d�fA "}��g�����b;�y��K,��{�赛 ۭ�b-qNi�.Lu��/�d��^)��,��E��*س��d�R:��sw�'����v�����U����L΃Ϊ��� ����&Xws��{d�y��<�5:����wMHK���n%�yj�������a�ɟ
W�u:��W�S�4����z57��.��w	տ6�_wnV�c`(�c+�;�B+>����Ql�T���	{�,�4�N��͙J��˙�/�^DBג�S�Jq�a�uG]����=��\O�c{�2Q��<�9a����ǱP^��Vo:���ac��?;�֦=w�ٹ��ۯ:_D�y�[��L����ß�`�>I�Ic�Z+�qՄ�A�3>*~�:�����gV��a�h�������p�WM����� �]2��OQ@�_�� 0rZ�a�C�x*Ĳ~�~�{�)����Ŵ4B��X���>u�஭o�cOi)Z�p�s8ϧۧ5f�uk�=3L���Pr]�C~q��tZ0]���V�}!Y*��xܲ��n�ڦ�9�ζt�/��|�	E��9�e8�MgO<VP������

�'<��f����:��_�ᣁ�DJ�ݠg���k�����/T��[��ψ&ɂѷ�]��ͨUך�iQ���,-PCz���"��+�+�蟚�a���m�o��Ą���jV<�h�HC��LH���w��x*��<�gMN�}�]�?ѱ��h�Q�vA�;���� ��4'A�x8��.][qtީC��c��n7/Cmak/�5�9�Wn� ��H�~n�n}�:!L+��368��4n0iUT��%��y��
L���R�����ɞ��g�BnZ�,��%tJ�c���!�чS��>��'���1ߢ�Zm�����nر���Q'���lO�;�J����R�Ap�o-��{0қO�#6��ۋ�@
�i2�?'�Gh���JvV�_�]3��ϛ$��h�z��+�%����&vu�k���1�EgȊ����*�-��>�A�Ww}��	���G�	�YL�mh������q	x�<��t���G�4��qg����N}��ŀh<o[�?i�?ӭ#��6ޡ�-r�	;�mm�t�؟B��&�� �%vh�P:F!��ߏ�)�g�m�"��)0]!�M0J`�'�jWQ�w��� ްAՔL�)�N|.Y��q����]���������0�!��A)���� �'~��5�8���H�� ?�w��tF1_o-�KW9�CW`H�@�J��,�+�%�����ƑU�á��1��`��(Z/~;c
t<��i���!i��O,�߿b
U�#�Ś���޷Z>��RlX�Vm��|���Q:��@�uY������J�J�a4�S(ɷn�}rǠ�QN�%�o��Z��t�bA�����E6��$"�^we뙚�Y�<��ҟ�����ڏ�T1�%!53�1�N�;��pWW���v���8h��f��\XB�֖�O~��f���f|dR��*6�f�I��-���6D�g���S��Y���/�{G ^�Z�(�\g]�����qP�ZK�f�a�@����_�d�q{����DB15�.-������ya�Qh���JSHR�|(��l�w5����(�cC`�(������f�8�d���x�L�����YЌT�@,',�64�!�'5�������_;9�eJ�DB͙��:\i���k�x��>��7]� �'������q����D��up:w82����"|f�~�=�=p�e���QJڣ0i��)�U��\ޝy��}o�約S
��I�0
Jř}"̍��5f�K�2����me�=� ��f���F��C��C�D� z�M�a"�"k�/�jJ��` �kĶO�z�����h��ȃ��JT�p^V�I��h�3��Q���K�e29C�m�<�����\Q΃��p���f6�[Z�Y{�"�G��9ŁX+p� F]#�U���k󹉳O���ឭ�.�<�ΖS�=
��e��.N�?�b$a����)b��2��^3�Ԧ�'B}��ho�Ғ2�uF��4�VR���M��[����$%«;"��`��	�A�7ҙ��Z�[Ǽ�[��à`; �.{� ��
�d��&	�JO�lB[:W d�(��m��Q��$�9db\{Q8\Ki~�Y� �¨�;��#B�)�v��B�$���VSaILV!����\�i%�W�G|h����#�=lv����χ�*�G����|?��b����S�Uec��/'0C�&ao����X�`F߃T}�Vڥ<<t�Ȍ,u�15�����F�3�|�^*�q��k>Y�:P��lh�������H� &͝/����Jy<�zʗcd~_�L���w&?�h����F!
*e�L'#���
�a��0��hNjD\��6j轨8�UĂZ~�(��Y$E�$���"z��Z��`$��{�DF#������F��|�����Οo�x	�/���eGd&S����®��Bؗ�P�I��,72���{ki��v��w�q%��f�����[I%����������f�����Eb�%�F\Fka#�� �2_�'6����w	�[z�k!^��nD#ͨ?�.^�SvMn���u��u�������	����i�1P�$I(x��(��a��敨I^�7L���Q� �������]����:���xRp�z���mHH�R���!TQɶi��fUs����M�%�N���M����r���{�8���-�`�}�1	��,���~n�m.U�7D5�mr	ݤ3�t��-O.h�6&n|8(f�@/= OA�a���~����<��b,������Yka��N�8 �΅�U�oĭ
0��5�,�*�y����D=�ޠ��t��(D�����c%�)��j#�e���ܔ��o�lT�~@:	:�m/��S�z�_b��q�h S�O6��Hi(\n5�E����Uh5�"�}����>����U��`k��oٛ����4���g�_\G�5�K���Ej
�<��]���E_͏���@q�>���Ҹ�@%�����4�����^!�Nvϭ�!���Y�ӇUqak�14��)��^�ػTd�Y�A�j$-�f%m����'�\z8V'��@KE=2t	Ҕ-�и���@��{o+�i�J�﹩[WR����]���� ���7i1��� ���n-<ƨ�$�����<�	�}�5���JɩT�j�R��)��N��b(/�f1L�T6p~Y���M�Z�.M���N��\4��!$mB��թ���P��;�LΌ�[=V��� �-%sў�� q*�WaC9=>�%ܒ�3H�}R�ّ�^޶� r�~������+����n��ls�$��r�]��-
��~ʾ��&UO&��l2	�[�9#ec�(�J���KkQPțJ��o���^R�Y��Բ���f����%Q$�J����8y�M�g1F�$L��m�z(y�ᙉ�Vb�@���<e�d����@��/ө�#��-���o��
#���2��A�w7�c��*�����O�-VC~�A�CGi?�77�x[FOl\��h),W��-����xݾ����;�z^NZäh�����v��}���R�>�v���h6������;�\ő���D��P�j�yHr|�u� ��K9ht��e� ;Cw���g@NIJ\��n*�?�co9`{i$�f�Љ:�`b�T�T�W@	�5,��n� ��{���w2�[�����'���9h��<����� $?�L;4*�עY]e3$����$'j���o��
�.��Ę�1:�ZB�߅��*�n�$�8�.���yMZ����[��/v�J6WB-�ʓ��X�g԰�O�:����'��_"?��Z�*Nj>��Rܪ�2^�D���d~!LkK]�U�Ww�i�H_mr�R+�����V�g���	��@x�bn��Ys��hL��eQ��J��Sh���/!����O}�Y:�g�Y�S��g��w�D��@���:��W��ps�[N�##���%�̓{(d���̄[^�a�"Z�H/��I?�´��)�R�= }݃<�3e3RŃ�������7�<,-T�;�[�gr5�&�`Vu��t���·�$ڑ�-[�Xzl�����{O[=ͤ�yRt����8܃wm� Jd��𬛞��8P�ٚ����?b�e���	�Q`}���{���ZI7����2z���(�A�(��Pܓz�[m�%���2&���>��[��8
�J�:ȗ��Ս�F�4�zk�P�p�M[��x�ϻt�2l��]�M����Z��!X���S)tm/OAC�.���/�p"��C0$�����{=����㡄JS�7�bJ��:�B�P���Ah�g�%]�I�г2�g�k`���"��,��
+Rp$Y��Yj7����6��QR�"��x_AΦ�'���m��5��Uˊ`_O�� z��/Z�v��Rb���^��������x�����Z�jͣ�Fӕ ��|ӂ3��Es�3���)��T�3��������Z�����m"a'��5t������5� *q�҇��*;0��FT�z�]D>�0��c��_[](yK�&g�RJLN_���@��8��8':�MjNd(�����?�6�U~�ͯ���J�e�w{��B��Ã=�Q�ϑ��S�����f~av����d+����Ia�I���_69ބϐb�S*��z�X����]�mR]"��͠{=5�����
�m�D���<�-S�T6��;�����>qy�������ƌ�٨�����NA�L`:�ē*X_l�	�}L�\A�˛�뫚a�M� �� �;
�g"?������%�F>kl�6P����Y+���L��_ѧ6깦��n6�/��e|�����F|��/�-:#������@{�C�q+)�f
 {c����L,{Q%�Z�B�Y0�-�$�D��ܐ��0Q�~��5�h��i�C�ZՀ]T�����ha��v<$4�k9A���b&�m���)1Fn���L��/o;5ۥf	q��(�t׼��o�_>!DH~���z��3��w�4����n<���d�=�	t����ZSi���	���0���TA����Xb�<���ڃ�' �Y�b�Mw2��W���s��dKj,��=<o�wgc�v# ����Y�:��"h6�>��Y���u�hN�[�)�E�.4e��2-�%+Z��`�1�c�F+I�������u�ǄT/yT,�0�#�o����M�֥`��-��Åkg�V��m�q�x e�c�Ք��[�!���o������ڃ��XuQP�'(>�y,�N��������4�$#)�0j���3)KR�S_+���R���[����[3N�.�&@�b�H���L�	5v��]Y�f��ޑ�6Hw�C���s4}s6�M;[�e�>�v�D=#�v�o"��+�!`����6�j)���� ��h�)Q�|Ud�0OeM^|�������C�BF[�P��h����W���U��R���i3�f��m�"�h�F�i�O"�IEcVة��ǲg�K���^�2L�I�[r�F;(.A��\?�7��9�B�_AB��W'~ca�����q��"�Oy�� �c�S�^�'E��k�{��Ш��&�xE|�=ꝇ|�����	븲��l���|� ��j~V�@!��L�����e�H����64!��:u���&������^�qc�Y�i&=�K���P��)��� ��!?#����L��ѭ�$�8WZ|;��{���=r��"�=�=nm4�HF��d���>�=��S��a���]��.Vl�Š0B>���u0���I�N�Y;�h��@���&[(�u�a�+�Qz1��Q��h����R����vm.mR8ƛ<��0iA��l�7z�
��3UI붻�C��e�f��� 6b�3.����Ϯ���;�IH%={˂\�B�ZMF{�xQcl�f�`2����'�ף����� �v�~(�tx.y�T>]������z#s�M�z�?e�i�=�� ��Qw�t�"ohq.PV�:�swB���27���ߚת7�2��ݕO���x�k�f�
ѥf��3�T��~������A�����5��71��kUX�\��'QͯCa�V�tš���8�c�ޜ���4�O�&=���E�1���ӽ��Tמ���~�/�Hbi�W��=�u��Z���eǳ`[/5%�n?�b.�d0�� h�|N|�����/��F|.L5�׆�;�v��/� �9����.�� :���?�`~�U_)>�!�������3��������
̙��b��L�㘻�{szT�6��
EO���bM�A��wbð���܍��u���b+KU6.�>���y�o`���L�^4t[�$6����}���PD��#�d�p��?H�%;�;�U4���(��"Y=���)>T�^�T��H,~�(�ն�=BR2���^d��!ܣ�.��xT�)pr��� �|����: �_ErisR��:5�
�t�g'd@���e#[s�xr�l;�w�<���V��g�t�T��ыx{�9�&��,�|0���pW��>-�U�z��_�<�5�D������d��}��UL�O��Ck�3G�)�)����7���>�B�g��9:v5Q���G@d�5&�˵w;=�)1"�eױ��'kN��������)�|��g�p�o@̓��7YC��K��3������3��G�����r܂8��ï�NQ��vޒ׋��ô���w9���|+��u�f�'&�q�'�l��!
���Ybxxfˆ��`^��KN�#Wc��:�0]�H2���$��$�uJ_�J%����qb����!�)��&�[J[������I�ċ <;����U�w�ݲı�Q���ρ��tj�"[��-�d�R<׻�1�>v?o�ܯ����^v|�b�vX	�N%��Yx��@��S���Z9�8�Dzg4�NA��:i�(���o��B�J ��l�"�;NВ�Ƨ����Rc�efºh�y��T��O�����$�8�5cH^$�:�f>#�gT	1>�M�n��a<�U���oy,�Tצ:�$f���T�T���ƞ$��Qj���8���mW/m��^g=ţB���_�ֆk�3����W� xm��+AVw#�6�E���no�����,�ǳ��>��3��V	��t\Q����0�2�d4�$�g3�a�t{�A!.~m����(� +����'��o�����������A�k���`)��z(F��tq��vZ��j̊bhy���cpw�p	����|,�߉^Ƌ�~�tm/m�0�!�\/	U����?S%M�f�nj+e�=��9�����0u���N��DF�e�q�GtFw6�X�v��n�:���֚�����xf�R�+L�.H����&1\߃(�$�p�:|�-=��T�o����0�=CR����\���P�Ќq	��]��M*gA�^��A�r�����cꩴ'AC�Ok��Z��l�~/�K-)�rdr�]��(G��������{6B&ȫ��9�k��=�>%1LiS�]�!j�8��{}R���d-�ᚷ��f �	���>�!�""��p���dD�06:=�	c�þ��K:�83<T��U)oNf|��7H�����z���l������J�x�Y����I�^]3��t7.�e���nJC�Q��jV��V�����pGv��I��G~�/�c���?�;���dI�ќ�Kp�5>���Uaj�c�@����6~����$�f	�\����N*�Ir��ћ�&E�����O��#ia�H�h���z���s��}Ҍ�(Q�'h�Ōs�*���Z�\ �$��O>�16���VN���>,r2<X���<`#���<�� 9�"��6d�އ_7M�o�_�W�MN�����!��	#�p���m�1Z�g�<$hB����f��]8!jq������{��{)��늆���pe�*H�ɖ{�[~ ��-l��_̂3�'�8u8�S�/0�W3�6�!��a_����l(�;�졒)'p��	��$���%QhiD� �^ۡ)�W{�N:�9��{���k<���R���-�(���H�~ђb�p�Aǋ�Ñ�z��H���N��J�~��k�+N柳����8�3iCT��n3D�FUb)!��$��/%ӧ���:i�w|jAĵ��Peٲ�g��F�ٻ@�T9�	`��(��BY%��G�->����x����>*��ܧ<�>ʹ�.��3܆k#J�6w!��[���X���n��`�u?-A<�������C��B�m]�OA����ق�2µ���4����jr�	ntx�ˬ?|Yut]kU�B�7-��gX8im�r��-o�����yS �W:�NOd�|��y�)�D`y:$�E�}{�~��D0jw�*u�:h3�o�?��7z� ,#��P[�#3(�d�ܷ�!nް�����,x��3���a��J�Ӵv��,�v�.��#�:0��s11ĳ����_.W`1��@�!�_@Τ�� AY�Lc`?o�2�J��ɯQ�N�g�c��U�w��%�VC^,�hI���3L ��ّ�y,���	~�V�\��To�ҩ
�hU  �^�v��з�3��=�V�C���1���m���u��&��#y�`�[�g<Hr�la��q�������c��1�9�L\�5ᕧkwx���d�����V�������v4�#�;��΋41��O�ԩ��/~yɊN�1�0F�q%�o6�3A5�]�e��d� ��w��@�r<�2����Ёئ����	�\�,��	��EǗ�h�~�D�N*��,B��jE�1�-tZ�B>+/eҸ��d^�ޠ��)�?�H�w3��Ă�V�T�2w��ϭ���!�o�I�R�)�Q��s=wx��F�|�TN6�����Oq�3�u�����rq�0�c�%.�/0���~��o0��&�0��]Yhg�=����C�H��u_�g�:_�"��^�pH@*H�-�>���G�� �d��\����C u�nz��y��+̒����Ӟ�U6OZzx�� (?L��8r<�X'���a�U/[��>P�ܪ�aEC��q���@mqmrI� �.�ooD(N����[����;��X�)c���.K��\d��6�_��:�q�\��B�rh�%����nDL�A�.�~��L��<W�������:�����@�X�9�2y�Ů"�ty��Yuݿ`3�*��^-ftڨ�/���z�����f�M 
���"�e���:� ڹWz����+��RJ�%��hi��>u�#i�][rx�$nŮ��p�b��1/jRt��Q��,\�uK;W�V�KMRJ��B�#�X��E�y�}�%�m.n[�
lq���`cy�H�ߍ5	��-|
�{\�HV�0QP�J�;{;��į��년��$,6о���ȣ��A��^�O��ewr��>�=�О�H�Y�>�\�G�ƻCr����s�dӕ,�,pX�C>}�cm����\�t��ջQ�c�cPy�P�ժ�]l"Cg��M�s$��?�pU�����o���@��`��dhc�6g���D���jń6e��'O.�&��j��v��3�������תV�ej��oz-&(�}N��m+"֛J�b<���x���L�7g\_��`�����>)ܹg�nP�޲(��}�%���J%�JKmĮ7��u ��J	虜�n'$vT�U��'��"/JՉ7�'�il��PUI͊�*L�����X�!�իs�q��<)FL��7?΋!�6*��o�(�J6�g�^��bpl�U���Q��*v�pxշ^�<A&͎H�hKwd/,6�ݔ>Bmc�_��$�7��B�� o�N��,er�P�H[zI�q~�%�ۨ�y��C��0Z�#ӱ�)4C~�����}�����D
�zn.�X��(�jhkw�M���滁j���e�=;[��� D,�]�UK��w�BDݥ���AM8L�FŞ~.ߔ4�ކ��Ot~��^��8����yr�����]r�n�����\�$W"�.�5x\r���u�&Y�[lu�
� U�|w�2n����J����I�O�Ĕw���UP��z�~������KS��m2��GT<F�y��;��v�i�ߦ��&5��������@e�vh[�Z^��p��Δ+8����䜂 �D�f�@�h��X�*��3QxP�.�A�?o?݋7c�-�'W&	���t����+��H�ᛆI��)�K��G1D4�|>��d��`~W�SS�j�ehfu�b1���4hQ�s�#������-��ک��c��KC�}�[3(A���S2K�Ͻ�h�Z�hF|�^5��k����X�8��rZ�1������M��Z�}(8M��ϥ���h�F�_cQ�z���,�Mvj���5�Vu��ߗ��"��'��`mX��)�0K�� �I���}zc�>����I÷��A�ź-& ���9�K�հ�7�<�c3~�CftUC���.���C�81�6ʌZ���@�r+�h��/��,�!D`�G"����uN��RKf����DF�Z�@���8�'Y�TvO��|��HV?i �y+�A뺚8湺�A��e�y��c�$.S~�Ho58�����l�!�V�k;.�Խ���_[..<�2��e�0� D�D-5��A��*R�6v�i�f�'�Z2s�����s΍���;�0kN�'l�ؾ+Ӻ��d��!������8�Y70z)N}`j��
(J՛zah��|Ę#Ќ463�0'"Ā/I\�گQmc��m�����w�Sv�@���iي��dy�zDX���`tu<ޡN/g�����[4%�z�����}�71)%��X���ݶDބ���9�@ߣ2P������B���>�/���Žd�3� w��B�7j��1�d�@.|qCiԒ8&�/����z4*�&���� �#l6?���{ �ET�~H�N���&H,-#,���7���l��-�*�ÝE�U0 2U����!��7�-d��]�Z��S��<®��Zl�+��M(����l[�f)(,�>>N���=�$���"���N^'��8l�$��'�gy �V����H�D�T�X��@�f��'��$��	��(�f�A`��9��_5Z��末�7�����"����J�aV�,T�����r��XS�5���e	*����)J�85�S�@�f9����Qk�;g,;n�
���=�8�J};���f�
��o�	�G6v�]�k5��v�G��A�Bb�-8K��&翳�0ZO�Ѥ�[�Hs���B��(#gU=�t��k����@�ME�tzN���@X�PΏ��i=���>�!�n��`���V�'�T�e�|+,
d4�O�~~Ү�by��uj/��+����'�X���-ݺ���۶j@��s[�kh����e!YJM�Q�[���1�뱒�P�Ձ��@�{�E^4��_�ƺ�9���1Sx�7�3Y�qk��~��˺�l#��������R�����Z�A)�.��.)kܷ/�)ZH���|2�7w��/�ǋ�쿭���~��,�j��XC�L�����d�ҥ�TN�~r�,ς�kx���U��>��cJ�� h�T����my�% X�4x��w��#���b�LdƇ�f>s�z���H�9AP��*��R�!����!t䝥c��Ė�kt��B��*�D���R2�����MPO����y��8�Y�Io�]��߭�N}������V�UҶ���៣����#�B.&���Zs��c���/�D�Q����aع�}�J8;��ߔ�L���8BP~x_�U����.��B/Nf�A4���{�.��=w��2��*�ފnf����W r����Ƴ�g\�{�A�ԅ��)�k�(���˷�!��uĄ�D����J��g��+��P�������+ (y6��˵ua?��i������$U�✺���W�C�\`4�"�����r�Jn�2��`}�R�v5`z�S��s_��'0���g��RԛX��P��`���A�g�3�|��'3���_��^����Pj#{���������z�$e��7���֚��>�e0�]��`��f+�$Ǧ��l�ު�����a��σK�T�9��WQD�s��T��k�S#���#4�Y��
����_)����pN���`�#��r�BQ��.�`:�쓺�ڟ�
�Uc���jN�p�Z��� )*��XZtr�����ٙ8_���않q�GwVƚ�,��a��V9�0���,^r��H�h����	t�v�p'!���|c��M�l�6��� ��7p�->��4i+��=�� *�H��_�jK5]?���F��➀�؝�'J3O$��Ō+E�e��_7μة�����t��~������^=�(��L�x���p_�"q��6(i2.�g�x*�f6|�[�`���^還O����h�"��X�u��n��߃�Wd�U�R�.��w?n=R�ԷP?��|�fBSH� A��h��q��QErC��(�p<�{�-��Q$&�$ʋ��:�)&L������z�!NX�@l�T�\�&F٦D0�(N1��hD�4�:�_o�e�U�"�7́9���@�2m}.����װ���+Fi\<��Z�CT�4�*�
����-����%�M+>9&_q91�#e���e}�p
/�3,+��]\���ͤ�\K��6�ڊ�H1g #
�~�h�A�5�n�Y�����r�P�3WlK/"n��`�J�3z��a��! ";�����j"|"_��&����g��+� ��nt+�BK��<K��L�')T�|�ϕ	�Wô=�YCص� 1/r���Y_I����XD�:�n��R�05��m�w�xV���x��36d�B�4�Q�ߕ�̉�t�ϸ��1��o�M
�q��&	�������$Y�3Qv��?�ʴx������2D��v�u���Q�4���DU�M�[�!��I��BY낍��9?�V�f����?��0 �?��.����v��}��CNu���1��Z��1d���aCt�t1��]H�����)��a�����jC[9������p�� D��*�S���)ۨ�O�;��LV�3M�/m�X��ذps�Fod�?$l���"�x�Z�s��+�5��$S��kݵ�H�e��y ���\_h���_��ט0�q�,j������M���.A�BR���sWBnnn8u/b؅u�gP�:��d��pr��{z(��AK%Ǿ����ϳ/b�Q��Q{荞W��e&���c�]wt"�A� �ef~� ��4?S�,nr(6�|؇��_�N`���y^?'$� ��K��1��x/�G�Cݩ�,�GN2�m��M���]�����o���7�$�t��9ǂkዡ��_�"O�2m��B�?fC��26��(����W��/!����[��l�J!��T�u���ے/�
Ib}Tt���Cj�-�Z�]˗h�=����Ou(����S<�TMTx�Ӂ��y��������/>����e�v���&E���2V��J�M>����WBl�M�\@�<�ي-iSiX`/�0�H�x��a)���6�>D"��bO���Ҟ~�]���R8N��`4���E+�>8@�ן�1��9��/!blb�vw^��L����d���SڧOHy�p���P�a����y}�ͯ��l̳�M�P(�Y	ov27;Q�m}*B�#�$��z������㠺��������A���DsR(�u[��o�r�s4��?�l^XƯB:nkն0�؉?.�Z���C�"2�6ܔľ�24x��⡽Ҏ��(IXZ걔����1��� D_Rw��ϛ3��q�E�U����~�17O�jM�&�Dl���tpŔaJ���]c#1�)Ȍ`��ƻ��P\e�Bc�x#�j��6V�	��AC�&a������8mK$g0>ydG��MR쳌�3�k�߁ �nB��a��V��#�ai���� �'Rs$�#H�~^*�R�vW���>m� Q��S1[i]1�qjYl���x���M^��>�%_?�2�a��R���?+������/q_m*o���=#}��?��7#�����M?ﭹ^��F`�I5*��6[x/��_�{^Q�Bat�Ns����L�q�?���}��c�S��B4"�2 |^�*����dh��_}~��L����w���{v�<��A+���H��G]���W���ةǦ��5X)0ꯜ2���+Ԃ��6Σ�KmӲ�v�}j4�)��O=�H��f�A����ِG񊍩�*b�6�n����$���˽�Q"Pu��(XӮO^i�����w�K�S���pwt)Fu=Q�Y\�!�oH�%��J���kxgr���'����b��3X���;�e@��)��J�$�@�4ڨؑR��ހB�O3@*�1�d؉B)�:*�?��\��Yo�d�#r� �Y�������k�!3X��y1�"������]O��nwm�9�Ke��O^\���U�x�7Hl>��w����
bA���)��N�ڎ�@����ל�(����g��)-T�0�o�yO@��j9����q�!�������#����k���H�j���H�~r�琽����3�Q�;����	����3���� � �
Q��he�T=����/N���>���,zpD�b�Y��$L{(Yh])&Kg_3/T�q�v�z�+�����0fz��R�#t(��@D�u���wLK3bc*���ո)��˽�d���qw�ń{7���)��h�<8�m5�^�)���m���iZB��Uѓg}�J�m��jIBA=�SΘ{ݝ}�U���L��t7���s�R�L^��5i�-L�=�i�/���(,G��Qȅ����HP��of� .3O ���E �@��E"l��p'ZTD�u>Q��:��ttx
��C���~J�)������RS?�L�'��h����f�b-���?��Nl���Oxx�T7˖��d�/b�6Ή�&r�>"��~/.�h]��9&y����.mrN��·b�h)
��\��U��b��v��䳴�qVi�,&7��+$�Q��#�&� ���$��=:��I�Wݍ�2��ב��n�}����9A$�K�7m�+��3�Ͳ_Ľ��
x\�B�b��l� ΤR��M0ݚpsd:�2}u����;)C9�Ǆ /���x�[��v�A�ó��>��3�� �$�� �)Ik� Y��fi�^�(��~z޻7�U����c�Ǡ� hB�k3��ߣB.+���kʃCʘ<,�_�b�G�N�j:Y���C������ևdҾ�O�ܺ��u�T�{�� ��V���(�.O`A���L��z��a9ɳ�Q�#��BΨԗya� 9A58��S��wp|5�+|W@i��:�R���s�g��s���R�ߗ�02�~�s+qEqOW����)K;nc���#q�I���:��!-���;Ӑ�1���C�����.��
�e*��z�c0 Eϑ"7��G3ez�:�m����4 �T����H���Buo�g�l3���>��a���5;d	L=
���0��k&����]Eju�pPu�@���m��.��Pf���@R����1r����c��9 ��w+ds�����!,�5��>R���i�n6 I�9�� |6ه����I�N(&����$|�%�NW�r��&K���%$�T{k(ߗg�,������CF���:.�f�&r۔'��S-��{cdŬ�У��z�G���%����P��O:�I���t}�;1&�K(yz���S�Y
����G�C��������k#�b�R�i&\�r�A��;��RO)ul�����L�p?"�m�<���ņ��@�i�Z8.6'#j�C�;�Xdx'�w-�0��H)�Gk��z:U�e�������w��c�$��?��A!�ܡL[Р2.�lgX�6�!ߌK�����-�gE+y�n��.��Ǭh	r�w*ky���L��s�<A�i} �'�U�e4�z�T����;{��&w�����+���6؋i��|�A���%t��NDf�2vJ#�ѩ�����w�����eM}-�j{\-Q̋�hB��7N���Tk���B)CA��7�"Kr�U�%��4����@�kƳ,����^�)�K��nM���a�-�W�:�)�NG�0�a��ıZKS��
�P�-Q\TMV�V�rL��+�f�y
��d������7������RǼ���A��VJ�k��?~��k�,�
��J{�r=�p��(�cj�x"�J���E�����^��V˽tJI l����(�8gwk���l�Q��I�Q�t�s��qy��7�9�F��|�����ͭ�x;�°_�8s_�8~�����ͲҢ������SRw،`$�,�p�)e����S4����_�~x�+ـY��<�OR��7�HL`O�r����#�wQ�.�gؗ�=�Et7�0a����|Xd�n�����/]2)�Ǘ�O ���m¡H8��5ޔզ5w��\��TΔ۳�/u����P��Y"oo�����?�����Og���,'���-���z:�̶ڣ[�5c���>o嶀ܲ3=��!�7iq�]��ђ7ɑ���-���G� ��r��B�)ϱ�ߵL�IA��ֆ��Ί��9��ʙM��X��.D5 ��ʇ3*'�/��6n=UQ�+/b�1-G<�a��YI`�1��jS���l�E��%uj�'�H��.�F�1=�s�K�85�K�����~���j!�﫹���*>��(����D�R/w@�óD��*B���}qHw�O��́�םh������@k
>l���A>hi�ꎡၱf�l�ì_V6�Ɨ���C� ��6��܉�kT��.��ǈ���'BSj"ߦ�$`_��Q�I:JW��߈o�ٺ�T]$%6��T�,W0�=|l�V�V�6��OEDR�:DN�Q�`�O��eN:��?�kU°�D"ܦa�V��/`rI��z�r�j�'�#X|p���	�zS}�H�܉�KjQp܄�!N��|^����Z�=���LU)���ѓ���N��: 1��a�l|{�FY��G�cSV_���f����������0��-Y5@m��D�����b
�Ā����?����8$�MӅ���D��͘��S&�El�d&>V9J���I�?c���l'�{��e�m���g �>��/�
G� �?���+�-i�@�=��gN�߶#b�l9��ޛw�v�9�/'O&�w���x�2'jk\���ˆ䁯7|1��d5e9��6U�o*���?�׊ҏ���+�Ŗ<F������[z���K���/==8�l�*U��lN��rG�Z���V�F�=���(C��e֡j�����P����zY�?��8�U:N�V��S��)J��������#ݍmb`�ѩ�)�*���dJ?c8`����IȞ@�c�� rl��gj��3�
�_"�Y�Ɯ����q{)moTǇ���\K}���85Y=�&����`��Yfؕ׳�3��,a�s�89���Z��z��~f�"k܏�HW1�y�_Y���8��&��Erm<3��0�qU��W�l�_`%��a�F��e��颕�I�c��'/�����4�G��0��p+@B� 2:��b��\�<25.���J�֡^�6�n|)[�C���2�5d���->޳D^�c�q�M����Z��:���$��/�x��{�7(�}�pт*^������n�,VOW^
��]!@Z6X��q�vާ9oŽ6�*%�y��B�0M�9^?b�7�BK�z>�(�|���d-;�66qEeD�a��谳R��q���/�֝cm��L\�(����MAZl���>�(������x�i��
oR�:5���@�����8V��2�;����=�5^�<��{n�8�W�d���K�|F, �GPE���P�5�Ԋ��a{t[2�l=$RAj�'�jE��u���k񤇌�|j$
��E�[�d-��1`��� z��-~��TQ�Ļ9��7�\sx�#�p'�s��$��xJ�|�n�$O6)�%OX�<>��|�,��f�=�B���R8�{�<IVx�=;��kK*� Q7�)TO�A��I��X�ۭ喒#N�#`�4]�_�y��R�r0-%�Rωq���A}4t7��*��+��X��p1�7S�%A�N�2��Ңl��}'đ���U�;�9�n����
dȹ�=*�	U)�p��z� ~"B�08�~C#z�
S������T�"]d�~Q0���n:�t8`��	'w;�;R��������$��C�����?��s��~�˓�O��$&_��ˇK���E���B��]�e��/���P�2����2�7�����Ѽ�a���߫3�1>�(��LT�/����u�B�~��nq���|�~�tFS|�!
B	��]Ss/	����qO�P�BL�-m�'*{x��	��>���wZ( 0��e�^؟�vPK=�3L�Jq�1����1b����'�\�M��
��,��9y`f,�B�$Ĩ"�j�筨�؅����8\���R%���SD4�S>�kPQ��۷�6��@�#~Ԃ4�2��&�9�l����G���^'
����:T�����0KZ�P짆%n�t���R�� p	�i�u#��� �G��m�k�'�g�u����8 UL�˺���(;�?����9x֦��ՖGrN�\���QIA�ӄ����Ϟ���m���X��"F�Y~�G,�tN�Y��k�-����"^�V�KP���s�:��.����3EΑ��Thzw7�9V�;�HEd�v�٫M�.�/����m/ċF�2	�3~��o���� �+ܻ%�L�Z�$��8��x�(��@f�ޙ�B�?��˽K�T��.z��I��Z~����e}���P����'��)��|>�--ĝ�����'����oi^{�iT�"�3����횗�n%�M����q���j�<儖�����,#��jR����-��;I�d�^� �7 v�,T�����(Q��Ϫd`�+�3?�*{J=p�����YM�*ז��N$r��4���C���f� Q�Z
��N6w�����xY�b�/��d4�M,Vք�[DU��f9����[�'Lp��q�9-p��*�5�ï��R̍���H�vw�_u�p�վ�����%p(������ժy��Ƨ�|����D󩎸��O?la�W�d����ŕ�M���.�Ы[��/���/¬�!E�E��TOs���k^ ��.W����n�󢎈5�(y{�0��	�����.��kЂ3b���$��JX�J^.���2���� &�6�q~K/��:�G?�?��TrF��%ܻO�j�x��	�>vSY�YLx�R�]F��2�ۥF]u�2�Dj#�<�F�]>��O/Kޮ�dh����J�K�[4г��O �AH���z�k��. �U<.�2G��^�9Ց�������õָ����Y=�����O���������Z+R�I��0z
r�\��B�E��a,�9�y� �k޲�>q�����MQAM��#��(�ذ�k�w׵���H�B���U������m(�w�1��	��=fЪJ�gΟ�X(�Y|����Hk�i�e搱"Ql$�LO}��7�*�F��"G�PZ�^t��T���{z�.�9��i-��	�Ũ���$���E\�>�R��7����dV�\�#�lH��w����5���7��?�gb�
Ԙ|0H5�N��_D��B���)|h9�*�w��X �F�T�X�"����$��ەz����m���'A/���`�$�R�������WQ�;3�Ǣ���x���<���^�u	����ę�5�Q�p\=g$ �hFD+3(��-������W�;E����ae����CpL��@X�1Č��CV��ef�^U�l�Rb�����/�e�n�w���ǭvr�xN��/�}9~����"�@��x�UDr��Ρ�nJHg7�;@�S&�adV�ŵL�h��o�L���{Ch�Y�ڍ^W׊�h�7*E�x��Y�	���iy.�!�G]E~��zc����$���iR^_ي�BNJ��P@�އ"T���p3.q���'��� �Leu�N�W�s�q�F�;y��6��
^��Y��I��������U=X���D
^]�Ax�#�ӝ�8�(�җ�;�2����������hg��F�vT�� [ʚ��e��)���m^h>{@����p��	�T����U���<���ۇ�ı"&�t�0�x�u%H���e� F�1��]i�r�􍑄��чƁF� d��t�f"���=��F@�;�F�)~�\M������;��YhHpo��Ǽ-e|��Yt j�o�g�Bh��,c^WpF;z�
�A������߸�=�<�~��j��H�U.
���Wu�0WTNӰvz?���<�=]�8�Z�*��
/9�H˔v�~�I���Z`Tk��%�L 
�h�� w�y�:��>�A��� ��:�|�}皞,2��CN��b�I2B����K�GÎ#�MȅT�7i]��h�,��۫2*}l[�Y�5����!�6�7LK0�%�_{<\d������4Ab4fװ���cA3k�"vŲ����I^�}�mnU�K+�5��y�6����H�U�Xl�a[��U�=;Ω�cA���Wo������M�kr�6ȦC�WG��LWo���k��d�V.�R�h�jq��%�o"���&PTZ U>ð�7�Ʀ��45�]n�ܛBNqHԨs�#�MP�Q���2:�U�{�=q���:P��ᾰH�9��9-e*lFR��K�!�^W#���������1�P����8@EA��`A��ߟ��^����^�$���h�-rYg�C��ZE���`|5�.�p`y���D�B댱=?��q�/�����5��J-��?f��^,��w�K���냧W}��p"-��]��Q�q���M�~ /���A��Z5 
���>>�� �Ε��w\�a(<�jL�N@�oꋻ�K��|4;�FI������(ֺM�m�p�N"�Mxe�r`�~S8��'nr�a�`�ld)k������q�ʽ���橄Oߑ��f����4%�H��S~u�~���ve���}o��=�Zu��箥#�l�<v=c�Y��-;�1�t��u��%zqKU~�g���>������6�
����A�|;GO�k��-}�1j ��/$�Hֵ����^�ρ�+�c�H؏�Y�� ;Gx��K��t�w��O��
��<���+_��kR}����M��n�#C�`��O�͸anH*�-�FDeб������[|�R��K�x|��	 �P�?c���ϗ���FH?z����y���Zw�����׬��GO?%ۀ)�M�����Y��#�f��4�1]6>U�>c�����?�X~6�F������v��G����h��j�w��<�t���8̿G�vF��;���>�1�d���ؚ����/� �7%�k>�]�`��-4?2�W"H>�FF�&�Tr`㼎hd��z��W���FIļ�G>�۬���6�`RV�ZI����^�����0�'��/\r]�o����gg�T�V�5!Yǜ2S8��'� x;�[��7���8U��5�"*Bkl�A� ��T���۟��6#���C&_w��-;}��;�n�ms�%OO�ݽ�م�c\�N��=��^J�n�I����p5վU�
Mx �� 1N�uSX��I�n.y�r���d��d�[��y��}{���Ȍb:�p|M9��?p.I�P�/��ґ�����j?�v��A4u�k��5��@�9����4Ȉ·�0���xЯ��EJk4�r��S�'�Bؘ�vۏ�w��+/o���wC1/�I��F����h�ر�ҽk(bt���;-��gI&/%oJ�����0`r�у�CU���@o}TU��b<E���P�	��>�:B/�)T\��״V���~"*x&���1D� MV��}����$n�0�0��rI�M���wJ��Џ�mA��r����`��BX��*��h۩�8���5Nު�n��aC�QM��?����Y�E�1D�/ow����6��_��5Y�TP��x��>[��$��6_3�|�& ��3%7R��h>z. Z2����[��%y��7Xk�X�(y�0;]$�/��ȴ�� y_f=܏�{ճh�/G��cM�����.v�˜˃<ZLxɑƊ�qQ�}��[���3�J����am�C &�m���v� )vYB
��Q�I��U���U�u����=�{��S%V�����CUd����D��u)!��w�1ۺ���4��/sN0=���Y�J��!5і�,� �̫�@u|N�X��G�d�_Î���Y����^pF�#�C7�S��O==Z�����A�M&���lw�YW��j��,W\�7�V�WC:T�����mY����ȡd�Um��خ�I�A�d_�����g�I��x�.I� ��'�9�	�6���ղ������q�R��cK�n�Rx�Ez�v�G6���~�_�2���Hl&����	�7/�nE�j��J����^u�ÆeR�d���+-QW
^e�����ꚪ��h4�z� ���t��D�dC��d�8��]��I�X���A����W��Y�|��3���	�f��F����x8O��=�iZ�7FʈK^Zgʏf4=��a�HI�c�Κ{���24�"��y3�Am��w(E1��Y9�S8�m�1�֗�
@�6�(K5���#���I�tP�7�	��-���% �q"�`$�'��a���2���%qoR&��p>ʪ���&{�E�=�CR׍,�m¯u>������Y��͠r��]a�ꋵ?�ap�|N1H�5�Q_�P�|%^�a��E�.W��H*]^Zd�.:o@�����ǡ�W��z`Nqg��Ԧ�RDic�(Q�S$��@|a6[�d�`FB�ށ�q1��7�Q-R�Rߟ��7�;�KM���GhtɈ�g�ՁbC:Ss�ِ0u�Ru�����h��k4S묂2O�XȒXQ��>#W+��%��ߌK	Τ��˭�A!gV�o~j��Iv�[p�`$���{}��i�#?�Q���~/���Uf��@����\ �е����tk+�O���
n�,7g��Ȏ��Y#�X��Y�E�y�t���,�`ݴ��lL���{Ǵ	��qS�u��t �Ы��'`��S�-w]��h��
B*~��uIs��b�-��JZN�ys��3��(MHƠ˪F&�7��$ ��kc�+�6^N��>b���c���?q�c�o�P���Q��Q58+�4�̬Y`�t�j�߂�;-D:�QU>��*��҇�M0�?�<W�Ű�C�8��-�!�NOv�ʘS�t�v���.��I½o^��8�h8��g�k4����Fɾ��f��!&%�ʑx/���Ѧ�2ҭ�������I^�~�fV�wW�Im#�� ��\�wa�jR�#����<��^�ә������4u���G��t'o�U�&��l�ӵj��\�d����Y�V�s���կ�]�	��w�%��cJw �1p+�����+	h��𵜹w�/z��0Tap����$��7/WD����+��#{�s!��V�>d�v[Ҥ�Na�dWR4Nx����h8��5e"u������M`9f��������Z7�W��b�4����N���|��;,��3��$�-�Ƀ�yoAs�4�}��99�y����i��+����F;�m��9
>��}j��:@�|��={-��Qx���5T'��V�E�3��5��{껚�k��/��LC	�����y0'�����2��~�H7�S��=�vg�������{l�d�70��z�d���jfΞ޲���(��h����kM�<��<����Aw�k�I�XG/��q�Ǽ����g�1BF�� 	����ә;"s��8B6����6��a��`�I������?�>���M������I:��t��)'x�`MOޔ�lyi��Fy�l$Ʃ�a�`��#�B���hր?�ʿA�F�1!���-�|��r`Z�X0Ղ�b��Xr���&@�j��I�����N�
vw�����]�N���ˈ������()�e��^�D	P
�zXv�R���[i)�^
� �/QjW^7}�*牞�R�?�
�!�A�0�Y>���J�
GI�е{��t$V�ptG�}���K���b��J���o[��v��?�3�1I���^�/6׌�^1��Z�="|��?��&T��8�6�>��������₤$�$���},ЃQjt�r�>� z	���g	��������X����n��ӌm�5���aw4g!G<z��4�iR���f���o�N�_��M��v=��"
;���ӵ�Oa���i�B����<Z�I$׌�\3��ό*��؍pR����4s�p`��$>��%X�gPؔ����D�����psY�4�SS`��ֽD�;��cѮ�e^���_#�Wz�Hf*�<��ZR�:�s�0n����t&#����)�F{�kL���v�l΋n�\��/���>K S������;a������ם�(�Dl��8�B�g���ϡ_kAt ;�[� K���ˁ�f�~
S��GXǣ��J�A��s��*'OR�4���+`�r�¬U�aK�^M�5!3����ztʫ�f�[$�D�\+b	���]^P=v������V���n�ݳ+���0e�.$���Ʊ�$�HR��<�,@�HI�$w��U�٦��>ۅ:l�8����j�E�p��ܔ��V��)�}��l셥?��k�_������VS��
�Ʌ�q�7� hQ�#�'�)�IQqa�r�{��OG�b��ڱ.	��ό�D���������@h�H�h�oҞ�R�s=-jI�^P˲�K�D�T5m���*)5֮�7��7��^������?Y�s�ĩ����&��Mѳnm q���q�T�$@�
�t@��hU��v�/5�XEx�ϴd�%��o6X'Js�H�s���h��l|��b���1o�=��n�i�HZ��^~#ަ-��� �'g�#�����o(r	b�!��d�)�f����1��x,r�$]%��hY1���GS���Ͱ�#e��>���o6ʊᇡ��A
d
�����O���uz	�&F�:��ѵ�!N�xt�� ���v�Yd��9`�1��Ê�q��M߉��T5Dv�\�mu늁2v��OlCpN��k�C�����,����'�W�t�����0{���/^~�^{5Ch��\Oq��)U"�ZY��>)Y��{��z�X5�JH���v_MD�;��F�0�O��b�<�@���������<X���I)
�\�l�F�>M�<Awg'ִ�Κ�"�{D�E�wx�=�s��>Ǌ=�m'��uR@~�s|-�ƹHh�|ֽ�(f�;h���:8�����F�D��������2]��o���NX�=�8L�h�� �,7T�<0��@�,�b�C��fn'��ha�� ����ו�4�x����Z��װ6)N0�� �[[J���]���W�1Nc�[����������0����0�́�10�&~��!n	�4
. �m�!�26���?������h��^�]����\��Ip����KvB��s�c��.�������C�L�6S�f"a����n��&0O�)`��k�/���lpa���2Z֏�e�HcV�M��40H�	�H	b�w��9����6'7>D�11���^���m$�����Z�d���?rM*a��щ?88�CO'Ud�LqX����`6�13�N��G�{�.>�b��.l;�D�|��KI���3�-#p�����[��)I��3�D�Km����A�N㟬���?w��'��O�z�%��]�M�~r+�2�l���uO�m蹷�1C.؝`4��:6#*��_XR3���u�[9�����ϲ��4˜�{�A ��0/.�|���5�,(�]��ldF���m�ƍ��.��Um�UE/]�5�"�lkS#�r:���T �tƮ�*5�e������؎{���1w.�I\���:��kH��2;�ͬcSF�6C�QE5E�0_�6:���Cm���6W��h�@�@ל�&�w$Ct�$��z�X�X�K y����xÐڙ���]�=׿�&��?���71�,7�.ˏ+@�c�
Qq?aI��$oB��I�<;�#��u��G �����d�?�����/�9��dd��k��W^���"������^M�<��Ut�Zzّ1�}
~�s�N0�t5��L�CP���o�&�J�����%
����qu$^��CD�m�yps}���U��+�yݘ����Q��֭����w��r1����8�&O+�'J<��_�8 1.��h�%eA�E�l��5ﻺY$hǌr�B0@�	~�p<���.�mG��C�j�!�DD޹�FR���((@�_S1�2�c������y��r��K�6A���,�_H�{͝%p��E̱ �;���(M�G"s���1��I��d[���*�l�'Qg
[T�!�y�~�[rB�Y��YP��#�Nw�;0j"d�G`U�ݴ��JK{�.��$}9�8*@�D�vr�w�.�]=�^A�~3���9�<B�vGU=��Z��O_[�b��!~O�m�F����ŕ~M] �2$#
S޳��1�t��0=�K��j�6!��T�IH��tlοB1D�����u ���c#5��v�t�ċEo1��aq��]����&���#�m�Z���Kg��	SR�{�1ꥳ]���48���*�Ǹ�iO��)������Zz��2r9��Ψ7��I��4��l��W0fzV�j�Vl��	��������-��3�}��aw4��M���>6�s.�s?��8Ue0��_�2J��G����ć-�$�A��C���oOJ c��C��u����!�~~��������t"R��4GI�j�x!H���vs`���õ(�<W\t26>��U��O����Ƅ��B]c/�s6���_�9}sgj��u�Ql\~���vd��NR�u�\��1nAb��Nz���2"Xg�K,�D�PsD�%w<P\1�OM�m�=���|���ͫDo�N2E���Gl�U�����'iS��hy��|���C�nM�M��O/��V`���;�p��ʂ��A��2p.'�Q�Ī�k��Ue'Ͻo���Vd��e�~>g{�;�@h(p6�HxvN�S�.�-�ȼ�@�L@�x\��?�:�)^�ׂ)�V6�6j����=U�Y��xw�6��V9��>4�lS�2��+ڈ�#ϮmR�P��W��M#9�+(X��������9Ua���-*����?�ߓ�%��18c�
�$C�r�9��`:�tl��g��:!Ȳ|Qk�t��ԢU��L>*�/Ei��Μv��&.4k3Q��i%�-�C�p�d��-��֦}��[FE�S@���T�g��9�0!����'��_^���	RE���%��>2%!f��~��P�㒴{�	ʰ��ɢ�Ӗ��=w����KSU7?�*�:�%�Ȇy1f�Q�ud�ik�n��E�������ׂl�����(z\p�PF�6��N�l{!9���IN�R�Jww:�?������U�#�p�j'�����$�J=gG�t[,�Jm4)�8�g�|�uS�a=� �[V�y�)p kxk |f��&���4�*ч̽��.�$>�
�v{�=E��!e�O)©$%��j�S5�\�w,�����O�<�9m��d��7K�yO�K��ȁ�Dޠ0 ����Ƴ&Y�B64ՙ=�"�
�q�"Ə&��o/Q��<�'��NZ���RE|/�F$��'��W65pOU/H�=��nj���;�?�H�b0����z9X=�\Hޒ����ʪ��Y�S�*x�p}$9�@:i��?g��T_�vj��{be�mAu�Ç�I-�?���k��}�#����j���7�M���$��t6��gh��}*��I;[+O,��a���'�|��b���Uc�՜N���̓x�����s�T$��?UP��v_g�rrF��-)���h���6�~��hI\��ɷV�hc�[��N6�:R�6a��ܑ ��X��0B�~H�8�[�vrV:ńd���,�\��Z��wshJT��3ێ���\r���C?f_?K@��[� �R�)�ԥ�n�mx.�/2�\h�W���G��T�(��NG8����D�~D45o��w[;��������T6��f�Q{�D�����).k�E����O�9���2�R��&�!��,��B�HP7�����]rV(�5��hٹdm1�\(�|��(#<*�+o��R�C�eZ�����,9�X���~���^"P��!>%����b��v"&)���K����+�++Qv۟�-�J��6�9#��\}�M��iҕhJ
�����ئ��>Ӣ�@ԙE:7N�'�Mﻐ���ϋ���r��ɿ8���1~Zn>����je8Թ\Bk&�S�����y���1���F�NU�d⽡��S%��yV���
�P��Q�y�98D��U>]4ק��1�Z^��AL�� z�-��47����ԉ)~�Xn�4	����8���L��5�I<���8�/�n����x���cs������#��F�d�@`d�W;�E"OmlC ��q���|���k��oa�N�C�J�����~Ե���@н"���<��z#>4$¼�s�tǂǟ��ޱY��O�%uY�t�-�@��!�юjJ�M�G����C^�^��2�����~�WIw�DJ��bH0�7%b���؆��CN&0�x%߭4Xe7 ���Gt������$Yw��p2皂��es�kP�K_&��9�A>CFNӓ�R䫆��z@��n8�׾D�Ry����{6�Yf��P���I��������\M0cԗ��<!+��	����\�ّ�Fkt����;5sƎc��ǟHT�U��[�XA3�Y�v,Q�A���#��P�m���zQ�W�s1�E��s��g��L@	O��V������(K۔���@�"��*oYH�[=
=DZ��)p���5��T_ė�H\�*�Āt�jt�y`B��/�<�u���&}���{�]��ɸm�t�/���gl�W����w�/fVe�m �z8�`Ʈ�)�S��UBt�PgUP>�źD���oT�jV����C]��`�q��b��E@��vP=З�ח����]fU=D�^��1��ً!	��%�2PQ��8"g��s�������T�x�R���*{�p5�e�b��P^��0�!�}1;MT��h��v�L���NM�o�lW��oLE�����)��bԴ�ݖ�eb/S���{:s$Q��c�r�[k'��!hԮ���lo-�^aQ�[6+���h
8���Lv8tm���vKLo+��"L.�T������^��ƌ�M�Ǭq4��*���`1�6��:m(�������Ҵ���+����K�q�ӕ'�6�E/8��V��ˊ-8�!�66�'m��;��u��&�f�H��O��K(�z��b>N�3�%���ޱ4�����F�f`�j�,d��5-�6\�B��s��r����E�y��5�`�t����o��߾#��M/�f�Il�L?e��u=@����q���H��s�>��s�'ܷ��]O�Y}�L����dAx����
[�d��7��(*92O���e��� �A��*q��d��4����l��ä��C��v'�@��F��k����ܼ� ~�'�B�����H�_w���¾ILM�jH'|n��&ո�G$�L���@�:��1�G� Xm
�;t|��#N��{t��p���V��D�d��b>� �� ������h̉M�,��	6�$�Z5*(d�vNf�D��c9%�$]]`�Λn��!��Ẅ́n�O��mkki����W[���o�ڳ@������@VH�]
���F'��	2��!<�l.h
�LZ_�oSH��N��O������&1���2�hg�a���ILP����A����>7I���r��zt;�%��W���Z��Q���~������\U_���1.�d5�[�����Zj�tE���XNI//šܓ%��{5���s���� �[�Ц%�DZE˰����qI���(?A@0���d���x�v��g�T֣�}9��?௏�,[9S�!�۵�����FF�ۚR�3�5E����(9�su���\ՅV��Oѻژܺ�=SQ�ė���c�pz��4*BZ
B�L[�h�Ծ ����,�	k��4���3Ȏo�:b�W�F`�WA�Q�?6����ܵkM���]���Xw�ո���n��|�Z	_t�21L�*B+̟��)6;�5B�k��Ko���3VC�g҉g)ݎ�pN�$ɀ$V-���H RXE�i����,��1σ�tT!������pn	^lX@/t?-����(��AI#<z4���*�G;�-���2���	ny�m��!e�B!�� � uO��JX��Jڗqm�xp�#�ȓM�/��#Y^�a��q"	5�]�L�qٙ#w�1ϐjI+n4����7��]�;K`F�UQ8�ı=�fť����g�3�i���,�3�� -K~�k�F�H�� ��4YV�Ҿ����w��/����W	\G�˩d���ye���zG�Vؑ����t�liӖҖo�8k��<�Y9@լ�̭W��=ɐ�QY�r�Ul�.���� $:�ڊe�6�Xkg�E
E*%�e�-�J�Im9�3{�m�*1�r��o���"�6�9s��n����� �ot}� m����-h�bM���Z��_����R������\���EZ^կ��x��U�g͵�͠��#sŋP1��N�����7ݙ�R<9e���(�����=��'9-�푢�Ien�ƹ��ƈ�=b8R_�z�ĥ�cY������ű=���S���QH���5Y�V��my\�e��&,y�3�:�Ǡ�ǩ4���fު�^��� 4?�����Y��%��e?�����[*ȠK���>b���a��Ӎ����-R������S1�0�?{�z�[�oEg!����Cg�l3K��!o��g��*�賕�Tg�ҕC�5�U[Hǡ�1*)��Ɍ��$��������w��T�67� �)��(�Ri.��\Nh�6��-��<���N	���#����59shD�Q�V�U;gM��5'#^
�&f 1m62��ۙ�%��P{}��*���ۏs7$�|�d�������2�s�|DN,�'�Y��l�J�uz�myz�274�VӦ@�Е�Bm�	�(T��2�B!��dJ�\h4vfl�i� 6�g��/q���N����b]w������b�V�v��A�L�'ة��+"��猡'n9L��R*$���9r�i�\|b�B�pm�Ƴ���V'�g+�̺�e��G�n��;]���؜���1����G��|��+3������ە^KT���,"���=�p��.Ȳ���K�,����v����ݼ����^�Xز
����4D�@�j��g��� s�B9U�G�Z%��K�c�#����t}
�k�HcN��B�[k�U�I�P�� ��.a�����ʸ��k�њ����I8x���(����@��V^٠��1�#���o� A��ѕݘ�M�tz;+�s�m��,��TQ��T���U�IR�������}D����74�7U
be�ˀs9H<�B{tE��C�Z&�닁��2X!=���%9�#�eF��K��V���q�l��V�E~a)�Tھ�A��T�#N��	2��P4��G�]�|F뗰�v38���S���sƉ+&�}�h~62���jŃ�W���������(�y��y%Z0�X������b'���\��V0�;�uo�o� ���O����E��ø�8Y�/��>/�����O"��?}B�`�3���l��H��~�?�U�����:�x��J�&�V���A1�V�dR~疹`Y<��IU�d�R���l[���r�C��}f�$d󊔩[$�a��y�G��8� ]�3V7$s�"�dH�������K�B��0��F&���x��[y
�U�=5�Ê�eh�x)^m~�[#;S��U
+� ��Rz�K X�f�le!���JQ��hg\�`]�hh�\�m�Ek��$����l���=�b������Tn+��J��l��*R
�H-�k�6T�"杄��S�����QS�;�We2(�52E�Ip�0BϜ�)���mi"�)�����M1�%S�����f_�K���C��a��\~3�5�n漲��+/�a!�>Kш��Sf�<�.M�P��5��71w�*R��{ �Ry���%�D]�KDߏ���1t��?�h�N#ߊ)-�o�4�s�q/f;�g������(�;zNl�k���Z�ݯ�/��d�nmy�PT�����{�����`��@�rmV��񵣖2�0�/n�3����s}^�Q!la���q�#�G���	GB��Kc'uon6��⃎����^�L2��?�͚c:��b=B^�I!'=���Y��6�=�G?˰JEe)��=��H�������t\�ZmR������"�f�;p���i5�D�*0>����ѻ�JH2�7�A� ��M�������Ayw�p	��M�UϮ�"�}��\��@�ñ�bة�XM�CT���BP���@�����J��vp:�]"O�~Fj��(H�<^�@����Q�Y��-���#�9i�ôa�Op��k�S����ϛ4��"r�|���!�r�y4��P��Q:S���J4�%�T�f<׭H!J�n�4W'�U�V��@�p���IY'�l�`W�C��^�Nj�@���q���q\�w�̻�����3��\'���꧊{>	�xM��u��Ld��k������R-�g��D�D��N|6���ƺ{I�No0��eJ��w]��,H�-��M;�\|2N�����ax�e�sy>D<�:�%�;̶0���t�^������h��~l_PH�� 7�~ѥf�h��Й����ao���t�#���c�vǊ��R @�DKT/����XdK��e�&&:���S��[\Q<�k��|�鐢`_ި����G�gѸ��{�k&����6O�v&S���W�\�n���Z?�y~V2e�M��֬��uݠ��iI��>�`�4D@]|9N���$��T<�$����j�POFc,+R��V���P���Ir�������A�&�@������E͏�r �8k5�I_��=ns2�?moŲ�;�Wv��������)f��@d�gclr)�c�M�i��!�Z��p$-g���Y�)t�q�{�R#��a~������C��?2�<k�2Y1�=6D�mUh���,���	��Q�6�L�D�\=Lȵ�2�<��M,���p�Q'󾭟-�O�J������2��R�0��h�$����Đ��`���h��V����P�Pz����{W����1����[�Ћ��b�y�7��ǒ���Ǵ�����U^^PT�73��H�@^��������$�r�gg?���#�P��l4,�LZ��*�Oh�C�h�Kb=����r��ۭ]a�/�.S~����جgVn�n3����@�r~�?�6`9��(��vO������U�W^�����(���;�M�&�'��u�3�1>+���.�Av���
��[~F����9��Мc�kZ6&�4Q2��?n�ӄʣGDD/���ʋ�;��f|��woG�4y�D׉��!M�����$f������e�Q���q��H%z��� A!'���D�j��Sel>�0ʺ!�N��� Cj��b��7�
��p�fϱ��AT}��^?+g�($�T2z/u�����v�c�S-�����R�-I�;
h�$��S�܁��#��u(���j\77�C�X�K��_�Y�E瓖�7�Il�)���6��a��h���y\���}�#��^8�4��)'�wv�����d^��W���;T�i�|������)J)�5dZ�Y�i!��c����t�ʖ��������}u;3�˻��uIp^:�fP���ڤ�������<������?�
���ye9�x0�:@�$�l�B�=x�z��|4k��k[FBJZI -�)�Y�$sn��k��)	�iYaKZ�)iq:	�<}�x�)�޼��������;�W&5f�.�c�!��K����
 ��5��d��
,��<�X�t��a������ʰ�L�������M�޸��5N�n�|D�[�@B{d�|"�+MH@���� &0��*O/�Y�N����Y��o� �;8`��f��p}G��~%���ړ�\���,`Ơ��=U��s�OQ��G��W�y����l 6�~MX�A_�8�sQ�)�_��gB�3��[nL���
ȅ�&1�.	m\`ӸT�C�a&~��ZlA�4&�̈́�C�b��I&�˾F�N���2��������N��N}�1��-��Up��4\t��i!�m��l�/g��`�v�_���`��<���e������o�V�LL6!bE���Ѝ���H(�n��=��2]wm �%-�n���t�b/Y5�&_�H�0�����~B@i���}��h��#^����p��v��DQq�zݟ

�f�d�,C�Y�ٓ��X>R��-1�"v�=A��&����	Dp�|>�tXX�h��dv��z�z�q�^h�1�'�z��z�CV�E�/�:Y�
2]��}��G��$}<s?�(�/_֊`�P$��9�υ	3q=(y�,������iK[-d������w��aq>`>���#�j�=͇��	�t
0v�F�� ���N/G;a���[�j���,��g?�.�����n�|����r\�rR�S�� ab	�b�Y�v;�x<4'�t�a�*]��1�k�c(�S���t�C8ߗ>/���r�6U`�r������(���#��{1QE�6��hF�g�@2i��UM�Mt��N,���́���+R��e��G�0|;�~��7�IVc����17]�	#0�,���6��풲��l�}ՠ��%�����58�h:�n.:p�kJ��ߔ�Y����>B��6�nX˛��s�7�E
�%��]u��ᰞ�Cw�1�E�fDz�����3@�zi'o�U{�7p�E5��=���Ab*Ƌ̜?|c\睓p�ȸ�`�ȳ�r������REs�%�	_�ҽ�b�wn w��I��h��%��҆
�Guz'�k%$ɜL,,z� �(	��9u �u]��;����uM��E,���ښ]2��0H��g ٸ+�$5���Q�[SS�=^q5�(t̢~�CM��2z�9.���K��,��p�b(���1��/�F�Px���K�;I�J���A�܇���:2�Z�4E���?�{�9�}�g�: +dls����.����Z{�Z�*ԃА�&�n�!�v2n�aXU�7��pcG8���G�!��q b���~έ�Q#˛�����+2�����,�p;f��oEs��ڱ�\w���Bn��w�:#R-��oJi}�j���ȿ3h���$&�8��R��s�V�H7?������F_	��:��j	��9�it+��2HV}`e賵��WL(߻��t�N�)؅�7���Ζ'?��a60G6��a��|\l�Z��;��n�ȴ��ڍ�|��ח�{�������n"ӵ������:a��?;�\j�J�/vY�;{k�+�'׹/XЎ�3����E1��Ps��͜c�x�,1yzq.w/��23w��>V����V~.����q}8ATn��׋:�9�OUO�=d��K�'�UM�A�=�N�Ǎ�^�lV4�z��͊+~Cl4����;�+�vB]��cUɰ�����t>��	XeJ���fY��خ8�<����G���S[1�i44��Q�+�{���K@�����B���CD^@˂�C�Hi�uz�_Qa���U�]枺�~���_��u~gb�]��wV} �V)�ȳ�1��h߮V��յ֨[���7o�+��h�4�4]��v��$فl���Db5U`��P[|P���<��sRW5�m̡�Y�Ъ��z�4|�*�ж������cw��d���Rt���c/�h���(i��Oej+4t�5݊=E]���+���û[��m&��7�d�PJ�^f�{4����k�n L>	՗\����=<��mD691'��Ij
�*<�Q�z���4���M �H�$
(�=��U�Q�"�K&�$2<��Z�5,�@�kEF�_Ē�3ev���!��;D]Ȋk����;A ^������Nýk�������%�F����]/�_|�s�ƃ��iK2�IQ����{`|9�\��F�`2�(��]%� 5�x��2W��\\~ߜ[|�2E���eε']�h���s.~���C�c�<R�N�̈́DX��Ʉŀ�Ŋ-+:8���
���_0h��FY�3uN	���2���6��$B �6W���Fd�x~ؼ�D��굀iH�e����d�;�csE� )
�+yv����A�
MC[<ҜI&�#�Қ�xd�jO�X �/	���(ST�򐯍��6V�iyбΓSo���q�Q]���"����m�>a���d�E;k���|��!�,��U(�f�:a��%2�9YM��qT�r8ac6��������X�8�T斋�we�֓V:-��j ���?b�|L�P9�8.�U�����9�H�_`I6�l��%:�-
����m��|��`������\�$o�X�CRu���ȹ��3"��;��ax�A�6��= �����*�� 0�R6pY��-�∅R�]�bŧe���L�1Њ̚U�?1���Y� d�
p���m�G�y�1똎��{'�&�2䥭U�76��֕�i�T'H����h�q���u�R�OR�%��Y[��Ѯ��6M�y!w{yx�������f|����B�JI�İ���]ц)�r3����z�F	b��4��@��|�G:���?(�`��j�E-������D݅B��F�������՚,8�+�f�w�J�
�`�DS�����.��V��2���S]���<�5�Dڿ|x�� �(����UѾ�~1X��;O����i3���"j	���BL4�����l�E��}ȁ]�j����[Yh�$R�[��25����Cm���"�0޵�\]�ώ	�������&���.�0�&0C�7���>	�DO��`>n��s�8%{3�����0�����_�؃*����Ƅ������p�ޙ��*��D`
�������yM�_?��Am�;���<{ -7>{],m��������*0����t����k䚴h2^���0Q\Mp����:�Q�g���dl��֩#Cb�j`��|�}\-Q�e����`�fL�>9��Ӌ�I���5�����;g xI�SE�cTE�ɍ�ם�Ȉ�Z��J��9�H�����c6T��CKpy&�퓊pQ�^�*rb��O���&Ѽ~��#^��^YM����}�L'�v���Y0Q�����t_�g�A�pcxY�-8�U�����b	/�!��H�n��ſ3`��Bc�Ubڇ���JtF�C��of�[���T���]ks3��V�ϙ2t�����`��KhOּ����Ѝ��c�%����w��<�L0Z�О
O�~���q�8A�\��9�������
�m��8��ss��\������v�kL����c�ǁ:�Jt���i�ⷂdZ��������7�8�:7x���$����'���_r�!sIe�iq�̜�:3_O�	v� �D?���� �O�ژ��I�[�A��V�$�K�b�3��A��#�h^� ��)E^�R�hHŗ�h�9R-f!���V��`cX4qxc\Xk�VQ��D '��g��&&-t��9�H�ΨT��	�k��5w������
gU�F[�_oF�;�⮰��;J-��`���w����ȇ�� _痤H�Xs��"�A�*W��9�+$z���E�U�@k<�S'g��PH�t}	���E�p~�͹!q��PM_9]�WE"�Az�?�7�b�Z��oQ'r����ʨn�L�H��~!�u����@�JL���~�[��"����������"���Pr	������L{�ٖ��.���|P��v�Eo�a�N�V�K��/)���|���/z��	ӥu;��%��:�O��T��揯� �
�)!��uS1O]�̓�.d�K�%�ޯ�.>�T�!y����/jE���i�Cμ 'L싂�G±�$�����wN>��m��2+�#�N�5�2���QW�*L�S��:����o��0��-��D�%��G�jV/(f�m�*W]/�}��~���fDE��z��}j�8P?!G��$Q��?�Ak��t^qw�x(���"#�TWb��˫���P�7}Sg\�pI� >��kץ>YKoi" ���%�]/l�P.��=2��-ԚF� y��>���m�
��CFA�+�o	~�°�t�p� �r��=Jv_���	�w�Z�-f��IR����ȑC�d~�#�&9<���h.K���KB���꭪!24��Ad>��ig�{kTtx���5'�c?]�,?�ѵ�k����4n㟗f�P�q>�Ǟ�/�Ĭ���N��!�u�5�Bk}.^�����0��2���I81�?%�[��m!��c��1���!��K���0��5�[	Z�����|����u'��%n,�z-�Ќ�rޣ��d�5�W|?6ma�[��q�/��b8}o�|�aZ�{)�W)�%"�es;>���
�k����5&���s�R⚠Ͼi�Ut�dR�uu�"�5<(QbJ��g���pj�(q1�|�̪,�7M)���G�j�>�d���j$~������|�eVmIpi9�:uy����{�mسu��%�(����Kv��|)�)Ny�%6j��|O���<��*�g�����oP�o|�3s�2�Jj4�cVEK|
���r����=�����6Q'3G�s���e�$�!R0�y�jA;mwok���S��;k|�zGZ|Ψ)�fRP��#�GlIwe_D���u�O�#�;#��ڈ���A��GfK���&�0���e@�ޢ��Gv|�y��c�����q�E��7����3�_�ݠF�~�")qe(s[?(�U��7���ÊjM��b�ӱ�I�%TUJ\$�i+2P�˽�(�bl8�� ����	}[!�'r���^���~zf�%I�I1�d����+_hG��O) ��D���
U��Jɐ8��
��5<�Q]ݥ��w�q&9O��wx�T�&���Fۘ|���]PS���<�]�Z��ā\� �ɀ��#mO����<����0��-�~6�<VZ�,K��3�h�쳂�$�|qyL�iQ@
�ZuM���Gؗ:��ѳaS����� �p*������i�R!�|G<�^XJK�^�<;f��P�i8J���uHL��\�릊�D �^�-��r8r^m|�}�����X����K`k��r�S_x[�
��;l�p�ׂ�D�uqEiX
U�k-�M<˸��	�h�,�/�)H��qVq|���H-x�,x"���7��ʬYl��d^Ey�G+�r�xfdg"�R�jD�"3�>�E�q�s"��ﶰ/K���w`=vss	"�\Nd���x�$��0u\�0��������)$��ɦ$b
���ËA���a�����w��s�I�ѡ��R���[8���~��;�>�6m���̵+���(t�_��^�Id��W�E���j��,�u�8/�[Cs�b;�dY���H(���"���:���Ya�4T���clQ��<���^_��1-���=����Pk�M��� �%��4�-����d�.ǄPA0��5���T�l�ho*��ip�e)傅"�>��uc�������*� t.�t��#��mF(,C�ck��Qơ�'�Գ�/�D����Mt�v��y�b=|e��+��v����:�'�k�_v^�_��:\Ќb���%Na��x�J��2"�'b<z�0��I���F݇��4؛P�
aR?0ʒ��� ����u|6�ߋx	l��U�¶�ߍB)9��Q������+u�s_�ɢ?�T��w�������K��ٙ�b���QeD����F�����ܿ}���|�+��Ǔ]8�N=Kf[�<v��K��d��θS�.n��bi)�I���P��`�j��5�y� ��V��݇vH�G؜�˼!E{��Mq]BTa��}Cbi������1IH�}����b�^�q�}E���j�rOpw3��!;v�e��H�Vc����nM�?7l"�I��Hf3Cރ`��7���z�)c4�T��9��b��44xY�(����,2�k����|VD��$?t9C��P�̈$�EO�O�ۭ&�0�|%�%��L�!�T�-�yjDׅ�����b�%
(�(�r6"��1;9/N:�>�)Cgc�\V��b<�&���B��C��}�̛�qw�<���Jr2�0ઋz��>/2뮷Q�9[��^֋@d��[��v��'��H�X7W�/\�rz	ڹ����e�&Y0��g��eJmG�����er��,p9U5��޳+b{G+��P�9T�b��ݼ�ki4�O&�,�.���Xd7�+a����4��Me��c},�:�Z9k[����W�v�7n,��c��Wwj�NE��+xUF^�0A,������p��̪������4q�A�m�s�=���	(Mv��'~��Q*jfK�vt�%��!%�.xr�T��1|&�e
���K�)/�����}I_�f�M~g�b�����*\�&�����y²�� S����M(b� �*k�A�M
}�����W�9ɕ��!<*�Ě����ț!�f�MҢ1�S���1��?F�$��k����ot%���﯉.j|�x��������y�<ZrqFT�0Lr�ô=�Vl�Q��&V����y}e�QE�ĥ'� wQ�'[%��[0���0w�����id��s{���~5���+-;Y�"����u�D�̐����,���MZ��D�PU�*��k�=��P˘ ���M��9W�9%�Oc7��l�]W24{�. .\����z�./L�p���&?�{���N�������pk������L%tSd�+5呺��*r�]�.hSG�2�:hT*�6q*M6#ü�nu�vU�kpD{E���EOm�V�\���3�����~�o/�Ap�
�6� ���K6��@l���ܻYq���D`((�D��p2;u����h.�_i��&���d�nA5��璹2f�K	�"d�s��Q����� �	�X�ƣ���hqN�໱��9wMi#��7+k �Hq��R�C! l��`������r�[���*x��D(�� 	��dz��\�#�/�@�W���gD*��X�������
�A�Bl����D�����_T	���	S��<4��1�jLMZ�$s�N$��*�!_�_�G_W�]d[&8^�>�����j� 0ݹ�OQ��U�K>��aί!w�#Fi�p"ϫ���(�d�!iWpM���w�Xn}A��$O]���*��V��k't�m.���V����B�i���R"n���7a�l���&�(��\'ތ	|����(���K�(WИ�]Jxt�VK>H�7T��Z����������p�
�x2�[p�7�;�hJ�{���;"�K���!mC8��x���� �1�{����n1���U{u��M���az�|r漑�5qX��&��E5R�S����9E�?�ZUT�P�4�a^�yD;�{F��Ց�`����Y"��.ߗA=g0j�����o�����mbf&�h��Ҕ-��Z��k/B�/� �ǰh���+eDj`���f�$>oE���:%���|Q�����.��M�}��YF��D��H�|�����Ӛ'ߊ���~<~s3:c��Y��zY��(D�7ǩ�b+ �r��S�y:y̔�X���5垤��6������i�q,�m3� j�h8}�%�����%�p�x�j���@:����)��*�j��3�ţi�N0u�f��x�S{j��ꈽ"�x�@$�?�H_&d�CK-�5p�Y�vzu�?�)��ޠ�ch�'ԁ�o��rlϭ�]�i��] "O����w�6�R�-A*�%p�� M�qd����V�V9�0��Su�]�G���p%��yH��65�3�>P�ܘ½��>�� ?���@%�W��T]�P�X���?��V(6E��}ΞĘ��~!�����uBK�֋���&�duƆG��ZC\��D��.�0iʆ��8ڣ���ݻ�t�{�,@���@G몹���Q��^;���q+���a�!�!�����C�6F�ns�j���/�Іoҽ�0<y����fCG�M�$�G�,�ś�HD>����r��K�g��nE{�)�,��%�5*��wx�=a0$+<�[�휖h�����q��Zh@	��?o�`O�e	s��8�D��J�_�(��6���p5��&�/x �^1&��'@��X�Z��FKUoC1� ����Z�#0ȑP�ѿ;��X�-�.[b.��݅�Q�g ��h~=��U��6e:pڅ�Y(�:PNh��CF�t9��~�� �z}x��Bp�r��zHU�a�V��$�a�oe�GUO�n.m�!.7�X5;��ދ��k�+��"����X�i��<��=���SD����)f-����]#Ѝ�´p>mk<�o�T�;��|�d*�(�����3Kp~��׺���-W�#��h�y,
�(M��ٍ����u!,[�\�̺�B�yL��H��\{IS�b�%�)z�O��}����v6��}}C�܉��n���q$+V��U��>K`��k0z4���=��@~;h�RO�)���q����F���ã����� ��Ɂ�<�����U���ա|�����L"�䞬��]��Cv.�8:�\&I����%�rSL�H��íB�E#�@P:��p
�D����khc��a�<����>�����x�Y���ޔ�q9����q��8��0yK޺Q��芑%���?M|r�T�� $fڬ&����,�����<U���(�:J6�'P߬5C|��1�v�z�ϛ-�Cԭh2�K���Ɗ�/��M��~B4��u�k�{��l%7��~B"mfNK����|0��q��ܳ{�ڱ������C�}�j�����j>� �=ƥ}��:�ߎ�"]]YsΣ=�_!U*I�X)��D'`t��~�#;{��^^��/�4����+��?XO���>M� ��bzt4��^��3��P�F��_a��Uv �x���a�l�PK���P߳�?���n����y�S�\Jr��L�=�HI ��� �]3�ЅL�?�h¾c���ld�J�Os[��=޾~�������G���9��o�9)�畜�z��9FyI�	@b^{��1��r<ZK�W'�é��kl�y��"d�������h��r��c�R��pa��? ��u���K 2�y��q�U��*Zʏ0�k�,x-��1��3�*�[9Əap���aoѡ���s����,��*|��jԝ\�� a_Ӂ�*{/�S��`�:u�N}r��ĉ�wz�6�Љ����!����`d>����?�O�DP���'�|���植$��'Z+��>C}�n>B��Q�	�t�3��-�Kh���r3	4�{��Zҥz��.�0���z�9�e�ʚ"I�f�Q��5��Ӂ^c%��V$W�/|����1`v{D�Sj"��#&�@*mL�S���9CvjB~6!��m��x�H��R�q�Y��Ѻ0:ln'�!�������`�����t�(F� ��g�h-H�T'�ƽ�ר����S8�H.�������ZJ�&%�'7����]��Fym�H1��Z݊�3���P\f=g���i�A��k,��!N\�ܕ���d��0�c���&��䗿X
�9�t<rZV�PXv�LXA�b���"�g��/�٪V���^��I�(&�^��(��c,�3�ܶ��������#�(�R���b��~sz
�$'��X���QG�fl\�b��ט��y�G*8<x��j�<���6;�$��S?z!Є�|G��:���e0���� �^�P�a_bR���Ed��\�q�䢉�n���q�)���
��.8Eh]$;d2ky�
���3!.@p���֨��
�:6��-�����\�܇��]��RHi/U͉�S�dS��H�#�b�%�Qehm�B:6l��}�(���(}G�>�+9�I�6��,�_���<�
śy�ɩ�+vbt���ܙY�3��[�{�ɪ��5k�K��O+Q�ʎ����J����@Go�驆I�c���8D�kw&���P'8��^�gnmr�愅@t�ۊ�0u����V�D0��/w�G�l,��UA\S#!��|�=u�������t_Cd+�CK(Gm��u�|ӓr.�dHP'���Ϧĕ������9�e� ���e@�������&���7-L��qQ�w�� \8��3�m��ay"���(�ꋭ<�'t.���%��O�~]���f9�Q�$�P���ZV��Ր��#��1�qUB�
vf��
��[7�h�����M	�zʸS>����IBB~����h�ԕV~�p~��̹$�9%1�]�y��1f^6�}�2Ǻ���d��oέ?0@.&>�!(�6$�~Y�l@�&��؁1��p�
���zR���I�N���6��ĳ�h`�̎�ms��e�@�����	����H�K�I�Ģ�b֜"�+����Z��_x_���p�ET���r��s�-֬$����_LQX�w؜FZ��"�AW�,�k��{`ےf����3�[R�ߓ�7�(S]J��#�r�{ IȢ>M0�'��ܵ��8�3�'�x͉%���r� ����!�pWo�b�������Ȑo�O!�BQ���E���ANg�Rg;ͦФP!/�c��nZ�ܐ��Њ��S+�(˴��j:l\S?�ք�#p��C��kQ��J]%G"���Y%s=���(�I�[%���P�[���ny����'/��GI�ә���I������:H/}`�s��iѓI�(��V�a��aA�	%�@OB�g
T��o�&�Pz�i����4(���|L����r0�r�~¨i��棪ZA=��Mfqh�"�Ae{�:�VoA}l_!�ѬKF���-�������W_�ե�<ҟ��,���Ez���.������,��2䏷�+ "��������U8��8?�>o�71�U�-G?�޳��YX4��!�Dj�E�b(,L_�+'ד2!Ҟ..u0���MKmDm%��`_���4�j��y��8 ��C���^���1���tt]�t��PcpX&!�[�v^�?��IU��E�*Q�Х#��Lʚ�2�n.R��P� �9��6C♱b��[���]\�k(��TI��+�RQl�3���#��h9�f��V�W�h��|��+��v���g6������:S漎�'pz曓$g�Q�!Qչ�9��?&��G�k8Z����L~�_I��|��O����Tsn�U4��7x�Ӻ��s��8r�i^GZ�̔��{	6���)�:�g�ε�Χ����aX��u�A�-��A=w��t8L'9��D�"�f�3��G��{"=��M�v�6T��*�2�KԜ1�#ev�a�9	_j��������K [3|��)�0�b(��[J�]����Ԏ/��7�\?V,��nV��&�;�&��E�j	G����}E�i�H�<j�Q���F�	f\����.�m��#	4�>*65����ݝ�]�݈�c՜\�9�7�ջ�^�P�`�\ea�mT���C.&fBL�$4{ڼA�%|����8G��[���4�3��°{��K���_������/{��ru_�I��.�������h	�;������Xr�i�c��3!���?هj�"��4���ۈfB`i�-Sm�t\�Uܪ��pܢ 1Y �ӵ��P.��:�?�Y\/g�����
���Y�D|,Z����U��5���t&L&��'O��~T�)^�Nd���6GZ2i�_y��Z��ï�c�˦��O���8&�4��q���T�C�и�(��	���r�f����u�o�z�\Sn;��d�^`V�n<]RT���%㣘�g�5��CE�7W���<��n��k��A�tD�Y�Jn˘�}Y���Lz�+������Q������#�������l�h\0G�`7�S���� orv��@_q��N���a	\�A���tmY2F�`�y2u�^��� =�����D�O�݂b84@ z��'Z�w��T8)1H�S�U�p�K$||��U�i�k�f�y$h=	=�!M!�qpz��'��fHM*w��4P�|����]T��X�m�m6g�&o�ܪ���� 1�W
�����)�Þ
>/�i���й����S�;�1N�P�Ɉ�?�OK�[�~�M!W@��/�ܽ4_X�q,M�  �2P��ɛ�M���cІ���.B�oca,]�h^Ǎ��㍄�x G�_j�27�N�Q�qP�����!PI��5[��R��HL;�f5��_�2U�6���bKA*�?.v}}C��D=,9BQv߃�0��N�R�@�ö�̸t\�&żVǴ��r�W�qiL�d�S��;|KXh��  ��cw�E��	@�����&���=k�jo���f9pʯ���}���GO$��|�C���̘{�S
:�r3i�4��$�� }��`C9[Z���D��ym<��)W}m+�w|һ;�{fx��&c-�."�~6+�aE��>�/Ehi�Ųv�!�9��w���  Z)I�8D�[>�A7� �FI�z��&�J	�mw�"}�盺��B(�� ����x\��3�>:N�G�w�ae$�^W��+�s��5�x&��^6���slDUi��sXP�Z��j%��9l�v%EUCv�F���4�&e8�J�O���<�q�\9��f�ͦ@}j�NQ�����y;�=�� ZOG��C��1mM�)&?��`qm������E�����S����
����G�����O#f�!�����H�@cj\�q�ޤ�SK��#��UUѐ6s	yJ����C:B�h����4+<o�y�J�$�v�� �Z�~{��݆�oƨ5w���KMO��Y#��(����d����n9%�JR�r��΅��n�Ic�_Q2T�Z�w4�'̥�j��?Sxm���N��	y�r #���?���~��/�@A�i?�>��an�VB~ڜ<�e-n)Nh�Z�;�٠yUQ�����q�#�4�{�Tj�� ��*�eȓз�W}�G�j��8�u�\�]�r�_S�Uv�����@׎ q��/r`�#��<�c��u�gN����2$ZcU��<�ȯ��i�S�+j�v�j�����o�Ui'�.���D'����m-��e��~�1����b�DQڞTƢ�Ĝ��@�dΰ�SY����k��/b�U{�Ϗ�S������JĵC0:���y�I�nM�e;�	�:YkQ-�:�"���:�SR��2�Z��֝E�I䄸�ճq�������k�$���ɟ[P?8+�������\N��o�ũ��饢[���"=^��S?���</����R���rk����"��H\�����l�Λo3�Hl���:ϔ���k.#�]���Y1\����ʏ\:o��:��Cq�$��?b��":��p��9J��91Jr%qT��^�\�;_��|�M!ZOk�<���(��Xl%����l_�T�ϓ�6�w1�f��]t����FS)EY/�]� �|J0��_�a��?�a!�.���%ަ�9?ʁrfhG�����Z:@Y�:!�c�4TX�w��v�k)b.щP�P$�s�[P*ǒ��˺�F�^�>�&�ւ�ӹ!B�>�m,G�/^BP�z�{�}f��������[���4��T7F>7�]��.VL2;`�[�����L�z'��o��Y-�{���j+�T�b4C[%�� 2A-�Q5�����ʙ��X���a�O��_r�.�y���/����Ժ�R�E�?z�K;�p���R}�lqko�:�|J�W�%��/V��O lOlͩ��WV� ;��%�^���܌�,�Z�`DA|�ZW� "A����pp9f75�f Q��/�/�>���L����;�7��Ԍ3~���a�dl�%}�,�,��=8�h>C�N�:��S�i�X�~c�	��֘��ve��U/�E���;c���ENe=���_3��w,I�YA�����]e�>^%�@��<�u���ɾ��^C�5j�3����S
���m�}I��D6T3YY��m���Ԣ@�����*���H�#a�TC��[��侀|���V�On��G��~����jЪ���h%�'KUR5�+2�S��
���2�.������w#�Ľ��
��Fӫ{�k�MK�q�V����#� ��oF9w��
�<7-�3Ĉ٭�&K�*�P��!@q��y1��������������l���y��	��߄Xjn�a��z�da�	��V>&]��~����#���[���/��?0.F1{����ZN��k:����P`)�:�{�ô�l��/ncFL����IGf��/���;4�-. Y��"1 �(�3� ȉ��A���s�k*qDɱxU+�� /��SJ�I�Kh��Gx�G&���j����4���J+4��Ak�xU��Җ���@<�����:��@9�d�N^qR��W����Y8���MF$�P1�@��䯺��Z����1�ͳ�|Mi�%�O�l�&��_brL# e����M�*�����ŷ;#���]���dݟ2/�(��Vz���ou�ԟѣ�4���"��'�)tg�-����G�%�W��uo�a�SÕ��a梪O0�o�e~���ĿX�|����Sc�aL do�ʁ��-��9�� �c�y�K�g�5��d.=ww!u����= R|�mGBD�o�:~�l��p#�2m�8��o揶��0��	n� De2$e4��.@ c����:7ID��P��4�`$�N�"�Cx�9�)>���<B�g	I{�on�+��F�$N��+�a K*ׄ�Df�� �!�Z�1i�1�S0�����Yױ�d?�T��p�N�r�M���LB�$h�D(���|�/��>c7'����|f
	�m�'㬖�ف.���)�s�����B0�^�$��4!���������G�$dZ1J��U��tX���,��P<�\��r�q�������y=��6[ȀW �O���o�4�H �D��K�e�l�����ܝ���b�7^��zA���J�À�Z�`�Э��Q�u��LA�f[8S�Rڴ����z�bEw4��ʐd�̧��	'j9���i����Nz^@��:'�6?�l�j�Z�� �8ql�V���,�N����N�ğI;=�{+ns����E<��-q5��W<��h)yD�
�I��J�fΑ���T�C�CZO�ͷ׈k�������܋��J��-�|���QS.�%�����o�k�N{��?Ǚ��7�5G0��a��o���G6���=�&���Q�>u�v"�@��D�����T��U;2C`���?�7gi���"�Z7?�Ku?��XC+��蠦�u��"�e�fg�I&n񙒪ϵ�{��)+V\�]Pْ�0��S7h�g4T�rEm]-�Óƻ���ռ2�����W��P��-�������gj-'yd��S�]�.<�`�I8eR�%^��K
U����Rl��	� ��1��SMi�7+(��ܶĽT��<��.领�xi\�b�$��1?}RO�B��0�oQz�)\-d�0��WCr��'��FK��x���\{��՝���}����� VsP��o�����ʦ����^�t�1�V?����T���>5����(�ט&��6n@�(Z�@�)M*�����Z/�A���R��w"��yWxc�=��&��j�JJ���*���9��)+z�ɑr4Q���*�م�O�ӵ�1^���S	5��(*F�����5�C0PY]bC�V,]��א��;f`�4�qC<�s䛕a���/����!6)cG7��,��x����QZ���
q/���Vv�a� �L#��K"�O�����Yw��򠁅BKAh<�f�*��)�*���xY@���u�����/�m<�x��s�;���JM2�~G��nHH�$[��V9���_���2��Z㘜�Z�,@"�^���S߿<�ć�}�K��0���Feޱ'���DXަ�敃A*J�S���Ʊg�pϘ�&�����V�61��w��𴏎4�f����t�S�_Pv!��/lV#����+�4����o]	k�Һ>gF��y�i�Uٮ�B��;���:����ItT�������r62K<R���'~ɡ�H\�h����)��`�æ�i|~�Zb�⥛��OL�w�Q�\�������ߓ������Ӄ:_ׯ!nGИ+^��AVM�0�i(BQ�O�:��r���L$ʜ�S�9�bs���Sė�!�%�@1�.:�v�?���:���=y�x���#����d��CmD�[Ry"(q�N��*K݂�'{�I��EQ�B��~A:/�;�<�v��2 
��軰�*�R	T��	����g�"P~�e-u�/�Qh���Ԟ�멤 ����5B&:E7��j#�u�V�t�7 ��L8B���N��#��9�W�4YF�[񇴩����/y�E΅B՝v+O����������&@ǆ`�ƽ��q�������{��ݾ]�Ⱦ�$X%x��'�=�-LI2�aط@�Z��MF��c!�dg��A�p�,��Z�҅B �d�Kx�~c	�� #	�_2�N��]~)�u��K2��¤�q�Иl��*G1��37e=yҧ(�R�mRKQ.O�*t.���^�'��FK'k���0-Ȭ����gg��KP���c˻m*�٨3�⣛Y��V�$q�����T9[;�	��vZ3�Q�V�F��w�d��Fu�[�	���������M�B����'G�g$d���晄��a}��2*:?i��(���u��|�%0,�{�[�� �T��ўoW�Ӌ?ޛˎ2�Ti�K9D?u/���s�쪾)�zG&PՐjY�����$�W_6�$"Ƚ��d�q��
ιU�W'1����!]NϮ���4���@�OzB����|P�ꂠb��.�b��W&�wBJǶR![*|
	�7���b�m5¹���]|��M�!R�p���)�xQ�yD�
����s^��F�\�ܴ�Q��V����	`����m����vB�lo���h�%�V�KV ��C�g��PP=c��l�_�aX��ְ��[IMHV`Y�y�ۑX������Ah���-:�ܙ)X?D �#(��Ux�J�i�+X!�o9E}Rԇ#�����[A����v����:��[ ��x͗�jk�.�Xu��&t�t��یgD��͑�_�H��������S�.�\�nR; ��%��y�iwÀ�BN��2��n�Ğ�,Pz؄�@ ܮ�8~[Nv�.8���ͼ���Z����y�tQ�>L�QcM��~d@z�0�^n���E�U_��Ñ/� ��ѝ��N��%lЏ-�Y�*��1��iVW��V�`��|�d>��;�Hojw$�����c�\�4��bT9k<���i��.I��qAq�u�ꏯc58��G�6ھC�W�@S����nї�R}Q�;�\�zO��g6�1�'S����k������.�opTR蛊D�{�AJ~sH�(��i�̖�Dʗ��'��S[��tE�`��>tA�sK�_F�G�� ��i�)���&���X��L�f�!�Kںa�!Ḳ��;}Te���IMQ�;�&��ل��(l��F��xR HZ3�@�&��fٶ蕾���I!y�BwcN���b��F�bFmY���,W�vڃ�:l�uY��y"��X�˼��� �cԷ,��>����߬�pX%�����C�����G�÷A#�J�ea��J�`�r���1(��@�Ă���$�UFG|)53G�wk�׈1�1*�o��4s�$k�
e�o^�J���������1/���=�7^,H�p�e�|{�[��/�_�jk���VHXh�H���H^O7���|62�dh��6-0�k���b�u'���Z̐2Nl�B�����P�=��c��3�w��WN�w>���IA5����>�-�{ #��ڐ�x��~�/�@��;�;	*@��Z���0���D���?f*�M�[;s����	��2��D�Ұ2��Ov�U�Px��4�J~�Fp�Gp���+{9tDz��bfm�l�O�5�� ��'����I����h;����a:cKT);�[>E�Y ��_#��ANrE�5�^~Bz��!>x+�a����Ț�f��iPV�gi�◊�̢ꍤ4���G.�X[ss~G`�8���<��	��@Jm]Y�
1�]/��ze ����eg�
6���t�T�TyМ��&���)�x��_Mo��hT�tw2Mnܛj,�-!����Y�[auZ���G���T�]�1)B�