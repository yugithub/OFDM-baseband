��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6I^��R�Ȍ� �r��ɻ�$a%���X�)�����NZ�(�D3�a��Z�����<��_���$��J��h�*�A{�Uzvy�E#A�	�����A�4\�W�$G7]H)���,j:�K�Ȝ�H���\��Uϙ���s��H�A)n�|��L��y���%�������x��!Sz�����_�-#�͉T��y��_W��D��.G3?�]�t�<t��pO#���ߊ���%�bZl��B%?dk����ju��/��ś /<�f*5��s?�V� >)�!-��Yw$�s�� �V�=y`��ЗO��v4����9�[��fy��fh֙Fb�e4|gj]��A�-���LA1NU	S�Ɍ��m̲f��u	ϒ�C���P���t(��aL1��ת,#��v�s�� �jk[��!0|�C���I�q��X`t�@�9\�_���q��U�K���Y������B঄�«s.W4��}w�<��h'������.ݼ�=��g?d�~��'u�_~AUa-�kцo_k�b���/�;J�B�⺫m��*h�z��}-�,4���S1����@�y�%�m)b� �w)6�V!
��u�~fh�ߢ����)� ���T�mE��E����/�G�@"ta�Wr="�d�� ���j�re��4�H�`p�A�
2 �ػ ��]�(Hj��q���Ɋ�E��$h�>���q-�8�<�ErQ8WR"j�>���a�uH��%�_R3��+1��z]���IҔc%8�t�� �&ۣޮ�c�F����d�(j���4v�tO?~��yp�ʖr��c���ֻw�6٭X-O��0��~I���]r*�D�	4�/1�w�-�3��2偡BI��@
z��ј����\lre�?^5����5���i<?�n�"��$p���^�>c֘�h�>lʸ&�,�t��~I�۔|=+>��d��Um�0���ݸ���@�w��6�<dN��]�-R�h=E��rux�P�>G��v��d���0�U�=.2�����8.�Gaa�-��i���k�Yy;�1��Y���!��a��K�!�k�2�K	�oa�MI�H���5�u�}>�1�"����<����~��@���g�^�E��v[�V��� ��[��oI�P����%�3fC�'XA�|�� �}��a߆46�i/Lty�i��������
��ùZ�$g{���j��j���9�vgWv" �vܠ�T�p}� ���>�i�5� k�I������\� u0�p}xs��6L���Cl��u���Ij����\�x�g���k�W�h@߇�"ki���"i�����f���STj�g^g�{���NF�^%����k�\C7���q�߫Fc�Q<�f� -k)�[䆸�����/�*�*-,$D�O"�~x�}��v(N�;UX�ȳ�Te6�R>��A���`D#��alb�#u�nO�'�.�+�� �k���U���b�~���ECFk	e@������Qg,��7���.;�����1����t7+��C�>�� �Ǧ��_���HА�[>Y-djO��B_^" O��8m�R,�}/�}�����ؒ��e���ר���\b�&��=r�i�ce}�������x[i��o+�>�A)�(��W.�� #���Ƙ-M��&�(n�<�+��N@I'l������G.F�yH�@�`�H$���%�VZ_�l��"Pe�&.Cՠ�)��"����������K�˭Š7�<�
D�&e@�^ba�	Un^�%���Z�5kZ1�*���F��0_b��F����� ]�opꑑ=5a���.Ss�-"��SW8����'7���oݫ���Z��o��j@F�;5��n���qȏ �Y�*������GS�HL �E������֭���#�5i(;��Wz�Ql�*l� �E��1'����8��Q��S��Z�+2�$Yu�U�,]lFv�?��DH|�:���*Q��3Y��B+�44�^����E�
޳�Փo���G�f����;���]h�T���[q�t�I���H���} �S�?a�Fw��
�;>����_�Ł>�
aP�灘�D�F�r�܎���ǻ����z��<��ok�E��~�U�)v��Tr
��>P3�iyw�7v�"2g,2Ɵ����q�]f�QǶŗ��e=�X-�Q�mL�9��e�Lm%M������!b�A���}K���hi-�������=�l]Rb+���D�y����?�2�����}F��o�솃h�2�P�*�r�i����<}�.�����ryp���o�2ft���؃�m#$,���F�KǞ��U�49� J^���z%�
RK��:��]�z��@#6��Ǣ��Dw�2�Di��k~�-�%���8����˜(�t��a�,�������{uX�JJ�<�u��&-.��*J?Ŵ�5X3R�P�QF��<������t����2�S��\}���!��=��龞����J$5� S<��5)]������W�,�4�x�K�O�����b���*��K��q+Q�3ݩnLZ��<|Sa��Z r=�E�]�i�6'NԤ�tM�8WX:�Ϳ���^�3W\1�{�[����A��L�R��5�r�Wݲ�MB���Vъ喾��|ˇfsX<����st�yQ�BOGm`��s����Ѵ���t�BH��[��  �b��.��\ tJ���7|�ġ��]o���q���j�_t �!8�����j|i�׼��Z� KC�A�*FJ}"��W��	�1��U6�����?�i��7Ef�	��Y��MC�?���K�"X�r
������9���)Oq�)<��T+����7�]���n�.H���J�F������_[��`X>T��8ћ�W*K^���N��ac|�?Vqx�+��|q�����s����L-4�~J�����怬�*�~�!�U�ޠl��_���q�@�A
��1�d{��g�&��YH=.l%�af9��m�[�������rjs5םG�̪Չ�H$�T`q;Q�Td���ա���l�����S:(:�a���.����܏Ɏa-2��tb��YB�!�Aaj&�KO(I��t�'�?PQ�3�8��k���Ij��l۵���v�g�Pl	�M�`�?������\��5<�B9k�&b�I{��X)^oԃ��lçC�5�Knύ�n�7�t� ��5�����U��1���7��a�[���D���Km�c���(��ߐ༐��p�/��W��Y� ���r��`��M�wD0L���'P���5�>�O���q��,�,�/�q+5���>���7�X'�mNR/�s����+ %^��1��WoU���������y�;�� e³�>D���L�����&����K�YD�s�Gi�q��t[)dl-!�]G��d��-�H^��z�!46_LvAk� g"Tn�DG�n�2̓hs��A�I�N	�QT,�d0���OV)l�wo*��&��� v�V�۰iKi.]��Q�����Ƞ,BĀ�{��M���n�O��I`�����"=GW<Ć��@D��;Z�ş�?�>���mq]շ<�b�%����ǿ�Ȼ��f^�s/z>�׻��'�J��܃,�qF�3�DV�?c-z1M7� �28��7/2iU��v��es8Q�:��Ę�|?jb_��-S��%F^u@��g�LA
/���������E���P���('x��[���w'��:ݾ��H��N4�(�d���F( 5��i���g�Ks1�*|��ތ)]��W=f�Z}��_����Q�:�֯���	��2�m���Z�M��3$�˯����%t����J�?!�]";���V%��B�$ς9�T������Y�߄��8��S�	(�w槄�c�|�n�Z���L���������F�mۧX�;"BA�&L���WWEC�'��K�|=r��Ve��KF���K)�
����(�Vr�x���3'�[ ($���*�S�M�;_��,�����VB+{ZU�v�;I���<�N#,�bY�#���� ON�*�H>%r�p�����6?fg��@�YV��ǈEr3�S����m�ۍ}����/y�ɉȧ�5�x����&��|�{Z�9����F��z"�ﴖ����[D�a0ٶxK�ل�S�t�Ǐ�vp�iL��7����:��d"����I�9'P���=����6'����|�Jlv�}X�x�B�	Z�D!�)�������O)�o���HA�L��G�&�b��jZ����Q<F_�����E���;�+����I/� �C�9�����Zw���vl�����<^8��
��i�^��&m	O�j�f��g�����a,c�{���"�)����i8 W;:��ech&��w��XsgI�a�xp�E	�@�����C�s3gy��
v���`JI_w�e��Y��+��C�<C}OI*��G۔���~+/-Bh�;r_��%���Tb{��_��S�G�������A�߱�H}aGIGʟ�N��#��vҒ
 բ�A�8눲�v�^�<d��Tø� �����|6 &.Yw�7�~�cN6��΁��w+�>Z?�-"PX'��/�fi��vY�?V/�>l��O���E"%�3��;�R�D`��dy�M3�=�՝>�[X�!�3���}������W��R^;�ќ6σ�I�b	�tJm��ù/��0�_�6t'E��q⪻g��бu[��,���obQݕ�F2�uh����������+�VT'^��ٿM W:h�9��H��"6V?Iې[�fdR�y�'��Î��1=�c������X�4,B���
/�iº%�i�7�ܾ@��� _��R��3.�zn�a97Ƚe{e�#�+}Z4�r�<>�zkl	o��MD&Q����=7�N醱��*����M�qu�>*z���H�ҁ�xjC�-��3��fß�.H�]K~�س�>����>O��kM(j�4~I^-����J��7�[*�\z���c���7�5��(e]~`𐰄�l���I���`�Fo�+��nʽ�S"#���ո}U�N�
&)BXju�GF��p���ax�7��us&%rd��%,�ۡ�5���۽�ho2]�ZO�������A}2:�% �l�lS�}�rpvǶ�7� dP��m����k:�91��5�a�����V�Ŀ_N�ࣝ*���u�s;K>1sI�v^L5�	�O�Hzi*�Eu��=��d%e�X��|Kq���˝x��]����Ɛ_�IU+�%dLw
�1����{�./mb34m>N��fp'Ho_\܏�p�x!���>ݥ������{�T�n�)7�_��m�n����������&";�Ʋ<?B�Žl��
߆�M�Эܗ��,�y��	8�Ͻ��M�۩��u��t���ݫ�t��_Z�fS=���+ױӜ�4`Y,���d��KG�v��~���n��fi7�p�91>���:��#�T�adWm/�����GV�����k
�o�DG}Z�gн��i�`Q27�w_MGӦ�+R�9��YPbT@bZ0��S?0j�E��"��>B5����L"e3��q|���on;�O3���Ӌ؅��GAeB����S�`2=� �Vn*tk�se�/T����`�
�1������VM�p	̕�����s΃�E�ֽ���O�ˬ28�f�E��5S!����(��"��ވx�rI@#�Yt���<�^����7� 1����i&!�����8�UI4,�x�}�֥���Յc�q���T+�V��RC�("����5��+�b���ŷ�p�1����0Ԩ����@޹�) �����7yb	��ct��rw�7��[�S<�}���)����}�P}��xvڸ���x,L��L+'�Ӡ���fdm�@�����'.�a�A���h%,�m�jW���v��l#U$b��<e���r�t8�I�H&���y�7�\��L��
��1!�b�8�c�Y?e2q9�<�o����(�
�w	ÂW���
j��zѪHWԐP���!��:�!���(Ge�
������稟�v71T���F��@8#Xt��B@ڣ������_*:�����d1�&X̩ ����J5U��^��#�t�q&!*'�=��C8�0F�#�Ec7TM0L���z5����:g���P�]��d����3~k�a��>��O݌'@�㗑6vp�:�����DC���f0�h�u,��� �x$ ���� ��r4~�P>7�s�^�n���1�V�/H�X�LfV/�܋�,oG�*����
螉��̔Q�G� nb@?�Q
�Yv�,��t>��1@�ߧû��˱5=͈3vf�m�#G���;�,�)ͦ����ReH���}%����ː�z-���Yȝ��߇[�,���U���W �@�l6��p��l*���'��aÕ�#/�%��J��Q��ϵ��gE°��OF#ۗIf=V�AW���w&��ϰ&[��cmQ*��[%�ut(F��r�h���ǥ��1���/W�-�-��^x�D��VN0>�I~2'1�!�!JO�v9�*T9cC��%�P�+&�!'am�v�d�o;ܯ<8��C$����tT����������Y�b�Xd^o�R�_�=�&���R���*����������	O�ۉ'K5' �����&��V!�V�m�������ocC�^�[L�(&�� �b�].r�c�G:&[Х!�}��u �� �Z��i&,gPoX���a��:|Nc����F�ܺ���kꭾ\���_�b�HF�n᾽�7Sy��������H�uX�C~�Z�!4z�����x{u�_�(o���x(��[�t ���f�����Svl8�#+
�����i0��n߁�w�d�ٸl]�$��1Bed�s�J��5�4Ĭ�ĝ2�p��gh����H�z���?}�*g���U��.1��eUu���N�ƿ�S]E�gGVN[t<i���"̶�TNt��V;Av8�s�G�9q�[�����C��]����r�c�?0�X�.����:^g2�c��8�<�h��H?3<9�2���.�	�#��cX��-��Ǳ,@B6R��Oh7);�|Z�6��s����V}��ڬH��t2��~�PY�R ��P����C� ���,S��"�L��a��1��<��YE# Ǆ��xn(�K\��S��N:�sm1
l�)]�\��yk�E�3�Zm�.Wk�~���J�m4MVI!���:���{ �)��1j{��\}���dk;� ��`�����?��HcL��^?]J:�(R������kP3�C��Z	xɿ +�F��)+~�~����=�\�KHGɅ��ԡ*�簘�3}�<���D����\�
"7d~�2Ԡ�z�+G�@����
t�ʄ���P�'�{S-K̥5�����C>�ő� ��M.Vݵ�Ō>��Sqס���%\y�l;H�w�����GQ�Ĉ4��̢c�������}�����k߿��3qs�X1~����`ݚO�~k-(��Îy��e��5uc�T�1Eֱf����n�&�(q+\�#�ˬ� �T{�8_��hr/��'CT��{�=N�Ƨ}`+VU��<̅{V�c��!�u�<�paM��t�q��?m���fU���"��UbQ	������/��(�!���r9��׋����Z�!ϙ�d���5a3����E>��7�kwc��,�_�"}�p�E}�E�zYf\���$ƪ����d��B�+A�aDf����o��ӐĶw���]�i�b@�)���`aLPV���P=�Î�[jP������g�VM?�g*������8�h��l-d(��QJKK(�	�;|�׶��y��h���$W0�k����':�ǟe����ZS�c�U33jv�Ż������U���akT�V~�]�%N٥�B��,����]�G�]�+i�Fl2�{N)��+�<yc�[�ra�RK�f���?���	�����ta6��K���>�)9[�U�D9 �!�8��]i*Q�yK�U2X5���*���p�fф<Z���u�,J���M;�v�Fg��ڴ�ԙW�Z�Q����@����c���#)��8T�]N�G��Uߗ����@�Z�
�����H}��f���I�a$���K�����LϾ$��&:t�r_*��%�s�0�o#�53{��6ͯ�_�Y��7�@M�e4 �*QÀ~2K��g�֥��,V���	���u��3���W
�L����G����z�U�`M�;Z�5�����Wp�M��1�SԻ ��3|&�d���@t;sњC9���mi5�Do@��3�!܂>���.��;i��]��������۰�jS�w��!%/�I���T㖕p��x�|i��9)������)�hOn[��3�B�5G�TM�C���u��&}�f8%=�����>c��Y1X5��!D�Q/������M�ưw�N=Ƨ/�N�m3[�ȄP�����wHӨVɎ�p\�_��_�+�n)�1�ǌ�c��x:]=�1�GNr���y�*Z�bg�O�˿���y�J�H+���S�r�Uoܚ���~���
$�o��_��� Q@u� ;f0�O�L���-��5Å:����r�R׫d��I�ܾ�2�e�,'�����d(��2$yx�
hǪ�	�"���Zi �=��~x�h֤F@_��;�6�P�wqS��)�P��͋�䬤��#�Q"�ݞ�=Md���`�x�<2���[$K�p֊5j��l�]�y0=Zo46��H���D:SeV��IL�����%�Ŷ!�I���>
�,Х�K,� -�2�hf:�oH/��
�ŗy��{��׈�u7hˁ5��!�Y�&,�^�Դf"�l����������m���<.�+��@�j��x2=^M �A�/��G�>���a�a@u�^Ir��f��^�&�)M���s>�F�7��Y�������HcZ�iARY��LW����[�`����݃Y\&�4�t���dzj�_��iܯnq�{z�~ 6��^75k0��VՈ'�y��徾�08Y��A��5�rO�ҏ��P�E��<����HQ�.��0�E��3��(���a5�ܖ{��t}�%^絓6�RN�O�1��f�4[���t*����M*&�Nb��lP�%O�j�;> ����z�9Q��0�!����º�K��/�#��;~/�*�+�A���2�p U<����3P����ǻ���#T�v�z.�J����X���u��f݉�y"�ûڛ�x��� �jD� 'T���%��'����<��w2��]_S�h!2��D�eN�ቭS��	*.�n�
�� B�v@o��S���r����q�$/��u��1h^�x��3���T�j��d@(pf�P�CG��S��g�R�RL��`Tc���;���?�D5.���%�Y�,�^�s�[ۻ�~����3f��f:�u�ey���j�;
V�EZ&k�I�\���h���'�wVC%%'qB�����kݯ�(&�꾜b�g+<�I�^��dP$k��V��J�ڦ��$.�^��_��q�Ʉ�Ɠ�i�/5f�!jg��
��L�#=�d�IQ��IN�F����W�{%qղ�U�+��
}&��窥����=7w���O W_w�p�i�+��3��&�Q��j���|�{�������p�q��`�4'c�f��4��ug�W���N'����G��Mf'F��((�!� ��O���UaB�*�N�w��i����Ɓ��W�>^�뭇cá�^S⸐/ u�FGU��6� Z
�l pG�_�o2�޷�@{��7�L�7��fr^��YgW(?`���[E�L�)E��M ��]c���K����乎���t;I��'�.ŀ�]D!���k䴌�����h�p�:�KE2���b���]�'�.�9?�8dD?$;}4�p��.�����d�s<�I����1�<=���\�����mv�<T�0�j��v��^��(����N|���~OCwp��*+kD�$��b�qq_�a��U9����4���p�O� t���M=�Rݓ�l{�Qa)�S3p �lT�O7�AB�^�W��iq�q�w���͵E�<{����]����56�����v�D`n�gm�*�������2"��<_�t��o�;�@2\���aI����3S�AtW&�|חD�I�����G��)��@Öuɓ�T�z�_F{�*�&M��t�f��]���*B�M%���E����ˉ���<�s$�<�_�����K-�+�?�3��k�#��Z"���1���)�TMe���'8)���m`x�R;;Tm��iÏR�F(�g14�}X{�3��g�ݎ�0���H�\ElR�y���g�L��&�ES�;�������D�zO�<��숋b���9X����J�Zd���X�0�S���H��ՙ2��E�+�N���n���!H|8�H�a/#U0��µ�z+Yո��[,����%o��]�e��k�b�ϊ�UV��u#0�L	?�Y)¸����IWG9՚Xl(�Jۺ�8% ��x��q7gM�TR��r�1j�q��8�O�����K�`j�M���"[j�8KK��h�.1;�7Vh��\��Հ-�1Ѭ���&�9�ڥbw�����{�XR��r��W�ԏ\,$Zt00�8(_~���[�ФW��
�$���i�^}r�Q�V���3O�߶���˟>�;�k7/�1��}[=��=(�7!<�{ߌǤ�������>�>׈�j�bXG�9���P֑?�����t�PgX�?��"$�U�P�����%�|.�$��5>����:�*��W��-�KiiU,&g�vA�0��3��2�M+�l?��D��5b�&��=�f��V�CF�!��Z��s������70p��bGX���Lx�K0����s��u�?�I�LW����3����P��|�@�/@���.|�c8��L��1E��OY3;.�Q��YqI�\g��d$
�,G�Z`j����;�G�|���c/i�7"�I//������!V���E��Q!��WŽ�`0��
 0c��+�z����l���φ����6/� ����B�\L���I���c7�y� ���Q�'�gﮜ�������o���鵢6��%%����;��ҁ%.{�����Dj,)Oqx����l�X�lЫY�W�̅�6?�ț�`�*r:�7�,F��1<�yzOA��f�SҎ�,�2c��m$�(�c�ԁI7��V��Y�|��mZ�l�1���� �"1�l�*�@�|"b5�l��62����Jdq/!����S5ު�q/��DIuVs&�+�����_��8u�Kw�� �7U}�� �����Z�Յ�x�H�< ������'37wu�&�j�|�_� �ŉ��ɂdQ޽��%(���|х���r�U���h��@۳��?#ԗe�K㴑�����l�( +�S\9K5���Q��������uLÓ������#l�����	��H��.4`b_��}�1���n��+~6$cj�E���Gǭ���VZK7A����vDB2 ���6����Fz����|I8�YW�R����$�^l�����R;��Jx�Vh:��@:����ͯ��Y
����Kf�2|7b�td"�b���(��t��e���w�ۉm<H�՜��J��).���̾X8�T�ם�"�^�{��FFb���G��jE�)�}ܭ��eWf��I�9�Y��峨Sv��ֺ@8A���`~yI��MؾӮ��P{�w0w[�S�F������:�a�d��n-�>i��2�����TW��d�(:�X���d�@C��#�R]�O����]��zb_ܼ��}��&����9���0�w� h�~�Jot[C�w�l��p[�x��kF��Nw^��F&��P,�A�n�_�4��81v^1̺�#Nc�:wz	 �
H�h{(QwQq���C��ء���R������8��P�O^��rO�喩�L�����ݷ��mPk�Z�i�{�@� �Y~U�sǈ�5����TK?��N�L1�a_��s��5��w6C��'�y�Hg�:��>NѺl�PQkx�w5d��P���1h�K?�ո�%��숄�4(�ޔ"����N��m��>�(%:Xo~�8c�a��ytdxĉ��Arp}'Gmd%�����ߦ5���ځ��a��w��aJ��K2�v�;��KW��H���pݧ��:^�3���-%�6�	r&������b�C�p�}��wY�O��wZmW6�ga��&����C� �M+c�R���pW�J]_�ɼ~�T�G��K�iO�����:�'Ѵ�Wۢ�]2��W_ItLᇽ�"��I�C�ȸ�~�F�������V*8�O�E�t�)JnR�E���H�Z�k�єy�d)Y�^�E=��A9輱��UJyY�0^1�2���:xv��Y�a_�q��
���&jxF�����6gqî?ӉB(3�J�ե� N��0U'�n��ou�8W���c��RS�t���=U��e[�a,��([��*�.���6�O�g�~PgN��O���֜��X���������0yj�<]�mb�eQ3ܫ��p�����i��ݞ9h��s8W��,m��ߒ��W�eb�~l���F�ˤK���i��y���2�)a��W�j	�C�w��vC1�&��1)�վ��l����J��M�NO��r��FmM��.�Ut�\��Y�����=J����p���x���K9@	elAI+P��P�%��*�	��/��
2�4�27��g�7��ȣ���M$��AY%�:E���;�Y�IL��M�D�G���\�oͶ��k��9�y��|O_Bj�;/�?Z��[{���w#s_r��e3����g#�����>[�j��O�A������r�;�<X�l�e�d��Y�!I��6�y�D��e�_��L��M!/��������T�è��h1.��y���:�����`��沍�45�{T'�O�w[6� Cx��~OQw�%��!##�Qɬ	�<t�|⌾	ݣj+��[��E�x��dŷ�$�� ���a}ܗМ��� R�"����8�c�k�p�6/��t��>#X;���)G6d�.�xmcN;E�:�a�B��(�%vP�w��>+��`�{�6WvBg�`m
���w9���ɐ�'I���\l��lM9qZ�5�B��y�clӹ>�����H����QB~��Q� ��B�_bHJ��#D�pt�b��C�i_0����Ƹ�����ꪠ�8����\�E���ە�cݧ�ct.�mj+!����h��h.g~c��1�V��1��0�OT�s��4����&�vǷ��|ߵ,���'y2Z�?m�6�� ����dYR�h�䊛ύ�@�T���Hp�Z����P 9�	����/E�{}p��{�cO|i�l�Y]��1���W�l{�;�	ٙW!AK���e��V�
ɔ$@N��V5^oM�Ya���I�Ke�c�[u� ���G`ǃ�5`�?�b+�j���A������Ǘ��%M��N�����Y�L�%q�f�DԨF����Y�&F2�B��{���Kxt��Łk7�b�|7Ne�����G�MA�C}���ܜ:������b��$����L�kَ#�c4VGucF�����8�P��Q��s5{�(%Ǥ��-�6T�X��Rf5��X7%��77�@�uHS�R5�
�q����%�К��E^[���Ee^L��������Y��V��(��+6	�֏��������-��nBG�W&������F�L��Nb�VVN�V�at�L��u�j��
:A�����������Ӂoy�۟[����"c�CW�x��4N�K~N ��ާ��ǚ�k]1w?�|C���5�Su<������Ǆ#�!��])���7̈́��Y���Hdn;g�[�)@GB4��8ʺ�yi�Ե`6��0
�`RDL�V��.�S�ۧ<��u�V:}*�^�̙�ps`[[���}2��g$w��wT 9�vlE>
i�#a�g�θ�R�&��,�mD�����er[�@�M��]\)����a�$�()����F8*P��/���Iռ��#O8�	��PȢK�ס����Z/��.]G�y�d��9�L�PrwM��b��	��!�BD̋�%
�?J�U��6��'��K��V�i�*�A������Ӑm��¥����!��g?�4��a:��n�]_�E5�l�x�,`�u��L�.Ӽ��e:�i�ܒ���:����}��2ϥ8�
�7̦��A�-���a����蕢�ny�m�y:;:0g1u��(݉Шp��g@OW͗��Te꭪��u_D=#�#-]��>?�]n@]n��d_�3�i_o���J�׊�P�B��02s��� 7����Υ�[�2Y$���F-�(� ��h�ӈ��`�Ӽ��>͹,~�'���&o�ʎ�26�	��	��w#��(;���~�jf~�\�7T!,l� ���pp��퓂2h�Y&�۰�o�;=�\��,���^�p_��vv�^�y# x�ca�J�*̈�vUR����4�3���(�_��P�(_����Z��ܹ��P��'{�3M6S�@����|��E1��f�Mp(S���un@�7k�Κm�W�n_��H�y��ő{.JB� �'5$B8HB$\�m�Z�OJ��' ��%���\�: �T��ק��ْ3#鈀_1/YU>6>�#��p�s�s?�Oc B6���ҽ߯_-�;�S�s+>�[:ݝ��	�����l3�U�����zN�)$`j�ιM�c`��Ӵ���)l0�y<��}�	���Xnto$���%ZL���L3ҏ��g����v�.4Ϳ�=��2�}�HƠf�i\�zGe��aj�:X7�99J�W�<x>�a(�cv�Xͱ���{ų o�4��\�`�B��CƼ�<�Z�
c�@��'�И�Ưs���a%!�D�
�7E��A~ �R(|�u��P����e�Z�h<b��F�S酥���=����P=�1b���+�($z��kT�l��ͥö��A��«06|)`�'�V�.��.h�d0�0W���ں�y$�P�J��9ͱ�U����?�e���C�G;���ԝ�3~� 9�VT�7�:��.��_����En��d���	%��_�!Kl��Hw'���W}�y��.��'�)��bi�2��aE��l� I��G)�L�g,�oJ��e�P�tmܹ��$O�:Եt[�����{#�抻0��O�:���Vp��*{g|5%�����d0#�����*Ғ��r�p</��1#��<�%��"<�?-��իO���?qQ��?��N����}����Q��n����8Z�>�=ԗD�Y3`yK$�5�@��y� ��n�(���ss��88�j{�6t�_2.-���}5���>�F�w]&]c���]���[1�0���u�u�1N!y����B�C��75�fu{��)0\�*��>�E��26V�6�}�9���P"�<���ɭk�:�@2U�K�'dU�x?Ym$��O*�S��^���$e�RK�n3��R ���&�6���wE��*�����!��+��t,a�FE�P�詎�P\8�*:�*�����a����IM�L��3|������W0�e�}�>e�q������`�E�J;�t�s/8�����8���~D�y���L65��OK�P�@�>:F 
pK��	�:u�_?�����v�mP�h���֙	�n�1z�%� +�Kl�\^�[�\Ԭz��ĉ)����@�	Gq_��{.��~u��?�@L&�x�[TGeva��x���k�@a�Dc$y<_ �2�3�+G��6m������Xq_��CE���2�p��a����"��g'xb��V�� E�_��7dDRcB�LB���[L{]a�l�'v/i�?*s��!u߯+K�C���S�"�1�͐~�q_����Çm��qe�.��S�!�_+x���F�y*ii�n�����cq|c�[�0�b�bez5`;��'1cذ�w���F5���g/��<D�8�(��P-��C����3C(�Fnr��g<+ӹ��-�am�L�V+�[���Sě1�LP�c�kSR4Cl�5�Ǉ0 ��Ic>����zp��D�28�˻$!Jҽ��)���Ы�
��g&F�9�հ�:�A�Fv���u�MOZ�n4i7�!���,��.k�ƞ��F,G>
��/��u� ��2�K.$�A]�RFX�ѩ���%��ė݂���qr��\�dts⛚���Φ �^�@0e�V%E��'����<"��;d�۝J��~=6�Ɓ
��2�
��ߣ.�H&-����X�)���Ӱ���p;����'mZ8�g�o�
m�x���:��@�S�&`:�F��
�js�)�cc����ۋD�_�=pc�S*:�^��B��3f]8���q�J�Z����~q�䘋YP��`����-X%�V�Y=��.�Ԏa<#y��pB�XJ�@�[�����z�#��>L�lD���΋�u�G}�,�0Ӌ���c���Iܠ���x����=`�|�'�y`k&�c�ҕ��{�u����l�~	�@d��u�p4��T�t�'IMq�"���t�FݒI�����@�'7�$�5��s�J�O�-��Lz9>(>ЏN��L�z�ȉ����f����*�[ɘ��DQ��X��<Ֆ���5"%��6!gY ��aǈ�T2�p�;�'#|$�W@"��b���TW�
��	z���������w���ԡ��W��r�#�f��yz�5��em�d���q���\�?vb͍Ƈ���5zm���t|�D���`������-��"]]�e�3�m���6�V���"������ڥ|4�؞Z띻����d�]�̰$V���I�d�@�J�Β�*w���
���"�"9=lb�{0����]��u]$Fą�C�[z=�샰p^E��T�gaI,V���h�X0*K��i�) ��#	f�#Rf����(�ĝ״p�/�4v2Oh�F�Pqd'O�S�Ai�i>�U��F�W0<�l�PN���D��ޕ82��B��O�����X:��z7N&'��غ�B�5�;\�lL�-	�;^{��qʬH�,{ޔס	tN�,D���� A�%r��p�"���}��v�('�VT�S�H�_u��e��3+�I@����=���Dq���zr�� �S�U<��"��-�1��tp�8PqB�"��6���Ja����2.;�$��ynzy�܀G�s�iW{m��]�Z����A�������V�N�F�Бr�(�$�������$>�vWT8��E��ٵ&w2�x����eGI#� A���g]������ү(]if���B���X��G7Q�Z���S�#�Euf�a��lf<}��<���;��ظ$-gA��Ba=u{X>^Z�P�����Rɗj�΄8tt��)��_4�o �p9�V����]�E�|?��./[M���HJQ\��:A��˒�KE�����N`͘��{Śk�Q�lT����ۚRϗ��1ns�j�"��[:py0�K�Κ������B���΁n�B��|���>��B��S�ÇDZ�vwD����Q�x�|��1i�	���v�w�w�E�����{��j��e�=kM�G��O^�8�{O�6�0�������$M�q}���L�/ge���ײ��#���X��J�L^ˉ�-��[Zμ�y�����rXL|30���,d�EH�3�������8O 毅�;&X�1�@)蒘��
��;H�d�rM0�	f�M46~;��g��֒"�B�a,�5>w�IGGL@�I`������f�/�4�6�X=<9Y��MՏ��y ���3���].
N�V�oպ����r�Ap���8�+�/ϭ��e���[��M�N�WlEk�>R���a����ŨcƔiE�*�SzO�+�R/�-L�x�}Ai��J��_:%�<>96�P�y��8w>��?��j9%ClHʔ�5����Ӿ�u���=��Y�Q�`.���o?5���tZ��Xة�h��@��"��X�K��+�j]',} ��"��z3�!�P(�����VD�+gs��-e���-F�kPZ�CY/`��-�ǜ׭���Rj?�څ�����9%5�ē>2���:����AB
; 3��ﱝ1��#+!5�a	E�a�G�Fv�tY|p�E
�}/w?Àb�\u��=1�Qh_�����4�樿~R������7fB���Yܑ���E����Ձ[()W��׮� qy��r��w��tW4@'�V%"�����V��҈��u�r׹�F6���2�𜜾��o�`����F,���ġ@GἨuD��9.��悁*��,(V+��D�C�~�n�`pںIԎ���u�n�a������6�i�A���I�7�v���3��J�!��Wz�A��v����}ap���3��VVtɨ�J��D�V����� �AP.��1ޤ]�ÆQ��Aͣv/q����6軎�㑖����E�K��2�C����i���%syLi��G9*(~ީ	}d�|h��Oh�q���*Μ�Dy:�`�+���Ҋ�N͓�>v6,�p"���;�z�i5!ro�Q� ��A(��#�TC{,u��F���+)��<�3`��S?#�nUȨX�~g���b�;5d�pJ���.���ſ�y����sMF7,Q�Ɋf��-��]�������&�+�]x�8P6��(������=��9��.PG����[	1g�wTjN�����^3h+/:��4����m�~lq�y�Db�y��;'�x:.����8SSR
ם�m�U����#�'dx{��r%|,�r�7�-�F~l�?Z��ב=�C �B�vl��铺�>M?n�$/����^	|�q��-��C�l�Tᢤ(w3&�(6�R���"ϬT�J�<X��d7���2,z��ʭ���ͨ;ڤ��+#'�P�뷊VO��B����'�@{GӾ��7p��Nç�LT`B�+�Gذ��;S���^	BI��)��)���7� ī�x�%�k��.'��e�.H�:J�����I�~��
�a/2�}-�yd�d�g�MB��5

�Ȝ�c.r-�&�����D�+����ם�Cq�u��9�Gu��8d�E5���@C�N�#)���肑�����Z$)M���BV��|�#<MG��Fw-:*@ ���p��Ų���?�4�^՘���
t\���>�9�	�,��u3�)2gJ2?��#�#uV�!j�fq�ْ�� �wI��XٞV��=]���%�;�>LP���a�p���m,=ǁ����VIx��$��M�+9�6h�I�8M��R�tǱ'�f�D~�Y��lK8�K��+W��Մ��ӕ���z]�0�;�R��,o�p��l���?�I%��+�G�DIcfO�[���%�\d1#�x�7q����'ɂ����Oao��7.���"1�=Nhn������S9BH�6H�^<�f�<�֭[��d��|�Z6z�8Fc{���f7��2��il�/�
���E�C�o"���.���iH9�j!��?�>�,��'F�˒�exO%U�l)���,������;�9�5O��:��	���u;4�d�g��_ғ5U����@�~n�E��J)���	}��Zu���ڽ֏��S�.'��o	1qtN��a�����A�����-8^#X)2���6tf��)���![0��PH.߃%� +h�p�S�=�0{ M:�@��":��k��>sKt�l���7��jB�7]'�g��q��G������O��%
��#^S��(����b�v�{x|�����q�wx�|�����}X�;f�X�X7��`���N�J���B
Bl�ڸ�K��!(��:��F9�E��!�=�[�!!�Y� ���yh�[�L*S��I���V�x��|�~c訩U���'<p����&��!�^�=9���t�B���bp��mx\�k`%�$��bL���f����	4�)I���9B��	CS�V�@be��|��Z$�e�>�O\2�w�U:�4�Tp��0��ރ�:��"�$1�"�>2J���_Ԑ;�ގ�kc��W�4��7_ɹ`�$���\��u��U���^t2���J��koㆃ����t�(d��%��ӂ�Ms*�|X2(��G�Ȫ���vN}(��W�w�.�1u{�~��!p9�	��#�mmR4�T:y�.T�G�sW|a���j(p���3Y�Y2Vд�p��hty���CUN�}ԺB^�΂:p3V��kT�ʮ��~��,u>���ś�6���oh�r���56�	\)�&����E�,��V�`7a��jw������L��=��kk�/w��]8d���^��rz'���`0�}�*��i�����%<D8d��G�3Et������'w 3��v��+��ēڨL�o8�ۜ�@�-]�߇ljd7�4q0X�ϒ�;�+�sw#�T�����\���魪l��GU`Y�s�X	�/��(t�v��������9�5YΨ½HIfO�"%L�}�����S`
��!�d���a�Fc�Y�3�>�ǂiJ]1XkAv�0�.��g����%D[Ͳx�`L`�gܕGUlq|V�<Vt���	��h�k.F���s��`}��Uhc��a�>�������'J�G8*�����ugh	BU��{��8���1�66Afى���������������I��Cw#kI�V�����r��.��x.z{_M)�rD:k��}cnuP�r�ps׊ t*V(/����f�էMt���0{>k$�ʎk�ߏ��;�OA8�S�Z@�s]��@L�Í�	�C�m�n�`���F�G(����\���h��`Po�$B���2�I<I�ֶ`ñ����b���K.�����8�.��R��E_�R�*��y�����g&���]#��Y�K��d����q9q���=YW?]�k�-��J;Yz %WS�0�a+��v�
�,kf,���R󈥻װ���HI����.]���������6���Ls"5okwyV��5��@��(tt�;]���(��S��0H�6�K/�Y_XE������<[#����F/�$k�f;:Ji&"�Sɭܺ���!V�fF�~\�ʉ���M�#�����s��E3�ap��;
�,��n�4CB]�'$�є��an,�<B���n�O��v�?,�?Z]���0�M���.ES�1m�[�k�\wo��L��P$Ik���#�6��o��@ye8n�az:ecִ*̂V_�'��ö�ꛇ6�B��˿0����kPe��-�5=�vW'�a�a�&���b��&��}��H�T"�x)���[@6�WĜ��@gr/v����Ɂur�p�cj	Z�s�8zח�N�_:ȹ�`���0$0H�x�i(N��K�
ϧN� ��A��=�J��kՁ�	��-�NJ�����4�KPO
�Dѻ�v����P.+�۫����D?�菾�:��6S��b�?��fPh 8r#��&[�H�\�)r�_�u�)6;HTl��V������S���.t��*u.��"KK�tY@���O� �	v&��!��V�$6����&֟�ⱟ�AL<�NKKZ wi��[*w)�0��v�X���ज़��^$�����Jo��%d̝�D.i��A�-���QG}�� �Ta��l�d���t�B,s$���(�We���_C�'>�~?��;��_��N�r��Yⳮ)�=rR� �9��:��Sk��:!��v;-�F�q �߫0RK�7�l)���Q�Gz{6FTm���٬i.*X�"�N:)�2&�����X>m5�h���0ǐ�E�Uam(��1���K��hm�!�|�;	�ecI
d�Cs|	p�$����B$�H���0l�:�Jp{��j4����ӡ�t��Ϥ5c�%v��D��o�}5ꜘ��{��Կ�}5/`���$�.6�ʵ����q�e���Z9������l�h]�l�� B$��"��vܯF&v���
ćc�"��kH=5Ϗ;������1�}q{�QM֯ڍh���̪m��5xp<XG1�8듻���kN�צH�/>2����n�0�Ν���+Z�K�ݗ�U(�2��|}5����)q�H�!ڄ����e����㇠i)���緲�1��;bΉ�/���{@O��t��2�!WS(gt�.�Kn�#\F���Fn�=��=j���awbK����ԚZ(GUC��2w]2L���h��ܲ�c@��w%�����ӜpM�,�<sts�2�gO���d�~�����1|@Z�H<H�)^S�hM㟺�ǎ{ִ�q��$��yY�u����]�F9����K�q|$Couu
(�l��Lg\列o&,��|��=��K"�gD��&�90��bPks���f4�NQJ~@�LJ�t�ȝ=�<����� ��̧�T��ԷG�.f��q���@1�1�_L��ލ��b�N��ܗ��L����K4��-yN�$����'Zh�'B��L�� 询��3m7�5g<k�n�2�H��������{�P��f�9�W�5�`e�?�����2�����٩V��_J'��ޒ�,I��%&L���r�(��C�Q3�,[j�H�m�/���䕗=���ꉦ��~���C�I�j*�/�YP.Əl2ȫ҄��g-*��za!DV��V����i���%�䞌9��\iL�q"�ق9v,���a�]=��̞���O�M0��Y��*��^�W�iSo%�.A�
ƝI�,l�ܤ^p�:j�B��&�x� Ԃ�д���;��lm�GI�08��lV�9�K� �d~��{wW�uf�#�Q�R�WZ&��iŴ3�|X�d$�H-4�n��"�>��&ì�||�@վ0�U�.�&V��!_�w�B��b�[�I<�㡊ʈ�*�_�&��.d!���`6�s_��ͳ3a�eG#�yB���ѐ��J���Ye�!ʋxY;���ϳ�b�n�2�Ϙ�n�2Ϥ�K��,3ÌhI��W
����F��]��V,�:ܼO���X����/��W�@r����56KA<CU9l�1Zc=�F��^��$�|\��l�y�W��{�M5����O,
n�4햵�ҡ��4�J��k���U�����-ynz�T*" �IPΗ{B�������D����o��n�⩋U����xg$�we�"�vr�ɡ�w%��E7MOr�1f!�!^�_���^d��S�'DU�?2j�&Q�W�R>7)d���s�ڪ�I��^���x�`g���o�/O���y|����<��6�(o7:��S���N,���f��V
��T�����i c�<r�b����w9�Uz  (��Z��ZH�L�Ϲe ���WU�|�������t����|�N�k�Sw�Z�V�Y�-x���F�𓷿�����1}կFK)��c�k�=���y���5/wج��Q2vs_%��Vb�&4#ȏ�?�i���C/��S �S'D�s�Iy��	��|�A?��G��@ߛq%�I��2�}�1D��.ź+3������{��|,�=�%I��I�+}y������[���I7A�g�pa-�Yn�'6��=�@е������wsAg	�U�" /��Ǉ��\��m��ݣ��g)gD o������e�n�@𗓹Z>+�A��i+V�]@��������f� sb��d#�b������ҭ��d-�pX����_m�y/ŖC�3E�d�l���:�ՉA�(������+�jQ�GA5���V]�R��=�Q4懜�X.3�L,X�$���yH�uS9��n��Ň�1 �vo�I��H�g��#�aG�y�V�*��-�noH��K(юF�`zd�.Qi(DX��-��������s��1�E��hM<!Ň�4��P�C��%"
%�k��u��ȇ�\ʍ@g\��wϠ�v�w�R}5��c1��>ӛf�q����Þ�Ħv����EG���0��z���T�K`3�/K�Z���R`�(����)�?���т�W�pZ��G�*zO�ǟ~�13tU������0�6�rP�>Y�r��=�[�����K�0�'����+j�k^5h��#�&L%r���|��P�tR*�!�X��;oS���!L�E�̡�XQ�����9�h@�g��$r���Q��F�g��:�����îP0V9Z��[�R�&�����9X���t$ݔ��f���H9I��5�]'!0�5�-V�9	�(l���� N���Nǩ�'�Jҩx�eF�?m��Qu�O'�o>L�h�яX�BE��[�G��BT�(X���[�L�<c	��3���6)t��B�f�^�b��ζy����0�I�(� ��Pv�@���j-,a��'����9����be�z4�8˳6A����8��`�)m�g�(��;�A�htB%��sK����C[�G��Ͳ=�rjiեh^f��zH|��:�1���_2N��i���&�J�H�w�� ��D���e��w�q�'�!�$�IP��?QO�"��ouVVl��(��?^*XZͿ�=�j���@@���������Rm�9/5)�Gu��F/�d)�&���N}P�����7�+5&��0p�=�f�0˰����Q0��|p�\+X�G�ߊ�~��9����c�5�%��O]�7[�Cu,��?
ʩ�� ��.����ú��C�N�{��>��$p����^�+Thqe�p��K��$��LQw������w$��������lD���z�zg��h��&��A~ج�Ի%�^�w��A�l�bT�6�D��P�k<�������Ԙ���J�,���諜I�G!���)����9� y:�cd=ug�Z���=Js�v�_F_�տW�K=�U��|��� ����˜.�)��M/v]�a;8yf�A�45�RQ�Ъ�ʹ���T)�E
6'R3{&%��C�7�p��ٍyZs�ԛ+**�yr���^��d ��1�N�t!��\���[KJ.���O��+WJ���3��@L�4hE�H�]Xk���?|f:<�z���?��<�ʽlU�{�������M���6)PU7k�X�r��ۂ-�����띦 -a�J��������X���]���K�j�-O��m�K�C�T񍯜Sc�s�T���MsO��`
��(��+z�M(u�(?X7��9��j��&��J�;��ǶՎ���Wѥ�%]�0����B��G��ψ�##�+'N�76.t���)��M�^iM��7W��Hz�)��,�J�='Bi&j'�K"eL�&3/�]�\~z�=��f2��ߚ��=����̘ϤE렁q� 	$�~FOP;Ҙ�zg�j�J #
���Qy�ַY���ܤ�������x!�*��<��*<��yS��yy����T;���v��-'~�vnA/K�p���@�R	��U���\�n- �3A�*<a�N1�\�ɺ�3�N�h���8����� :s��nD�;��)i@�r*ph����|^2a�x��ԥ����Cf��a��e>�Oc�JړNjȕr�ág���ES�쎝�4�
 ��/w�K�r����#Q���x{�R5�[�M����t��We14Aw�P�/,���R1�ҙ�ׅT�J�X�+6q�]R�߷3uM�����|�<Γ��Da-E2<�"��rM��q߼�Nʙ�(�wȆG[%!-��������=�#@KG�~*�,��H�S��`��p|w�Ƿ��yww	7���_j��6���Y������< ~�4�6X��<C���fN�|���Wx���D��Ú�p��Z�����9�uF굓�
(�)�V^r�K�Mɧ!/�Í��65Π>]��ǜ�i盧��HR�:�a������z�3;��l^�E�A{O�LLu�������^�,�GL����]|B �*i���E�9����4��~!��c8۰y����r甯)b�d�����ŀr\d���'ٸ�`6;�1}���#����i�<x��#�� �q�K�����X�0Ot
��Jď��ÜJ�Pw�2<:��'��� �A��m�&�����  3�=Y]IE�@�4�P6�a��ޢ]�v$Ƙ��l�C�o]�a�J�]��+nz@"N�>E�a���2)�,FV�B 8;V�`�@29�|R~;$�'������Ո�UFjYʅ�����*~o��&� }���}z+;7��@$�������e�C��A�+����ʐ�Է���Xo�?T�`ki�ץ3��"��(�
e�\Z%x��Q+�Aa���h��ԏ�li�����4�{���Q\�DJ9�ǛЯR:����)��6����8t�ݏ:Y�E���Uetʁ�FR�̃|s���A�.,�]����������ك�[*�[l�#���F���E/��F��"|Q�l`.x��{��wv���0���7��ͽN�u7Բ�����8)pR8)����	�����G&��*��!��)�ͧ7�-��8��$5�Hc��7��#�R���%��`����� ���o	��\K��(��Pe�R��f��A�3��Q"�戝�`�H�Y h�X��DA���9���0Л�@q*�[���b����TQ���y&�9�í{�w�MF���f��U�Y<��b��*_+;I�(C�jm�	5�濾���+��󲸌X.s��GA���'@��ns\_FYqp�L|�<]M\,��� �������n�c�� >[�p�N�+*��
�lp7	�@�>���A�ã��Xۡg��U�� S���N�&b!�+R�ݢ�>F}L�y�d	�>պ��(K�a�TBx�m	��G�9]@���2n�>���'Z�=�� ������!�8�~��1#�4s�lJM�\�b�G��;q�*��bj�����2&?�u�O��6G/�����E�.���g�����h�9�˵70pڝ�g�^�w_4����"v>�Z��\8RI�-@X4�>M�4�sO���P����L6�#��IЕ�.o/��J���`�/�r��no��dp��y��
:�lg�3��[�P�90��:�s��i���K.�x �L�ސ�Dӏ-?�.��������46��8KS0hΐ�|m)m�C��fШ�4�$�;��T�}�������=��l�!aÄEE����}������$P����b3M��l�j�7C�/@���=�U�\�cI&�����@���e0]oo���x�.���y ��9�歖�J���Q�=���q�u�`Z�<��\���"�����S���n���6�Ь�\nf���,���1%�s�TOZW�.[ힸ����	���Ӣ�?�5	0���k7�V��=[���&��~U7|���Ao�_M�1�e6�V��V��OX�����HF����о$G�1W̛|� ɘ8�;[ꕰ�A�o �^W��[}�X����f�H,��^jz���H�&_�o�!����C�O^�lG�N%_"�!v��U��~�{]ha���+�6�m5S1�:��u(awrF�r$�ˌ}��g�ڥ�4[�u�p�m�56���aj�h��7B-&�\�ɥD�^�W�u2gZ�	�ݗ��|l�#{_:�N�E7꠵ �HhshLrHh������ՏH�0��*�&�@����B�e�0;� ����1�[�L#���i�]�"��l�A2�ÐJg�V�3��6.�{��a2�u<AY�-x���JFq�X4�gXF�'�&m�EN�I)�����H)�+ه���|prb�);&���1g\X�Xb<F���8�uv��+�&�6d����j�I�"x3^��D��227��L��ǂ)��o⡡�����p���g����sV�B#�C|�����}DV��h:}L:��v,�g�E�l��p-�F}�^ی���f�?�S@���)��<��ղ��n�h�"�Fw %���r`�9�Md�so��Y'������v��@��u�}&C� B��Y�Nr�~Ͼ�~E�j�I<��R\`iB��͍�:�q�S����H�y�Y۲4�4YuH�{]V�h�6��si8�a�C�+w��
h����}�w}Klӳ�Q�w�JD2�LdMG�����"�X	|5��q�o�@�L���c$,2D)~>�!�����YnhE Q�JЩ�Vt��!�d[�L����������x��@ѭ���뇢y���3�Ϡ�T���ެ���@[+��.X�����'���O�u��_6��U��w����F ���|u15�x�@I��ez��D�M�9{�,�-3�<�C#���-K�ԡ�wWʟ�6�R��k�~ц�tPzD�l�
R���B���Tô�Fl9@�����V�@�,~��>���+��i���߇/�����?&��L!=k�.)�$b��)٧:�d�)���L��f�/
#���#R��*2��#���G�C��k�N��VoFp��b�����myP�?��F������	4�(�03��gk��8��%�꽦fU3�D�6�UY ���BEʍi@O�Y>>?������`?�sjMt��q���ɫf��d%+UL�$��({.)�Psu�2��jVt���S�(�q��j��2�Lp?"�7<�(�v"��O�l�&t_W R�:J�����R�E��G��������N��#��Ԡ.$qha��Uj��#��q�E�g��(˅M�7��k4U	�b��OX��ͤ6^.wn�p��)��iQ���a&�J>��ܙF�K)T��#;A���_O;��j�S��-8����&�h�O�B�/�}�;+����^ʴ��|��B�Ӄ�>�������n��� ���#�i۹�S˜p���ᇙ��	�S�����//�4�Ό89:�9>D��Q�Cy��v�o�)���>�EX�7���øv�����Ÿ��A	2� �P����o@���,c��M��p�bh�����D�.M�=��՜%kg�7��i��?\���:��a��u�q��b�4eD�R7C�|�b2�!o]�9uAm�����>cI�s�`9�C�T��υs��K�|��ކ�[�E��_��?�3�9�<���:���ܥ�����}�ng$o��A�lǳ�����G�XOv"�}���0�ȭ�e�:�ױ��Ir�(�������1�Y�����]l�,ϛ�q0)�FǎҀP�g�!}L�T@�W�O�K6�rcl��*��u�y�_��fA���N����[�4���iǃy���#`��8��¼*";l{v(���K�<��:6I}� �>E�#�:�p��j�Q���dA��'Hȸ|�����ĵcs0$�U�!��u�m�تZq�_��H�X��kv��4(���{� �X��@��2o�*���R@(�xjKΣ9���(L�N$V�����7�K���{�^�)��`���$����oN���>��,���k������o�rT�D��ӳ�#��ONs�4#�-_�MjnH���B�e��rVZ=ɣf����n�q��V�0Z�=��{D�� B�E��0��Mj���'*TF����cYt����~�<kC_꿸���O���(w�\�~w�4P�h|Զ+O
����9�>�ҥ�L��
.ҟ?��zH�{���/��q0���lve�sǴ�g5x�P�e���<p���:�]��ʌ/�8�Wy�)AF����/��J�0ի�%�`���=WҢq{��׮>�pg�!v�x��A���yJ�T��	~E�{Hz��g�����1����Mjx���ύ� ��V�H��9>�_��O�p�oV�1S�Š��͍Y}�ɗ�-���v���l0ta��>Yag���j�����60�s1��e��fA�K<+ �FF{'۳i2�&J\�#k��%H+��1% �Dߓ��s�o$�z>�г3Ѽ�ק���a�Ŭ�:�b�9'�r���>C�Au�SV��@Y��8£����D3,�W!���tPQ����v���"�n6�ٞ|�,_�[����_#=��ߘ9T���!xF���-=�:���оdX��
���7�K�Jo1��k���!l�����ۆo���h2ʆ�dݹb)�J�x���)6��
+=�b�BN|]���gd��V?��}v�M�^iIy�D��e�P�?�6��;G%�t��^ᄠ��F���D�ƻ�g�;�����g���"= x�r��,��|�*����aب��E����u�v0���c����{2m�E�{�p�������J�%�m��͚CO�9�4n�U>j>t����F�>���{���8lv28�eU�%xf}^xj��׫k�[j�ah�C��I+�����S�-�A�Ͻ���.�P������zJ������#O�X�5Q���pw��R(�c� J�?�σ�w&�,��g��)��I�����]�)���8��ϬbA��JC:��d|jf����R���Ý�-{j$w���������ߊ����m?���\|����;$�>�8M=׃M�����:�%��5��(�n6��ȷ�^��gr��e6i0�h*�E�**�0K�N�U`�W�U����f"C��h_b�-���/��n/�0�r,Ƃ���6��߬��-�"��F�K�{]���	�C�EEen�{�,E�>�b^��F�[�DR��B��E$0�Ⱥ�[��Y��Я��.;?�+�][��tG��m�>X�z6����[�g���5t�8���]J�+���P��{��Z�1Z�4/]S¼�QZ��(9���摸?��H-Yi�`�P�m0^�!J�������g��=��@0:�`�z1�1A������9,��ꤸ�޶�0����}� �qTB\EG��/#fw�G}'s�:�A�t&�H�$NQн�����v� ^/��/���*p��.x��H�1��{s&��� ������J�ʼ;�uȑt�^b�ݗ�1�n	�u		p�ѻ:�SʫY�z�M�HHn�~B�q#�Ӕ���)g���dY��� ��m�5�=������Y9�����= �F�:Z�>����O�a�n>����z�K.��&%�=�.����W��G޼a��^�7%�{;↩��ŵG���g%sX�D�bv$O�j�W/|�N9 ���hƳم��������n�Q�L��^��at!����]&Ѽ�V�d����V�,�_G�Dd��(cnd΅*![)y*��/�{�[�/��Gy�����)�ݏ�4���x�֛�X��ZMÞ�y�u�t�qD0�JN��8g���=�A��ڣ��N��K�����	�0��9�_0���fvv��%���a��V�u�#UO<�%��s�-q_��5����Q_��~ڝ���.�$�b����K�B�9�蝦�.`3��Q5�5�˗�x-��F����|VS'ζ}U]᣽���	x{�L����1���Nu! ��Ɨ�22�/+�/qK�\i�K �0�9�@�gҐy����� ��z��,�㦚U��f4������p�n�\_UW4�=b�,iR|��|(A������;(Ҥ�8��>L�hv��Ԝ��1>�BwR�� �(�|��Yl �asR���xT�<Gq�<ƛٺ@������O��r�hѦ�n��p�c��������e�oZ�����jf�-1Ȕl�̣�>k��gL1���k2	s�ESKu�NRޕ�	P,���Q����eM������C]NG-��(�F�,��Q�ɨ.�[��m���"\$v;���]�3�(��d�R�;4����|�ЕH�`�^�&�c��w��v)��@޶��Ss���aa���&��s���o@�<� �=�$����c~���|��T�z��	F��I!l�C�\=߿�u�z�%�99U�Z�����e@���`��JRP�a�~���]	l��jԃ4 2;��X8m[7a({ m���&��z)�����+�v����7���0��<���[Q�EL�.z�; y�*? ��^�3��6��`P�{}%.5��ߣݕ\����tB��~s���oS0��~�H�������2Z�F���"�U-�'�LهǝA֧Ҏu��������{��X�p��IǉE�N�O =AJbi��ǈI�~,�>���6�����O������Ev.�dx{D�[�lt���78Rj��gg�7Ф�����<����	y蚶=��pE�˾b�����l}_K�z�\��Mb�����لf��)�ٛ�c��^��襈)�p��oWtk+�^
�<ϒ}� ��ÙGJ�g�GR�~�������h`���,�>�$6J��w.�#������;�l�Ҷ��j��������7��T:���['1�Gr)�����s�$�K�C��6!�k�\ �D�U
��'� ��&�2�F)2��i6c�',� �Z�M9�����t,�7��Vr���/���Pn�:���މTQH�Eqp�͗�f{��1�aM���XH<��)i����̹�я��������޳k"�궍��Q��_3�um)�K���o`q�^~���7��\�C:�d��J��tu`�3��g��"1P+V��Q|�ei2*��:�DrSb����[�U<�ʅ*���ԇ���C:�k��K���n���c���}�;����Ṝ��}x�}� �)�~�rd�9���8����3�G��p����ChP?�5�k����)D#Lz����<y��z�$�>��g��|P�Ǫ����E���|��	���5&��\@K1Mvv���dhDUR}���
d3�WrAo�M?A ��UY��R��"TE�Ѵ����0x���g�4��x��1�Xu�L�+����u$VǶ����Cz�D�������ݾ�	'���C�Z��@K'��;~ȵ\����?��|��.ś���|�a��=�;w��$�;�8�?�*߿�<se���	�/�hҪ�8��>o�����K5�_��i��Q�1�.5���� �7�c�1�Lk���YP���&�h��@�"�����|v������:.d^�
�8��M��\Ϩ���Y/!����:�1w���u\�痴lWd���6$Lab��ht�� �c��K�(2��n��)�^��n��P#����4����%���_�M�g�����$�XK�UE<�9ΐ�?�HQ�8:*��v��Ξ�t��n��<(�����j�/)C�H�d���&��r+���|��ǋN8ٳ��O1�S�s��+�""�p���<2���g�1V6H���c5�+��ȱ,9�Ȳ�y(B���Ԥv��ĆoA@�R*��<�f:�~��yQ�%�A��EE#��&�WJX6���52��w<�ƍ�M��
2L��4׆AF
0C`��t����G��u(��׮�uLD+���![�����hr��E&��?�WG9.�q%�TQ\a-�3�Ê_��;C�щi%�����
O%Zc��i-�)?�_r�2��f�p0F%�7C�گ4�����v���<�đ�8i�y��WX��al�Y�AV��p�Qc�L�s���t�����<��	�����_����Y2M��2�Eg�Z�a��%�B���T�5-�=2<�ܳ�	����9�y��\q�:	JPf�*�����+o}K��B��>y��˼PC�#����Oe"��0�F#�'���8o6G͂���������4��5x�A�P��%O�������{�[�G^�14���ߟZ1`�^�o��9��T���Z_}�8��H̩�rՇG#~��3��.��������T�R.�W7!Td&k�"�*��V�J�7v�/�a�e�Z����Kn����3�m�<�eC}���kxY�E�gَ��� u[�X�����|7Z>��jd�ߊ�ߴ�A����~#Z�����2},Q�C�~�(㯗8��s�E�*&Q�jr� C6
T��$�� _K�XЊ������;V��S�*s�t��E��R����@��������h��]��#��z+�E1�>�G��	��r�4��w��
Gp��i
},<�ʟ~Φ��ԟ����>>zIP�}�P$�ܱ��ڌ{jw��cJ�#>�w94�
l�1�oS�ѓ�0?��6'�+����Z����s�Rڋ?�p?��6:��1c�&�]v}֪��"rsr�L4�{G�IGB�(Wo�G楋�t��w��IU7%S=E,93p��w�!AF���槯�{����9��R6�? ў:5b/��l_V�=+��Gj�pOe���0�L��P'1�]�g+��H����&��|����?�_�o�Iş��7>1*��+S$oEW����ż99�Y&�wq�(�^������.�%�����qR����.�=;}��>�}կ�NPX����&���ͱ�Q��^WpM�����:E�^�C�'a���y�h�5��r3e��Z̓��ph���h�E�`S=W�kI���|��5rt '�NC}g^�7�LQe��W��B�M�U���4�4Q�yF���p���[oG�A����f�$���.EF��B�x�j�xkghE��ϲ��i���t�
U�熉�j�k�N��qݧW)=艓�U�>A���+�[L�J��am�PN/q�
�V���m坽O� ����:f�(ܨ�q0��3�[ ���R� ��E�|�sM���͉' �Z
�G��eF������'I���B�_��d�μ���^V!@9ݡ�Z���>�D��w���J�e�񎌃^���5��K��0���K��������ڍ��p]�iƵf�q�����J�p	����5����B`�f��d[�I~��X[!(�W4_�L��E� \�?��,??Җ�?r��n��@[���it'	?���h��.�=��� N��#�d��h�b������y�R�~�䣂i5o��D�^�+�I�����l{T�2��-^�����PP6�G�E�R}=x�4	!"�E�Քƞ��� k4��3p�V�X f�X�[5+�,��LS��~���Ϛ���Ϲ�Ze9[_��@��'~,sB� ��t��YSf܏7p)�s$+Y��z��A�|<�lZJ�[!Vt[<��v��YͶ�)��}��O�w�.�'����r$��o%��o�-�ua����%�2rJ��<h_�b���o��PO�f0HҨ��8���m��lM��AV��S&M�	�E��ƈ�=�������&�Pi������DW���9�vB:0�T�d��G��3Y������[Ku��}�Y�%��������j�9���(,�$�xF��W'7��Q:j�c4�:��L)P<ӜE���t,<��5��Ĥm"�tʚe��Pn��*Ίׇ�91>�W�2�n��ؾ�2�
������Ӡ�����iK�1����U���i}2��=���p�Y��_���ȅ|�wX/YȾ���D�M�%gwV��8أ��~��5�K����ȍd�7<�?�IS��f�/^�r	��kw]nU�>'�Wc}DKhC�9��������wP�^���]5T�[�'�l�T��H9S��xПZ����D�B�J���i$�nq�{�p4"�L��\�䑉�%=��6�(�֬Q߄-��rS)���=8�lӦ��=���N!�B��]DhlA%���P��
�����g��u��C���8'�z㣍z��%�:�g�(�� �.��Q��*�čЌ�� =�!��*X5�}����x��P<�M�"�]�@$ �<s��xI���Պ��X}��ݕߠ�cؔ̂�T?~8��Y�.|� M���%b�S�+�UL���GoĒ���$V��n�F�� ��!��s�����iZ2�E��0LԪODn���:Q
�J9�a��Π�!:j���}Fw�=��O�����貈��|�(~
 ���r��� ���ߢ�胒9���$�r)ձB�pC�R;�ӷRCe����3���އ]l--���qf@��r�}Q�Wݗ��4w|b _;~6����IfR��7�QK�lŋ�Tam������!\��Y�bM>���5M� �c,����	It���w"�b>\;��a{@�����zd��H���&��xh�u���GH����c[~Z*E�Z�e�u�(Y_\��Rn(��T�)���]�#p�2�5X�d`����O�\9a��Xj��[0�{�ذ��-�D�f�l):8����5\�6���e7C�s>s��T�K:`�ڄ*��8i���s���}�=B���/H�֐X������m��.B�T=�F;l�`����k�>n��uÏ�����'r� �{�迨�	��W�;g��4=��X>\��Y6�;��qS�k����+��ߺ������:?x̯���Ě�uXW%����"��4'��h��+&�l�q=r�͚��(�/�B�w�=FT�:�JU��Sݾ�J̰��~ޗ2�m�2���]\]��NN&��\QRXq�6%��=z]�Q��y	�Ê��ZUfկ��y9$�R�Zωݨ����;���ՌNu�@?Y�"��x��%4=�7��\o9���G�>�Eŏ�	b:	�N��c��ZƪS�T��,UsPL�tB><�GC�yu:��:�q�:.n��ga�i�P��i{�Wǘ�/�l�'X���v�\�֓n�~1��돷nh�Zl)�-�α(�8��qN`��8Rt�Ɂ3de�9�Y������|V�
���'�{ HC�_��Eab^�޴ ��s��7�#�"��z� ��~��Yx��gpIM��6�O��^}c���[u�-��=��9�a"��0��YS=���ǒ����ū��k�ݡJX��xo����i)ʩ�+�O?�r@��� /NoM9��d�0�3(�J��9�.���l�8�c����ʏ����U@�"�C�����1�W���v�f�����ČtuIlv��0np_��#��h�+W�U���%m�X��S-c���iTh����!���e��mTR2��=�B��-ˆ�~I���+�[-�����h��w4Mm~�e>���z�����
�Euf��m��>��~P-�9�P��6@����k(������_t*��wÎ	R�!{7Y���˯+)��'�v8��C���SQa!w��Q�ꈀA��e��?8%��h�8�'n�mA�kY#�֤�~�+��5|�#�T�̶7�H����6���d6T���t�>`:���6,�8�N�}]��˽�H1V}cWr�f�8��Q�ty��3�CJ5��� ���Q6�M(�jRYN_�� r���|���:����cP�ea���(�ն{گ��d�:`�~�96HF�i�t����b=7M��?i�SA�<U�1���h�8��M$Y6�����j����Xk2U糣���j�czX���2�"�cO�:�y%�+Õ��P����4V��#�'9D�5���Myベ��i��HP�.ѫN�k�NZ��������ܧ=�P�%�f�A�L��dY�pq�]Ys\)�ҭ�3�*:Ng ��Е�m���D�8݂.�ڊ�i�)�n/#���5Xú��(J($ݦ@˻_�_����	o%pO]��/�:����!T�v��k޻����J��Ͳ��S+�%8?b��e�=SC��.A�$�i0��B׌�-��T�׾�Z@���J���ؕ���,��3IV;Ķ��RE����\�?�J�x~Gm�Q�[.������Z�G��4�t7k��|r����_r>��Pɡ;��z<��6���*�8�P����|�v�Q�\���"�:`i��6\�5�%q 
�D���A�+��9z/c!����&iU�|S곤�+��s����$�\$�g�����1�\T �jWY�w7Y�>%�XgA ���.�m-�s�]YG�*����J�kh�qM���������x��U��gD{}`5_H6���������đ��5�A�;�9�Qh�*��z�,i�>��Y�gT��-a᭲�&a�i�&���fy�z2�� �b��R�W���$[\�-�Y��������F��_�AEЋ{�l�ĈⓏ����6�l3=�MDyf�+I�a����\9��������|�+����`��z���f��w
A�Y0�D��)�$a��$ �d0=r�n��q�B�H��~��k�,&N}5ʓ-�y���	�&�U�͕�56O�Ɖ��L��k�^��T���N����@i3&�qX�v�#�[�$�ެ�z6�eH'A��X�S�~� �LV)a� ��[1i��I�Ї�/y����1�������]|������$Âdګu���D�=B��5�y��(񏻝+"��Xڇ8J2�&�����%N����q��"��"2��у��'�v@ǩjl���|�罽v�g��2{����'����mG�/.M��IO�Ƨoü恎T��)�T�L��3�u�xo\9�*⧾I���Bg�gB��ѥ��K�߶dv�`�R5HvD`x	����!l��)9�:ia��T�On'��T%�᧦*�\���M�\�P�������F�5���Ī�E���]ʍ��(W0��(�~�[�:w1�Ē���m�6�G�z�mK�ރ;�NlUT��+`�M�Z�5ݚc=H�� ��x(jS�%+�[-���GP�0��z�W���	��EM�������D���B[���=	�����ɮ"��^�Ӓ�����2�д���q0
=��o�)�(�������q�d<�PZi�v8evƜ-���������R�1A��R��2��}�,b�D���6X�U��G����mE�=p51�����YX$���th�1��g*��"%�y�%7E�?�A����_��b|��?�#L�w.B��A�yQ$W y4Gt����:@[B�9D��O15���S�d��	1�-�y���h{2J��w�ً��gΚ�+4���^ߺM�腥q�T-�0$�!�i�e�x�}b��V�G4�@�-��Qa�4�㏶�ҧYs[��n��Hu\3��#�3K���B.��G�f��,n;r���� ]��P]�0.�J����l��_G$�՗<0QH��!��=��������dg)�i��\��1���8+�k��18�R��y�p.f)���蜽57!?�&���#ip�Z�	��%k0��ɓ���^��X �d�t�X�P���ڳAE%���օ�ݘ�����d�4IF"P���~��[ݢR��,��pJ����$�ե�)�̓ރ���F1�	��X&���~���!�/��(��<l�W0
ht��o ��'���n<���E{�S�Lg�h���䗎�i��������e�3n��(yć�Q<���u~.��mؼ_�zg��sx��)Ro,;���U��/�6�8	��^� �ʤn�|�q�A�/�mW]h�<����1�j�P�+6���E���#ZVBRN�^�ؤqX�H֨���"x�R���+��0�RA{����2�2����??�d����ml��Ɔ�[w ��o& �s/_t�%�}D:o
l��B�5�KFLw%+X~�!hV�.RK
>^���X���e�.ɺ<��м=��hl9��px/��"P��+"����M�����d���C�y��čV�D������V�ZKܧA������3�h�γ�jM���Ȳ��z��Y�M����Up		
��� -��>��:\�Y߱O�1Q��p�-0�x&��@��{���od�0�ӭ��.v)��`�4wyP�J$-�T�A�,d���˭��R���sHP9k�Z�����f�ղ��q+��8)��)w���]sӦl�an(��-����(g3����Z���K���pI`�nQz�!��x��4P3h�3�Z5��|�.J�q}��)_��,�r��?�d�:��M��� �a�G�@.��Ҹ��n�Xw|)�
��y��IM���0�}�G�Q(�N������|��--�%m�[��`�|m/�Τ��h��x�J����eId�nP	�}Z���V���Y����J0�呋y�	1������w7Tf����F[���L���~7k��r�!lLE?�_.�+h��"~��q�-�O$���y>�_����  >�4-���*�x!�Q�p����$O����-��-8�q-U2��ݑՈ�Ǘ���ns������8�j��1��S�j���Y,5y��K`ѽm��u0�&��#�`�@޵����먴ީY�×�����k��ޘ�ן�lC��E���"�F�@����n��uGN�k��vn_�t����7r�F�1�3�JMdt0<�EXw���;��"�S������b+������ji�J�-U����|g�eoT�<�0��Yg���4n3m�s��G�H�jY��^^�-7�����*/)f�����6OR�Ҫ_�LK�Q�䕁���O�"n��Rc!�+�"K!u��{T��05��mHr눃�ơ���g��W�c�%#�J�(*��)ƾ��þ ��}9���z.��>���>ZI�feY��b�n��'��ef� |D; ���nް�U�4������	�$��Tʻ�k��T�@�q���h�s3�yÉH���R0������ߛ���K�,�{L���-K	/��7s�N)2Ξޅqyi=�pQ��v��:*_���h{4\஼Xxէ��~���@��s���ӿ��V���m޹'������L��L+�܆0�ؼ��q �{��c�H��%��y��T�$]��T�N�q�c ��q��:�7�U�I�]�=f�;LqT�z�u{��q-�V�e�[j����ۛI��h��ݍ0fjBĹz�b|�$��-���mgd�7����y���a �/�����i[`n�;v7���}����s���y�t�𷻑Ө1�s�_�F_���i:��%AH����Cj��\m��8w*Ꮦ
+p�7��k�X�|B|�[����Ue��A��X;��%���/�b�$�U�������I�Sn��?��<W����ݮ�u �tTaZ}����k�����*�Dڸ�y[�u�z�OJ�2е �8���//��:��4�e��1�X��(/�8��p~5�AGf~W^��:��[ �c��^٨7w	�����E�ߒ�����\3UY���Ў*I�J/Q��w��2�~��²SVHo{���� �0���.3�½�F���������eg�E��p�Q�^x����,��6� �'K�r\A���x{T�t�!��c��v�1�*S�2'�ݴ��`<c���C'G.��Ц�5I��,a3�FyI�U�T����2tI�5�E�J���y��G~Oq��a���:>047�uomV&<m�\����$��)��>����Z��p�V�),�l�FA!�m�?�� ��9g�t��X�)/��{���N���A����>K%N��h4"m��|KY.��&%����,�O�) �1i���
-m�,��֑s	|C���`��9=N�Q?�1=;�E!�?h�߸��~��c�8�G�$�V6i�*O��"�&ސ)?�ǎ�oM��`sH��:#C�2��M�mMD����������c&���-+�K��,�$��g�U	�c�%�35��L��&!�����e�>�ߗf�J���!CY��Wu~"x���YTq̲��丮0���@�s^$�i�盿���I2_�U09l�	��_i�"�$yv����c���G[�J���L��/�KVd����B�5�5x�i��D�'W�Dm�!�?qm�M�ɓ�qJ�L�TC��e�-�������[��W6w�^wH~�π+s9;ƞԁt_6���ɛ�a�&8�t@KR�[8O��V�Ts�V}����t�=����0���敔Tbs��#�v���Z������ɴGE���; ehE����-%�"͠SR\�K!�#��9=����9�i|�C��_��R�!=�MR}jQr����� Ú�gU��,l�.1L'�%X� j��ꉨp6��9�b���:�td�nF�B7>�����-�CL�E�	���6���o)���L�'#Ta�	DM6�-  ��,X���o*'/���Ԋs}ӗ�� c���ur
�.��f�[x!��_�{� ���٦:�!�ۻ\�6\�È^b6}��	�Pe�ޜs���v����|�v���4���s�F�̬j�O��8Ƭ.�[ǂ�����1�:2�@rxv9T��P�3�z��?F!�Za5�7m��\,�4G��Ođm�R*���9��;s3�2���EQ�ojp����?��ѿl�&	�H���&�q=3���Ͼ��������U�|���i��M@�\���\+�V�Κ�'�c�K���EI�x:o~K�o�s@����U��Ⱥ�'�6�_3��)��'��Uqݭh����y��[�������ĳC�q�u�m]��wy���
{K|~+تCA�,�9f�k���ZU�q��uC�&�.�9w��P���Ҽg��*6@/�����5C�^ͣawu�֌=����@��@5�������6T~9�D�>h^�:$�������^$(��ejx�f��]z��PٛIƮ�\y8��?ZV-��4�`�*sd�G��j������M��7)���e-�Μw8:�4q�Ш��ų��qB��<ى�f'�#i�.�|��%�p���B�NT7�e�������qw�r���?�ǡ�b�B���gF���#�р��P��������y��VL$jg�4E���ٞ��&�)��47�b�i#�>�U��n>�����`C3���`�$���A�Z�J����K�q��E�R=Mc��b
G7��<X.�]�[��<�01�"�b��Ń�iY~z>oa�Gr��ۼ�T�����W�d�z?N���u�T�i��������[��F�}��\�d��*>��)�V^eʥ�%�_@}'�"�## �B������/�E�l>G��|�Ъq�ۣ��l�!A��IG�f0�����^�Q/�$C2`u��¡���&"-{�J�X�h��-&�*�_A(P�d�����+���C6�N~8^��w�W��aށa~�5/��wg�<ؐ^�ٙ&0��Q_z�ZG��Y�8�������xx�(;�b�#��(q����悙�e��{���g���!�4��[�76�W�����5@ң�pR9S���L�w��,y�8����grj�§������b%����rk �(\�+=�'�HrzC���ĺ�_��3�;'� �1��{����"�^Im$P9⨏9�/s^�| le�@���pi�(&�_�#d�E@g�f��ZZu�| ��&�A�N�k.���H��ɛQ�ݚ�&:��sX~	�>1�r �E+����܅�2@����l~g��A����'4�=i6%l��������8�����}4�b���6�?}�Ӟ]]Q�= �o"h�P4�ݲ3�{�5T�o>O���]\�4�y���z�Ì�%Nɦ4�k�B1�ѓCl��.�t���@�T&��Y�8������;�$e���bT�Մv7���_�|��ܪ/h���7�y\w}�L��E>i�E����ܒ'�7{�����L]��-zE�	I�;A�����w8�I�٫4ߡ�䕺��&a����PY�K�fy}X�A�.b��X�[Oѣ\7p/w������Q_�ET,?	w΅�ݩ��Ȗ݊^�4s��/�&>2L-ӌ�tt�C��=0i��_���D����6Vh[\��n�b����+�~Oζ">�0uɨ��/�B�l���3[ݾ24R��(�����T�O��c��P��D��y>1oH��@���H�&�e\y]�� �c�7S=�g��EI���?.��Ɇ�.��xv�zB&�~��f����txEX]�n��>�sj&A�����s�V5C=#���Hld6*�t�0���'�'���Q5�L�V��tus��\�*c!?f�t��S��Y��< '@��Ҽ%Eʐ�!�'���xFt��Bq���4����hy,EC�*|2��c�1�� ��q3a++�����!'����ȝN�f�]���3ޥ����h��g�J�D�bM7���I�ڀ�!���%#�rۉ����1�8�ợz*�1:�`X�,p�o�ӐV�������)o�&���x�mi��`����bH�-i`�`�N7��_�6L��9&T�hGO�����ȓ�pyOuʳT8��(���x������k��YV����o��~�!Gԁ	N�FPh�GH��(uڟs�(���T�%���ѷۣg�^��$}~�"�������l���d@E��`�F��#���c��	�����=�@�2��Y�@�������6Lǲ�Bade�d`T'��Z�%�J�'n�QG��a�Im,8�SSp\5EZ��U��~�3R�ܾ��\ŀaP	!�EA�e8�j)�������{�A�G���5����MW�+dl�n�M�����Y������h<����˝�t�l9Fm#�{�H��h�;�5�@5�A��'f�~۞�n�'�1�����y�P9�딙R4�VO-��ve�F����z���{B�J�U��Ǐ��r�P3.��N��*9}���c�R�tw"W@��X-�cW�DK=�ݟ.0���X��4���e�>��j�=Y��t(��F�^"��_b��V�Ƙ@KTy��L��2 ��(���ے����D�����F�k��Dt��f���u�W	����]q�1�4��n1*ǽQ��:9�:a����k����B�ѿ�{�W�"�pi����ݓ#:�=�$���#`���gs`�R�:�|��3�@���e˫�M�W�F�"�>����Kg�4�i���v��7]�]�]�.���4���S\�z=ZA`����}c�0��+_���v$�_o�V����g��I��侎�\��,����ԡ"�����E�j��t������A�3�_��mp���8O	�1�8��zX��`�.z�o��ʹ��4GX'���OW�*�j ��!Rm+/[Å����ףS:x>������(r��T�쐒�Pl4�ք7���I{�����.��$Zi������xs��n�Q����O�/�G��窛�lk�]Gz��ӥt�oM$?m�o�J�7
N�\O��Ӕ�&$S�H��z��0cׄ�7�^e(25M-��dd,��!sEx*�tZ�4ǌQ4��nuU�k�ܑu$݋��s�]�R7�� ���E���e��q��5I�-���Ȫ4���9��<�и�7x$��?5�V>�#@�Z�K�?�Oj#�寜R\��79w�_��gj�k[y�e��R�g� ~c�XC�'O�!8ٗq
��'%���+�-�:*m12�������N�i��>0gw,3IF�K�4Վ����	}�`�F�׋�����A����0Y�~�K�*�������\�� >�L���Cx}c5��6C��	�61�tw�:�Z@Y�X]o���u%��$���7o�֝�ʰ���H˼"w֭����9�l;��g�"�J�$�BI�u��Ƭ�g}����M�0��'�J�;z}�qbXڅDm��b�^% �F�K7d�b�͆P�O}�x�ؤ�0њ�~3(r*Dl�&:��M�A����I����$�dZ�dT�]~^R<#�{?�kJd�zVs��x6��t
uI�)��E�Q�����o�+��p~5G�� h-椋s���
%J<J{�X���l�ʨpl�[k�:"?%I$g���2�F?�s���`�m�Q1�s�	�U�TrQ�z= ��O��V���CC�!�E��C?)p�'�-�5���.>
���$Ӛv‼נ#]ȸ�Y��W��wY� >ʕC��N�k\���Nޙ��n��;%(D����$�9_jK"�a03 �@���\h/��t��0���;4���^�W���q�vt��_ӇC�I{ ���R�19�CG6ψ�D�س����Y�"M
�@r�IvI(�����E�J��+�^���"��e
q��zH8Y��hrRn�oe�\I3��;��*ٛ�2Q0��ٜR�����ՙ����T��C��� l(��m�&!�W$ q��O��J$�=_5u�kv�K̓��N��&Q�
v��~����h�//ל�אu_\��^%,]p����S�s����0�?�q��{�0R�ԯi�^Ǳ��X0�M|��S�����(�.nl:
���N؏P��n0F,�8�[;|���t�#��]�n��������.P_�g�#�j�M��;�'#2�\�$�^/Ir�C:X!S��&�+���-�&�����ܐ���
~�[�sGB�D`�ȧ�wƩ���n>7HKU��%����� 
/�'��ȡ;[�,���a������EMn���#�����q�[ �71hi��ʊ�)�΋X�^���7=��=�a�Kie�1]�j,�3D��lZ�9j�?l���\?d��l��M�v�OK�e�u�������>�9���K6_�{f����j���i�/��ʬ 1���c�c��~q=��͋֙�N��x۩uW�T�!�\��k��h"�]��}�x��,���
 ��Ƹa	o�L��1F�]��~2i_��§7]��-���N��{�ܲ�u��_�Jby�d�CG{4a�I�2�0�Kiw����xZ=�=�{HK�v�*j�5���$�����,�=�r��aa�5�4��!�0�uvQ����H�.�v�s��N"��Yzf��*�}D�yMP�\
�����r]�^���4���G�����BZ�X�RJ^!"{v�;� �:�5oM2��˦���6���;#\���MP���e���L��c�tL(�Ƈ6����7&�R$�=�q_�>D��h2mWŬ�V=T�����ڐ;�5���"���ou��}��(�H.�����SK��bP\ه��it��,z a����}�S%v���ԭk�NbR��#>-'�֟/E<:��L�ё�c%�%潮��T��h���?§=�]�L��'�ݹ	�&$��6������m��,ȉŸ�����2�٢�o�� ��[1=;+ǂ��j��5�������-sk�Y�J�WU<�*��|h��y��&4��v2v�ڲ�	��)�{�ְ����p���*r�)��a �(���^�j~��I%����f4����H�ֳ��1�A,è�2]��Ƞ��{Ǖ���(��v-:"o���΅�ȘL@�����?{��q�{r�FCdx�|A�FrHN9A�Bs�zPneN�"�j.AR�6��_#��`t���b��.m2��D=���r2�$�S�r� Q�}=�pK��y�}�����BR�Q�?
 �7��}�'�1�> `�!������7�L��8@t|`#:�z����G��>J���.�]ś�������4�� Ϸ����2���Mf�!�#�
Դ~��:��֭�QJOC�~ʝ���ҀK.����Q�`;C�������T��uَ0��"����ۼ�(���7M��h>��vG���W��)�������TL�$<��0�-w��ԭ��Y�.Kfc�m��xˏ���a�P�Af#cT'h�O-��D��#��N!�%|��|��<��g8��w�g:��U��

�*W�Gζ�h�qUڍQ*�|�0:�|��K+�U�o��2ԣ4�3�"�)-Ӑ��X�=ắ��uoub[/�_�%G�Dp.��AKܮ���U�bc�:�����UR+�F� �[�԰�<֢[N�o�̼k���^b��şd2K$ +Ǳ:�h�f�f1p[�`��&J]+#>V �"d���Y[h��E� C)�c�I�T��^C��B֩U�	�~N!m��@3v>,�h�Ws��Fml��O��t��i��]�Hb���;>�A��9c�A������/{:�Y��S`�O_ZA��2�ϡ}:\=�_�[��!0z_���|���Mܞ�����҄�KPh�?'!
X��{� ��p�����u	U�S|#�k����Ք¦���;t�@'F�ñx@4�oy}c��}� q��]'�#ӬO`/Iѱ�?�h�.���z�Q��v�5zը������Y�,㝜�ֵ.���w�C�-pڼ/8H �Z�3q켁��2��I���
.u�>�ԭ1J_�&�2�B��'��-@��jPq������Na3����D{�g�sdBq�N4�O=+�Q&dΩ�xb��uvAxQ\X[��j�!���\��eO{t>��%U.4�97d�)���Lڔv�Hz��p��ƭ�c$\d���?�I����d?m䵃�0��Su	1���#ϖ����ݵ7�o�> H���ȭ�x��h�.94����Fn�����9���c!O`y��܀�Ȗh�M�?���Nw��d��`�=��v+#�0�Y'�]R�Na/vB_N0|�Nvd�?��@ە|;!�Tk1�����?aږE��y��Wm� s,���q�DP��_���M�g��k����$��� Įx�����
��U��z�2���8�yq��#",0��o�J����#ȞE��ѵ�)8E��o�CH1� �)@�jp��%��K'��l�����m���m��˽��W��@�.!q���D�i41�`�=�[C�[Cy���R��a��|��i!�B�	h��^J���ͳ�	�TwܘsM��  O:����T��ʁ�����|���Ə���9]d��~�?�`�|,9�O����_�V���7҃*g/F�5��'Q�������� ��8�q��V>}�^.��G�� �6��g�x�C��kWł������5�%-H�~5<U�{����8k�m2�W���c�ĵ��O�mz��vP�XG1���+��a�lwJG�I%-�N��UGF��^�����=��O�&P���J�}�o��dZzw���R2�"QՅ�6_�W���G�6�;pQ�1�}{T�wZ�n����`/s�W.��V����(e���	L�<AVj��?#�rO�z��!����:/�e�~�� *u�$y���?����)���7�؈�RA�=U�[��%���1i��$�.���e�(�ď��o::F+Tm�(/�� 9n�@5�:����?@�>A;��.yz�|��:=��A���]>�pi�����O79; �Q+��l��O�B��O:��ee�W���Z��>�?!��8p��C�m�W�����r��=u���Zu�_�����œ�7�Ï��J1<x��-�/�ȍ@xxP�\�}>����C㔡�:��9:��1��~Y[��:�zW�ţ�4/SE��{����x��F!���N���/��<D�����U=!81��s�Aj��i�����  p�'��e[\���&�AC�}�j� ��aؔ��w��!�#-۔�6 ��IV��pzM���C�����$�^s4�L����we����_A��ĸ]�΅��_��6� �W&�7O+ؿӹZXtM��WlX��aJQz>�E�@Xl��A>���#?q����v眿_)mfd��\�u���9�VT6�b��i��\^�BH�T��{���O�ӷ�P���R�H�1�)���{�����E��t�ӕT��-�D_Y٠/N�������u��7�+����3[�(��H<�΍���%p~7;.�~w0���"�j�K�A�9�h�"�1�U�d�՘�JS�����a� )���X��w:A������<�0'�x�:kIDK���_"��d�Cg�Z$�����A�Br�u�bx}:%�ѕ_�.ƕe��u<fm�Jd7�~��H\���ذ�"7.{����g��f��J,���m��ֳ:Z���B7&�d���T���-��fэ�\:/�3��q,k �p躙���9��� V�7�C ��JF��)��a��BY������^� G=�f�1��#���y����i�6�����y�h,�nX��G�����+�Y�Ī�]�s��O��V�.�̂���)��{G@?��N����O��r��׻���Z3?�$�/���_yvޮg\�����ሔ�
�$b�X����s9�S�ك�3��}�t�2I�n��B�Oo~G��[�{�8��^_�O��7�&9_�<�1��_F���8�4/o
z�RNX�֒�~g(ҷ���#-�U���_pL:f|��,[˱�HH0|�| 
Mu��+����x:�J���g\��Y�0B��72�%���&U���1������h���笈�y�ݛ��cs`o�Oԧ�=����Upa�����/q^n!7	��Q������~S�K��[	�Aq����3�'��T�;Q�W��U��PTg_s=�Rű[}Gw��<��0R��*�eE�ۮa�9���r:`�-N�/��2�,���ޅ��W�������1�s ���e�V�B�N&��y�Ӕg���#�����>-k�F�î��H�ГH�zг�9��c8d�#�јAP�����Z�w�^Y_̆+%��Rh�}���#Ӊ�8bl��!Ѧ�e��ix�CO]��[�Y[�-��ع��a_ ��"2
, �x�
���fl��9^W�G�&��y4��eC�>�T��(��.r���.އt�/ik�� �'�����?�)��o��ӰX�]�q	���;؟d�� ��?�t� nH{l)�h�ђ��љh�t}G��DJ?�<N@J$,����O[�\�h��-����Dhֵパ�n���h��[�O���v�0�HI.��oe�z�h��g����S�C��c���Cn+Z�ЄX����U�������IB���WY��e�K�*RZ���~૑G8)Lz\!�DUN�Z��ZTՈ˂Ph��;��Q �Ɂ/�>�ы{)4s)~n��o	B�W��_�Y���.As"�	T�������^fZ�?��e�{ے�V��*� �p�y��l�~ʈ��R�m����0P�v���gO�	��sJkR岿��,N��v�?Ѱ]���oM��LM�<�s�}���R����^�O�����bێ�LNՠp�ô� [Ɓ����	�{f*�>���.�I��Xxm�Jc���:}��ŐxEs:��X��_/��x���w���VR��[�Sok�kTm䣅��D$ٵ��Ҡ�R��K��M��F��_;���ks�0-���$A�/!�X�U�F�;���y']�uaw��"�cl�g	�!����,��Ø��'qӞ7g�<�l����	�"q 2�.q����'�o�x�o|߸!������4������F�Wu�P�-x�^ハ�v�,�hjf�S%򡙆w���Z�à��6�8�P��t�����	5���Dj��������N����;�OIv�@Ԧ	��8�wX����Y���ە��%��b۬��JPR�1��J�e$!J�y�_A�c5��4c�8n���3�-���W�z�@[����[Ҋ�ڬ5M/����:[�����?�\��V>+�(�WokZ
���TnaP̐v(�;oP���斐�|xK��eH��
�|��%��O�. V��,�m��_�=��-���0�y���aS��xUv��#P��/�~���	7��%3mհ����0�{i[�"=�R⿻�e�P}�i�_
�K���0oVb��	SM��Xb}��@@�Ή��]��Ʀ3�_]��rs�ct��� G�E���x�]��U�ّ���}8cƅ�"C�!wtQ��b�iyـ=J�<��C��'I���.G���=(Us��ҋ�`n&Z_� �l�������<ξ�܌ � v�s���B����z�(U�xF��M�J�;�L�,Y�z�#����%�?P��[.��}vk�������3�'��b�A�u���'ۊ�:��;9.&2��^C �K��O���; ���i��?��e�,����(]l/��jYs9ycjV��B��zCt?>tּ��V�K���(�:�}��� ��ɏ��w��v2��_n_-}Y���>��m���K�Ӫ0 �7�*:H���$
F���gO�(���zV?�}ͬJV"��'�~t�?�uNZ߾r�RpRi`����q�;�ß�BT���U+��`�P$���M$��,`ᖓ�S����Ǽ����5��4�	�!:����z�<��	�/�V�.hh���K�����2G��l �:Z�4
ʒ�UB��O��j{#�(|��u>�������`��U�|���e*Yk�:����<��<�qr��m@J�9C�w����C$�^2B����R���Oey��lEkK"�g�T4�&�ǧ�ڵ�s-����u��t#�`��%�v��Iyw��+�x���h�0(p���'�ʹ�k��ҏ��Q4a����,ܧc��ꀔ�qS 6O�H�\B���xf������Erw#��1�p�?��z�&��J���n�ڟ�厇��D��v�2���;���`�q��\��9�rWM�^�70r1RPm�0S?1���\�MN���LB�ץq��Ptx����ފr)/T�)�s�?	��q��*��R�b���w��f�����+fko(��Z��R�p���J^�h[0���K���i�S�TQ�� ߗ�N"ѩE}��H4d�W��Z�UA��Q�%՚���~�<ꈤ���OP�O��2�v�Z���1�v������֪J-+Э�
��xu2 �1J,�+%����O��p�픗�+?5�����P/�!��L�R�um�V�b����m'/CFi��\:e?��"D@��ޭ�Ϊ�Ie����M���C�[k��fnߣ�7^��^^]��:��_I��\���s�F���!�a ��lu�V@D9)桹,&��f���?��hC�Ӆu�\�}z���\�ql�#d���*R�Ui �|����Clu��cu��j��/��0��B�z�S�G(�y�u$}N��S��N.%�Z�����,ܭ��m���>ѕ��Z�����գ��oe�Z4���h,3@��eތ��/Cg��C�aT��Q���$�w�p�>�l�	đ��:����ڥq�Sv#C�un*�pKJ\u�:8;Nu}57aΛȬ9l�y`ѳG�p7g���6B&?%v�>.���fU����ɗ��XC.Z���q��*U��z��z��ܤ��L�h��������2��3��E�������>D���z���cL��E�\�����R6�G����V�=�~Q>2yW{۝�;"�q哵�..�A�75_���%�Ezf[��w?�o���y�k�����Hcu̶)�E;y-��ަPoL�6�R���r���п��
;	���8��5�Y�#CZp����Kg5
%ތ%E�]6.�l��͕_+H(7��JW�+���%��:�S���5��x����dk��I(���&�R�dY˳���9j`7K)�_���u]:\���S���A6�Q&��!3I�a�iI8��=l��>��6�8C�Qk�=p��sp�̟���r�ũ�B:���k����הl"���E��<-,�:\P�NF@:�U"	�^r��K_C��7�\�a��倏
ūb2���dh|�x�������SO�@(_!a���e���r6ʠ��-�8�y�����̗���&(��
�~��r��0T�-�z��61]�s�k 	C�y��&Â0�p�e��
L[��ک�����r%}�a�nk��]˱Oi��J�#!���{W~T�W����ҷp�0i��v�����Y�4ғm����m ��ϥ3�n���}�q�� '�M]C��w�T!9�c�J���T@�Q:p��������H0E��?p6P���#�N*��j�E��!���5�n�n_�(��h����X#��i3�Lj$Ι��t��ne*� �)���`���I�Je�s��.��E�3
l�E�Z�.6���-���Z�����<`{�7�Zu�)�T	2.�'A8����"����#]��fr�E�&�Om���]�2e��hJ,S� "�|$���c����H���[0LW�	#^N4� ܭ�b�2����p�>����i� �ܫ��t�O�<覾��A���0i���J���q�Q��?���M�f�V��s�Yw��Lw;�IO��zG�I���9GƤ����a��e ����Z��yE �T��xz��~<	C�(=��9?ˠ�&�(�^�̛G��Q���)�E��r�К�B+�*�R�[/�&ٷn�&�m*���|]]��h�l��.3t[�O
2�(�y����qD`�o���[Mt���ܟ����E'��0ă�Ȗȅӱ�X�����Bv-K\�����J�2���0]"�O��z�E+[����B]C��(DD���YH�V2�ђ��Gd0 c�L�.N�כ�Tٕ��}e�Ex����T8�w�R%����z*�f��9
��٤��a:�4���H�c+��c�5mܝ�~(�g��j�������y�M�r�@3�M���@�����6�7�m
�c�_"�fq��;S���^W�D����žx��q�w
��b\,��(|=�{`�����S7m�90]�b<�2�*��z҄Q7��.[�&eʠ����ǯ��<r�$�!��X+ $�o7�ܼ��z��o�sش� \{�zV�#��~,nIfÂ0^�
E���7�j)�B+�!N�i���K�4��d�	���⾊ox����J�i���3ݒhsJ�s5����5�Σ�g�9�𥉉�a�;���f�i�-_�9�|4!;]4�K�]gF�ٺ`��~	��fE���m�y�����T��pO�W�$�kw����,���R��a*En���-Q�W�ŖTI�<հ�����8��M=�ւ��j{ڈ��:Y�-�[ǭF���\�S�AAZ(�����	k%��x��6��"3G��]h�,�$��o6����2�0&�3u�Kă���C��Q����y0o��'�_q�@�!���⒛RR;N[
o?�8�X�/��x(����s����QV�F�����_Jk�!���Q7� T���ut�vCd�(�3q�s�Dh�*�c�د@��OO�Š'J\,t���d�׮!�|�w��-	�>��0\�Z2��y^.	�8¢�C��1~;��PZ�F�8�����������$��6��E}K0)�l�џ4E���\���a����ЛW�/�pK���Id _-V]�7�4R?0)����	$�ͬ�)3��s�ؠ�RХۓ|��#����}�\Gjt�^���n0��Gٳ?`9=��烪T��F -;����IB��W��G򫒢Y���u���;	��!�z�	#P�����]��);x{2��K�
vT��)?yzi���>����X�����2�B7e�U���H�#F�>t��)?�)��M)}JE}n�<	���u%ƙj�}��nf$@n���
�W��f{t G�����e��+�`�In��C2�:����7�)ߟU�7t��h����#<�&�O�*G֨`�ˎ�L�>|�1�����OL:e�����`Y	<��cb���,�%%�Y��y�����/xبn�3��{�/߬|��[᥷�!�tk�0�)gA��]�xD���[�Yˋ��m9⠛�➅��_2��٥�m+E��]����#��������]��`]����X���D�T�����2�t��f,���u{W�u��Tw
�?�y�K�F�ej?�	S��w�6�C�����!i�C�-!�O|I�	Y�{�O����z@ ��/I�ku*ϙ#��pɒS��ψ�nX+�o}E�om$R��zlt�E� ����g�4	�)��BZ��Q��4N��D]�X�fQ}�2��)�f�Í��\{<}�8;��o��}���a�3�R�'��NC��y��DYK��3�c�F�ǔA�Qj>�ܪ��}ESԉ���QUCT�/�V3P1�����hp�!o�Z����)�bRW�a�����o�����8�{�W[���?����`{Uq�!d�lYue�vתDK%��%�H�ڃ���_�@%�L'�}ܝl���`
�}հ ��_�Զ\�}�g�9�7������`��2A���P#�l�@�8\����^Ċ)�f�-��L�SD��z�ý֍��c�'�����8/;#i����j($���ܳ�(�|�^�������Q(�9m���`sJ�0��1�E��A�P�{�sp��o����VT�g���IBS\k���'�C�s�� ��a��.:tQBI�QK՝�_䠒ؒc�[�n�v_�)dL�.�Ϡ�,��ʽn�Ѳ�U����a�z�R�d���<m�ד�����<��_<���7���'�����Ͳ������;.�E"=�'!�T�: ���4pj�������؇��\� s�gk�z˺`����n�hwZ�̊����r-ᢗ�F�D��P�ꟚY���׌��]�}p[�̪��EГ� {�{�è��m����� ����s��h��c� �3ǀ�a6'�錘���������c��BlQw�� yU��(�VQ���D�0c1�TEf��� �Ǩ�F��*/p99���MZ�4��,��o�F���`4Rra0Ԇ!���>�A�N������]��3��k�ʱ !MV�0�O��e��ӹd�������PM�F�aP�?lQ���.�����t��&1����z��C`]�����@����j��ڛ�T�|	� ס��&����e��O'���"�g�B��o
pY<�D�o��W�U�:,�B�	�#�p����$#-��p�g$�����h&NH��a��ئ#��x�+�"b�8q]���H��0��\]�@��9+�	L|&j�%��aj����a/��|m�������_H��'�*-��Y0��d�'����[��M��]��rE����e���L-Rڔ�� �����@��2� ������?oV�.�h+6��j{{�D���/4  x[_��t�%�UDZ]͞�D���b-�9y���W����唐��ba��L��m��,���:W]XF�u��~���wX{�>�����Ea�kx�s�M��E,�ia�YJ�r)��LY�WI��s�\��p���W�EZM�$�p�����uU�A�4T$��B���]��tq.A�����Y��D,\iF	�I܆q[�y~�e*��_1[���2>�ԥQ
�q���e�?��'V]������<����.*#�3�2���@zVg��ŭ�t`#�;��Ԁ�Wbf�8�$�3Aaam�������R�F?������i���u��T�^+
���Qҹ��3+T �]|{�$f8K�	Cv#�#�Ћ�w�P���ֺٟ�U���Yc$�WSۑrKh�fn��R� ���ez�B�}=�3vZ� t_����\��|hxw̹K#��P|=b>����fnZ���bY�-~ �'"J���΋Kit�L����O]��ܩm�)�l��c���!���b&{v6kk6�	㏨"f6�y����T`C�HY�c=�O��x2"+m�8^{�Νr��Vx����|�s��X 4��K"E�����N���˿aN� ���n'U��䃟{I*�Ro~E�ю?�����M��z>�+$��< ߉��#�p�$_Ժ����N���[�M��N��}��	��h���LJ�@�/N~���Qėj�����Q��D��)���}����(V����KA���-n�D����=Ig���(Y�j�GMWa�(�_��*���v����7��rE��ݝǹĒ�X���$T'kA�$�tYF��Qs���Ӳ[�i1Й9Ǟ�̀i�7]紭�!��sU�/�f��S�D�8N>���J��ʷ�_\�^��
��a8>u!|��l�y*Rh��cB�)�XU�S�����C���'l�IFj��Gc�J9��^�����s������Zo7��"�������g���bx��f|Г 6ձ�G�>4��ȘS�65��F��D��	z��oӥ���z�;�9���|�� �a�G� �j�b�ho����5�h�ː��b�Ħ����Q�~&�6]�)H[��
��`�2��^k8+Wo���8�H��z[BY(4T��A���8R����"׸N�=�Ltu�:<�|����b ~:�
Q8�k�>���Y��<�6LdE��oZn�kK��&}��f�v�2�L%���g�F�*	X�T_zt���z(^�Ҽ�o��=�"n�A�rD�Bp��>	�~1�|QI;��&��*��*��^��>�t��h܄�T�]�K��]jk#'�E�U�d��W5��p�ky�t�1��M�o\B�U�]��u<�3���AR�@f?q�B�2w�g�������D����j^6���o����ʽDC�A�&�hg��%�;<�ȳ�A~<���Xncֈfg��'h�ť"�?��{��EՀ�̜���Y�z;�Gu�8f*�.K�����<B�
����l�1�r�s�Gd0��F��K$�78�Mx��U��f�7���(G׶�<�R��{��7�z@�[�xp�ڎ���<ȷ-��E��%��f)I4Ϫ�7<��u�S�<mG;aG��.uK��fs<��K�~<�pDo��f���:�~�T(z5COkc'E����$��ش6��mj�{��qj�R�XM
a�.��?n�&�c����݊��>N�;�����2�(nQ����V	�׏��8˭'�=�J#r�(:�0�u,�'� 1��� �`^͓��?��i��j��U��M��O�QVh=�[�����J�S�U�4�w� ru�E>���ܢ �KCx�����M��!���j�R/��l�9�k)�dEU�S�,Yvh+i@ǲ�qZ<yYnq����0��m?(Ov���b�?9bҰ���N�&�0���G�k!�����W��р���c�KZ�ѕE)�K��9���K�"�7��������I�- �*���_�C�P�#��H����,�'<�@�B[s��������a�1I����ր��8�҈(�0�l�sюϘ��׀e�l^�����l�	���նq�Y4��,��=+��Ŀ�f�!�9��s��_l�Jl�8�B���[�W�նTt����ͮ��8@�˓=�F.Bl�F�`W�8fJTS8��)+ ���%������>^���b�J%[C�����?����R�kr;��`y	|R^1���fګ�"�B1�b�(��)4��J�a����W��؍x�p5;9	74|gx��������7F0�)Qb;�u�����J�@Lc��ߦ��Vt	x��SE�ó�D!�+��M܌u|T�&6�>�!C��iV�/1n]S�HJ�^Wt�,��Sn:�e�-�n��Xbɞ�G��p�QoZ,1��=aXA�XK.�0����x��)�nP���=1[[��Vk`�\�|�����V0K뉕�.�w�7?�s����(�X�2�4T��gHW>�������5\�M&}�� #��=|�*T��c�*�B� �ش�s�WV�[K?����|��|ӳ#%\��f�y<0V�$����
L�H(+�b��y��Z�ת�f�x2�!;W�ޮ�n<���0n�Z�ⴢj��� +��m�i����q.��GB�ğ*�϶��\m�[�P׆^x���*,�d�b,�R�x ��v|Y~����V��jp�u�VE�[
�b�X�6�P~�F��;�V`�N!ԏ�^�α��3g2\S��c	���o�x��V�N�DK�,A
+�K)H�O�2a�m�q��B>�3�{���f�sg������]!mc1��O�`C���I�+�'7���Aa���5
>HI�D�'b��ߝt�慇"2���f`�T��jep&<�T.NB%?�	�e}��p��H��_Y���p��J���ML���i�	-8N�R�:�]}�5\�H���3u��R����S�\�N��_��<��~9|(�/�'>�dy�`�;��X��0rЀU�Z���bOtz��s����&��[[�}ܣyG�
�4wF:���̀�5�T�}0�h�Hx�B:��+Օ�
�e�bV�H����?�4�RC!Kf��u�(#�P-�����OZ)bmt�0�^;�N�oA���_���I<�ՠ���#T�?�vI9�mI��?vRa]R/W0�py�=�V'!|I���7D/H�K:\�|\�ޕ����qb�vB)FkR�����~�&#�`5-ß`9gh�;m5֧of?~�Ѫ���+�;�ʆ�!��:�>����;1Nm<�s2�@fP�{xUF����c����S�0Z݈���Y�p��C�i�+��-�䨟Y�tx�?���B�*U��i�x��P�aj��fg���剜%eR�j5��̏�VrI�ʯ@bi���)x~�e��.��kOrL��SY�J��Ӓz�ʼ+�	�1.����F��L��Qi����S@!WQ�D%!2�%`�gf�3n����O�%)%�Y�<i� �r�@Re	m�B&,�9v�"JN��܃��"y�)�����Oh�x!N���o�C�PH���<5X��v��6�Gy;d�Xdmef��vӻ��.�ؖviX�(^�w#��*2�ă�H�=����v� ۃr��{QJ�՘8�ռ:�n'yf�7��6z�~E���;seM�5L�p(z�gB�
VP(�>�������d=i���y'��A����@t���9��e�wP�JV�iHW2a[y�C�1y.\�"�[v>P�:�қB�r��N�L�[�9�����Ɖ�ya�����
������s�Je#
fC���H�}Q���d�t}��r���'LO�P9�����	bS�'�ʏ�^K3^�����yef)-��v�+�j�x���D�Je/�i.���be��Ni�OοS���h�������o��]+�M�ӢH�������|N��m�����J��B�N���}�*��#W3W�8�>F�0����KUC���L��$��a�.��7!l�QW�����*�`�F ��P���gO<Š��Nj��8h2n��ԉ<jF6-pd���ѕa�E��X�[Lӭ "��7��cz���U#ѵ3](*|�B ��3���cO��;T �P�!U���m��W)��ӯ٪�E�S{f���D�H��I=8d(0x�б�Ĩ: K�$�C���`��T^H0�����kgN�h��t� 
	R¾�W��=|�΋z[B��D��\���bK*��?�d��Cқ��whF@
�5��,}L��P��}4zT���4<�����<?Wk���ԑj�x�^TN޺��.io�\�P����fV�"��5�49�D�/�2Ǎ������
�&�)%ƅ��7��>��7!oT�>S+����=X�l[��52x����a���qA@�A�lϚ�y�/J�L�q[��晙[�INHU��b\y;�KI���/��|�	r�T�)��	��&�~,�n/+��	�h{x��	�n�zL%�l��j������HS>��)�, �or��R�ݯ_ٌ������2Q��A,���^�p�⋋$bC�	���0.���
��h�l�Ԁ3�v���yl�? ��_�
����M��������t�m  �㤑^r�����j�S h�ٕ��<�#�N0=�1E��-7����U�?F1��ʼO�ň{��0s��I����T�f�@C��\g��S"�rڡ�`h��X��ك�Σ�&G�*h��{p�`�37��<������_%gÐ��9��r�s3}�ܲ'fHD���U�d:N$|2�;�xX���Oaˆhmr2q	���YK�&���Q�Z(�xsWؿ+���U�
�@{��7�ឧ��:�B���8>���x�̼"�dcCO�xh�����6��a�B����X�'a6
@�ٹ�����Ft(ʐ�$��`�8��Ѵ����s_	���6E��d7:p��3f%��(��a����bT��k��s'�*/�>�̓����_�.�{��Z4�S/�d�z#�a�LNPo��4+P&�W�ˤ�"X��w��i.�ٻ�.n���NdZ+�J?#���%�+A9���Og_���[����U���<�7G���V��P�U���؞����3䖮�m��Lq_�T���]&���%H���Ϧ�9��<ԴE�ކ	��dz��E2Sh�T>�|�C�5���$���j&x�u70�*��P��t=q���	Q�!���=X҉�W�~BR�e'���Z��+�dV��#��O�5`�~.�v��K���8{@�@�	��y�bY��^D޺�(qo�+���]dj扴Q�F���v+����W{��'�T�9����q�Ih�\��]t�|��(��g	���hd-��#�hC��
� 5���\��.kUL����GӺc��@\�a��Oe��M�*'2�@tTL�6��:�C�N��C��=�'F~���՟�Kż��j����?�0r\�JԤ��t* �� ��c0��rDQRY�qO�Rˊu��9?�w�'�fm�P8�)�_��	�U�p/J{�|vN7}��g��xE�>ޞš��:�1��+}���V��1��<��+�6^��kq��~�kf��6�>�W��4�����h�)_\;&ś�ڬ� �u���e�'��ȧ��O��"�A��6C0U�~Ł��s��ܐ� m���B#�3��gՂ�N*�Ԥ!�W�4���e�z��},}m'�����-���^KlY�ٕ����g㈓�Y�3�����u��EV��:���:��l�/����@�����2��T����x�C�83ɲr"���Ju-�g� X,�/i#a�]s6��C���W�y~ֻ�>Z�|�$v���tk��b��+��.��mC �$ΰ_�����,d�(iv��kY����Z8L�0���7�v��Ew�"�D*>�ǝ����N��1�n����Br��x |o��
'�:��+�V����.����9�R0MVa�{�	#w3K[�`{J(��-���u��ǫ0ǋ2�O�����/�R+������/XNq��2�i2RP��!��6|/p���[%�lE���f�{�����*ː�O��[v�<��dk�%sC�~s��5�o�-O�TL{�x�q7]��0:a�̀+lN��2�[�{̎��n&�~�0�
���ƭ߽G'3�����z��#�c6��=�{8�ܒ5x,�U�2��s�?�C��v������!�_���,����<��(�÷愑���P����I��*�*�B��1Q�t��T��K[* .����OAv6g��O�d�:S܌�G�59��P�`�W�/<���9��H��ý�6AeM��ck�h�"gP��*�6A�Y���JO^��#z���}�{`'�o��]��\�7�a4���'�n�|M�����5��ŗFY��\,V�^V�I��	yI��e���������xy�hJd�J�kR��g�``��8_h?��兙�o4;����	]�Pw���9�?�e�'���8wW�C�O	$$ �%���Z�}@�G�s��)B�mg�iS�,�ur��ERݰM�����$)+�ü�Z��˱F��S��l�������z«R�
i�H�r��	�f�%ۥ��s5�jVl��f�*��9��bhF���;���?�T��}��5f
U���xu3!4������S�����{WŢ����Ó�r�wS|�gӜ�K�[gBe�}$�����B�ƼT���ŧv���\�<ƖXu��:�q���
�j�2[�q�r�.pqk�z�s�C��|�s?�W����z݄ �l5��t������T��=u�z��G��<����n���I�Z5��[�_LHf�Uʲ=���H��"��+��ܥvU��N<A��C�d�؆J�Y�
�h�gV��`���6�<�q*�`a]H ?�×�G���G�G�gJ�&��
)�2�7L�xfN�"˝X�e-��[�@�NKE����d���5���ix�����V�x�]�I�E�EO髳.f;wc���W�s�.�S���� %���ps���j����fm@w$�}�j1�O�)Z�P�}>��G��(}��J�t�pv��0c��U����O�{"�yH�m�?R�Og��`��Ɔ�K$�a3?Ovpw�h�@��h���9�-�NM�]��i�A�
�ڜ��3'[��Z��)F��GI�s��������[��:���~�.�7GbK�IHd�."�d"zT8�==?��ZU����c� ��u+�w7��������OTn�ԩ�aI)�n���z,�8J$��n�u0�.��%Y�_�������O��pS\jP���:=�0b���ޗ��L�� (�XYn�%c٭�^����4��ꮦ�%B�p$�h�>$��5:����"�4Z��A�$����Z\��m��5̴B�fXM���� �j�$B�]n%���O�~��P�kis�%&��.V�3����4�7�
��ެ�2�H��O$����W��~}�:ݰ�С# I7|�̩.y��Y�$Q	[ ���P�t*�\�yc����������6
���d.��u�C��g�K9'�(x����c�z��`�h_�8p���$�Z0 �Z�7��b��A�c_�� �&���&]8�E�Ϩ ��ٽK�����C���y�o���q�C)��_#d�^�췡��	
�퉴��,j� ~�I�W�+6�ў�i>��Qh���SB,�p0��xdU��� f�x3�Ɍ/(�z��~R�%ס^o��\ބ0 }-���Lo�\�"���-��k|�^��ċ�����Tt�C��2"҇����^2p��?��f��}:T��F�,g��ZrY�W���xX+�*�\�mY7ʟ�����8�����o�k�	5΅<�l���
6=@D�뼵Ӷ܌ G�E�E��|RW+ٵCU�M9����R�	Rk�"���a�R��/9�@�!���z��S�R�Q5�$�&�q����}?�b��[�f�J�w��Fqˮ���>	L�&�FK6(���?%�6�M1=i��P��)f^?���5�p��ӝס�b�����i�Om;�������J�]�<8����9�_E;�}'������D@"�KAT����aן�b���ݸ=��:�4z����>�ͬ.�^�2Z��Sy�ݰ�̹^zTY�� $�$�|��Ξ�NP� �k��ڌ���QTE˥�X�g�b��y@23A���Ց�k�nkl��3�f�><�pV��F��
Y���+�ȡ.�!g�D�PTJ��W�#;;����Wn��엾�ՠ\�����{�~�6�h�8AA�7;bQ�?�Wr2��f�$�����P�M���Yy}�z��oӚ+-1�_���#[7m�`*?�J�����?4]���я]B� \��:��
 L�1��:���^P+��5���#�M%���d���H��V��:�jmz\�w��~�{.e�=�7Iz	}/�Z��X�A�S�M�3}�V?L���
���r�%��m�7TB��eXI,��ه&{�ʽL��^(���f���'�P�p��HƝ��&��}~r�x&�И���L��_rĠM����}^��g6��8�'xg��b�Ԯ3�?��!ۖ����mvu���X{D�=�:H��ā��ǽ�L+p彦�h�ρ��Д;�^(}�����]�Dm��O�.l0�g0��'�"�Zj��f9]�4��>J��E]	�����%~��DM�A�dq�,7�|l45(2��R���C���Y��?��v�q��/{
U���z%VR�W���v���A�P�٠����,���.BD>
:��^�8i�cn������v���՚�S��ӳ�B��!��;}Q���f��-l�'�g
�US�1��&�%O{`^����B�	�*�!�d8T�;����8�F#z��cP�#C����{��JЩ8�B��RG����+�j4�CHU�RSH�5=:���8��4˅k�p��c��{�<?�ͳ+����R��-r8�V�`xU$-+.|5fS�-��v�v2H?df�g�����G�� Jf�6��2��5|�l�W5�'*�L5�d��i:�ݢS��D]�t8:���0$fM�90H�hTɕ���2�[o�</�c��?���s�b�WoW�}uO~�vW����"���!�^�K�\��9G�6b��?s �_"�els�# <�|�{Q����C��n�
�R��3��ai#c)-�W�#���d��d�ƚ�!}��1��`S3�L���P�@p�5�K�C�oÆ_dO��ѡ�r�{�6����}�ڗ��)2������UF}ks�.���Y���%�8�r=V�8����_��D{��8I����~u\�ǒZ��ؘo��2���Ď�a�\+~/��l�ѯX���<�b/�-J�I3�ذ����%9�ϛ�(����/�EV���j��嵊R�&�:��z�V�s�܋l(=K�g��x��x��̎�u8�-��m�H��`�h���9<��m����׍Fp�w�t�����&�o��"_��PSZ��'E�Pu}�c[��vXWGeR��#����.��P?��ޟ�S&\;5��G���c�? ���D�J�ʗD���|�'S%M��6�M�E�Az���q'z�1�K�~Mz '��K�U��r���g�?�&���ok5�8��c2ĿG�m*�_zS���(��z	� �Ld7Fr���)�D��'�z<��hz5	���8�,ܸ0�;��Ȭ��OT-L���sf^�B
[ݔ<LG9��F�f9��
��ZmKdDK�f_Z$P#Xr�Zʁ�}y�.�Q؉Bqb��~nfO�\'}�A����9�T��j*� q��F5 <�G6y^0?�9�^]�ؼ&,3��o����$S�ܿ�!}��
r��Uf����O}X�cFGիD�PaTL)�����#���'`Qa���	���fE]�)���%�M�D4���p󺂰�|HMՙ���o�cT:��#�sR��Bt���M!ń�#q����B���$yho����mg*�;9C����s����)!&r�f�#�fmɈ:��K)��2h�V��P�&��MϤe�-����:�����E3���JA;��=�H.�fb���-���i`G�Z+sQ�s�(���/~P(��ak���F�#cW�ge�i ��Ϲ��r�F6�鴦��{/ږ!��
mݍdi�̍>��A��m��|s?Ψ#�HƯr`$f\����yf6ח߲�����8j`��{�Й���M�p!��� �o�v���������0��H"�yK��*��_\�HP�Ա� �*�9p�6j��DYrԈu;փv�p,��P9SI_J�L A��5�8�iq34���KĴr;):�DO��r� }m���_�P$�9�����j���B���6��?��[ fTZ���p�D&�(sA�Z�'�s�&b�ϲ�֮�C�#�sK��1Fc(���45d�ڈ�Ḷ��S�#�m+F��iі�+�hJ_=��Qͪj6�K�]Za������dG��}�k,f�S���-__O�����%���a�Bx8d��~��:=��_�g\�+�O "��������Dj;6�����/�b?|G/YN��i�� �%����[|���JL�`b�$�]�Bz��F6�8�ǌŴ�؆�&���I��N���%j�L=YT���$�ҷ=w�yZ�z`��|�"? (�4�5�KK�����д�#.Xa��%�U���@�b��*gݶ�����s���>��
�@(�'�
(��*�dT��U1Ԝ�C���>C�+K��A�m�S�@�n0y��^h^�rH{_�F/��i�8G
?#��9�{�;��ڻ10�bU@""~/A�Rz!��8`瑚�{:���� j�P�:��0z^���s��OU��HZp\P�W�⧉����M�����lyˀ���E6�T΂[/��ty�\��PJ'<�բ��R�ж��:��q��٭rT(�������O�8���}P��ģ'�,�n�zU��IF�繦��7��ؾ����O&=QZQ�=w�J��9U"�Ʊ���=�Ī��� �$+6��T��AXv��s�i�9�_v�֑O�y�G��n��l�zl��vw5��3��/�9C���7�@ۨ�0o�.	C̎,z+ש-��=2,��<�͐�Ɓ�q@��Zq9��	�}�ȏ����}O/��&so"��/�]�rM���kX�j7:��Q�S�]�O��Ka���P����} �D�$E�ϴ��ýzEc;?T�Řz�V"�ݝ *����G���Jč��w�Aj�+N�4cM\�[�Ѥu4IJ4����v䎦Dac�˘]�V�X�tj�,@��e�q  W(���(y��o��G|����s����/�t�c�*�V�r2ą�؇���d �ˇ�Y�:�M��\?�;j���P7)� r�yf�A�{'s(7y��0I	�)50 �[�Q<^u�-��O�h��_��.�M�z7�R/3O��h9�B�Lg8����K�܈4(E���|��4�=��	``?n���.ڬ'�P&X:L��M�����6�K����O���~�eG��-�D��u�6K�}���B�o�K!/&I6��8��c�������M�C�^�p�+}��oD��V��`����كOX-���m�2�Өa����Ƃi���y����@��T{GE�f��^�s��"����Țܔh�?#Ow��-�P�>]2imj��0S�BTW�����gQs�H���B��d�&��YZ�$b�*%�]�=�"�JF!�&� �����;d����¢�W~��dw�]o�a�X�E��y4gb�����̯��S������N�C��G���J��E�/?щş�>����*+�heWy��t�b���=��~��͌���NKd^-�@e�ۧY�'J6 6?ɥ��K)�+<�̂G`����nA�c	�t��B9%�9PH���j��B<�!g�����"�ܱ�j����-qe)��������\�: x1>�${��3��`��#O,�%�K��Jl]P^+q:7�}��J��ŏ(��:庈'�8��{a+'z���9c{z!p�.m"�<7�qS26+x֨���+�	��E��l���wW!�${����7&�̃N}���х~����Q8�è�^&�0Wپ*�=���T�$M����p�,U�RD_,��"3@���i�-�.�w��|E���j�*ks;G���S������S��)'j�{j�j,e����J�?�Ѯ�,
��֢�S���{e	k�ǡT7�?�����QL��l*��X�8��Rކ������+m"�`C4���龈e�����w���r�cL#�&�^�R�O$[�K��7Y �#qW����O�Y)��E�����	޳!t�FV�9�Y��3��2M�����Kh�����n5�2������˕�vd K�"��B��G�[�%H���6�,R���f4�.��F��p�KUM �g�0�_�=%K�!I��Z��_ �N�N.uJ�������ckt"!>���n<�k�2~�I3:xi�n�~r��$]UB�n��C�CyG`�	�����Me \�p?�|�k:�o��+眐�D�P�F�QGk��P��� �C�Q ��lG�7:
pc�#0�93vb�ז��
��[��8���z�8P^�~��z�z���ϖ#o}�b�ÕRYL�8t�<)�r�#E�)�#R��*w�J�IK݂�I�A*�N.	��������LA�)��0{P�T
jh���8ԙZG?��芇NQ����D��e�S�)���pM��5A��n�i���-fa��z0V�\M�^)��͛����܍��G�IM�Ә�(�_�n�V�jz�.��v�'��L�XV�݁�8������=��cN���|S-���zހW��ti�Idq^+0[*`����e�? ��o?ƌ?�ٿ��Z�Qg1/�2��G�3(Q����3�I��.a�	������PB����Q֜�ܦi1�e@^k�z^%y�����#��l�G�	�'�h"�ѱ���C+�瓿f/^s�u�����`;"A�F��D��1����Z�o\`�, �SM|C�'���@�����̠������D�v��I�1�Q�[0��<��kw�q���F8�זhuvr �b��-]fd���	8 ��0.c83��(u��������}��aΪ�t���x��[�r1U�����N"K�iEI�ތSA�jR7o��2�x�x�]�[!��PX��:"��r0gRQ�[�B�����	B6dS����H�������J]��g-���;��j)�������[�=!�	#�hA �]�:Q:mɘ�*ƱO�q��2>o�>V	�8}~6�����TR�W��pه�|߽��2�Ri��m;^zf#L���uH��^�:��ݮ��6K�9�;-=�ȕM�{^ͨ��茫�v��r���/����� �-�g]����X�D+�K�z�UyKk��5��3W���|����3ہv`�K���� �/�����F������)K2�=�[���'���SO��1 �s��*�=!!�G�r.��j8r��^EX�wm��QΣ1Fm��*.Oёg5�x�����d���ٜ^@KJ�= �v講����pm��~Շ�ͦ�ؐ@�	�KJ)����l���B�O{9��Ҧ,1a��� O~�A�]��dxc�@"�󈴔��Џ��;�Kǳ} �)Qc�>��I��� *=�@|����B���� ��8���ºJ�`�\��#��;����Fn<1�I;gq�	���s���y�ں]��^ϩ6��gn3
���%02��*�
TƁ"�E>:MpGo,��D�������3��E�t�x�6H��c�[*Z���fM���sk���ZJ2��5�IP�۳@k~�B�:���ܴ������#��t%( i�u�fp�ӑ�1K���v:�^Ma�y"���눯�Chj�Z��K��tJ�	ԥ�Y�;kzM[_d�}e��|��o��獖s���YO�΃�g������
�27_!�/� ��y���ݿ� ��^9ZPI1��zpc�]�o1A�?}�+q��uC}�����<x<Dד����7 l3������+.4�/�!iW�i��2K�}ʡg)�Z=�� gb�/i�+�s�1�G{�] �ʪ�"NX,����ocҟڝ4N�)T�n�:o�k5�Z(S�ؙ�/)�x� l�Gnd-�7����bb}ک-}Eꯍ��=E�R�gr=�C��0�4u�:�J�:"f���Z\�첟d���i���K�*���3(�O��w���ژ`KQ��9�Ѳ�$�e���Yn�0�\[s�R�ٞ��&�(�s�C��U�_����]G��2�ؿ�q����a��Y�o�_���-M>H��#��k2�#D�p�_����f���ޟ;��޲�۾�RA ���"|+,���L�X�`&��RüǑ�s�r�N���G�qN�l�%�f��r��vz�����g�t����bW�6�?�|XNB
�ߥ|�#��Ώ*%Lۏâ�,��R�v6�k��K����x�F0
�#Ms5S�,������DR�+�Gݑ�S~Q���,W9e���t�{�~b��$��1Y��T���P�LyNW6�������T^/ �� f�#���*yY�(��� �`^a�Ǯ��hli�f���`I�Y��M�!����|]}�w�D��}�-�d�x�ۤ����L����}_�Hc�8]K���=�4/ KgՂ�g��W:M����F97�Nv-ᐧvD���P95z�#[��=�N��b��f�Ċ�m�,�� �v�d,�w�rlZ���#9]1��hI�\���b��2��U�>��m�<:�د�Z�ob���;WD��F߻;�};��+9S*�Ŕ��QP�ǘ�Bj��������78vF�lEq��fm��رf���]S}��+gAd�;��`���`I��#v��b�[�\]���%S0(�!��qe˫�+��M�����l ]z20l9�cE�*҅��7�4���i�y)�Vr���*�X�@����Y&�NB"K<y���RCr��B�Ő�[�~$^�V�g��H7�HE��d\�{�7b�lV �5��ޮjp��g�7>��x �6�;C�e2%��g�2rl�I�D/�E� �8����X�/�g�x�j�f��������K��=�f���a�zEkܹ�:�|(��+"��S�yr7�AG�\�U��^_��Hf�*~���ύ>GE��ӂ��`�x�Ȳ����X��x�<��[|����/�c��z�C�d~co`Ğ8j�����+�<k-��'lf��C�d�Hr�T6��ǕX@�uT^f��c���;]w�;N4X�_��I��5Ɲ˳TP�� ���a�#we�6ٴ��n�P��;��A�J,���KOj��glhpY� ̵,,C��b�E<��������\e��4M=|+V�1��*�z�g��>N>AP�ZG=n�s�,���t�N���+�45^�0MJ���R���+�/��aT�3���@�T���y�NA��+�i����3���1�n��d�r:�m�*$GaeÀ}�A0����BY�l�O^ưN��`�
��c.l4��r��-$�F���t��,���ȇ��tѤm(����Mc��q2�����g�9�Bp{��� ��@�(�"����{�	f(�Y�W���}�`b���\,�K�Q1 |3�5��$�ۄ���	�u8 '�_����XR;͖��Y3��\���
��7sTSt,��ϕ�J��V-䔮c,���;O�=�����b��GKd�؛�o�z��">>������x���";��U���d�]rB-�aԣ6aX��p#4O0���1"�n8�&�q��
�����ggT�@\$:-����o�~�b�Ҕ+���#�i�&��S����VRUp;�$�g����O���pwfrzI+�P~e�~��	��GA���:EG�Ѧ8`�X
z�k����G�roPS-�9*K,�:����l���@�1�aQVv_P�YN ({�i���	�R�l�C6��rI9�h8��LQ���e�`�^���V���	��YXj�዆� F/��ot�����Q%��
�b�Jy)��+������҃Q!y b����U<��w"�1|#"��.��Jƴ���hqbY��J�`�_D>�0�Ld���9:z��A��a��9����i��	�Lݩs�:
��~e�Z3���M=6l}�%$�	B�!�6&�pF��u�a�h��/"A���2�WLF%1����S:�f�3<��,���<f�����G�J����:�R�A4p��<����Q�i�L4Ti"��S3�6Τ��P�p�ρVxy���Q���R�e#;A⎇����'���G�����|K>���`Ⱥ����x��Ah�9Z��$Qҳ�q�z>��]�K�-#���VZ.�c�4������w�su'ǧ�!��y�P��v5"�Վ�NP���3j�:�ޙgt��^
��[��kO�F	��&�I�\���)pQʞ]��s�QV�N1Nz��=j��զ�U�@�H��Ĺ,�A�y(���m�X&���?M^�r�h2^�^��D�����)�Þ&΍�����yh�꥛�Lhݺ�E.yP)	�ѽD�s���6�� 6�Ǉ����=M[k���K/�v�'ǈ�N���Mt|l����	����'tpD������BΕ����3 ����Cy�< �ڃk/�Wr��_W����i�`K�D%���-#D4�·�K�([�v2�~��;�z�J7���F�3u����EY��[;h�x�v�I8Pܬ�!S>�:�y]{��xN�)[6Φ����&ıQ���q,�<�:6r���5�.��&h�KENc`���LW�>T5��ǆ�?Y��5��9�'  YE{7��������ζ�"k?:��sMc�#�δ;�֗s��m0ֱ�ɴ1w 2��F��|̕ɨ��G��4w�U��N6_��8�Y}��s]�!t?��}�����A��j��% v�@��>��[��a����( ���=����}�OX����L���z�@�������7����}d��u�4A�媇��ǎR�ײS�CWI��4�o��n�����4��Z�����8�iĪSS/c�GS6ZʢYoi[�/�Y��$��&�\��#�6�oY��n�S��ۿ�N�x{$#փ�D���|���@�eC�|ϛ�pA���[��ӑ��A���-,L�N%�*,C�� �a%���Ѐ�K��*��i��S�ø��Iϛ3]��e�ȥ�
���hpt��dǒ
1� }������;�kٽ0炮E[!_�X +]���`	��Sm�Kp����Mm�i_�e�v� ��@[�5R8��29�}�p�W-�=��D�{���9B�q���K���z|����"�o����pM���e��!Z���%e�`m���*"�jbW����H.��j�1�ɱ�W:7��>vp���]fb("��P����ȥ�)�?��!��l�̤�e�D}?�瓮�g}��H�N���j:��}�Әz�4]<_����7P�QmdJ�]��"l��|������2�8bzt�!1|` =h�̣��#K���M��U�
�����*F����*:ȃ�M˧�3^�����#�M��;T%Bb��3_QP��7��I�v@ᓓ.��SNѡ��t��V��@�������32�&��J!�t1��	:��^�	� �*��#��^��b�`������tK~����Dj��<@��["ߺi�F#��J���r�F-�7��������M5	��E���Q��04	!C`酡���vF�O��h�u.E<���˝���s�6�N��M��⠪������c�Ҡ-'��IQ�;�3@��mAͯ���J�����1��"�2��������k�l��Z��a%���}�EX	ځ2�E��]ԓ�
�yv�6 ��7�.9ɿ��5^��ܺ��E�	!�}7X�_+w"��L���~e����D���6gq�Tj)�|$ķ:�y��߇w'�s]|J���me]�D�-�����Uې��Po���1�~��)}��b���|�ZP?�UndZD�So`7C����Z�&M�[�*uIeI��V<�.蒴3�z��(6��eG�?9ou��DT��@���M�(ꄹ� ���4ڐQ�$}]}R-[�5w��5�w���#3-�V�����	�V$����v�*�����o:�f"�:(��_Q�{���'�i���<%����Q����켳VO*�B�툎�6$���>Kgn�4[���#t���1�&�k�P�|W�Ф@����>�������q$=�jL4�3����� $"����g���r8�`$[����V����0̜',@����Ԭj�f,��\cQD		okuM��D'���R����6��[ e���֯�������ַ˞��N!1�����=��J`�d$����o�#e�VD-][��������5��s�+(���fo�í�(�#����qwC��t�Y$Ŭ�G��uX��#3.��5K���Q]_w&�r�U��ّZ:�f�c�����Jk�l���ヾ����I�G���><���<$��zp��r��Zc��� G �v��3�)#�������# L�GT+�X�f��R@�)��N�P�w�=���>��X'��H����Am��I3Km/t�_Ú�z.�|Xk�����%z͋	���27���q����	��*��q�n����D:��̻`::��]L��6�o�{)�����{O�U��lӹL��ZŔ�����ľf����!]}�@�� <8卑7��Ŭ�P�B>�87��r]-�,�-
]=k6�֓��<V���憟���ߢM��Azw�V�{N%o\(�Ӌ@��O����8@�?g:�ދw�Q*
1�0�I(�[��[>��n�D�t�W�¿�R��W�ȴ?Mb\����@��ȸ�E_�}�+4��_I�k��
�;8=�L>��z�<�E�d�2��n-����,e�3)�۾2E(Q�u�N�B���(�_��[�P��ER�#|���>+�����ꗷv�p�ڭ�r1'-� 7�G��;�~d�.��iB�}�h��+���M ���B3L��j�~���_�r%��~�
u�ɨ�b{/��L$���M�`�p�%#�L�#�n&�d؋�͹Y-;��*9�L�#�C2庝,~ċ�8��h&�)��=�n)E>@��Fa���,}��Bעv�;T��T�U���>�#���D����9`�q+1o���ʇ2ˎ�8�j�Gzw%�t4cMgu�]Q/I2�re��� ���Wcٔ��E�
��ٓM/�%����c�$���A1�cH_^J9�vs,y���T��.Q�I��y<j1�d|}��CT�}�>�Mhk�]���U'�>���o���[�!��~FB�ڧ� �$�r+80~�d�.�
y"L�QI��d�si���Dg����i��B��vD�κ���U�q_�i?y���p���/�
i����&aإ��١����i.�-#�u���^^��ˣ�zAE�w�ʝ�}'=�m�2�ԛ��XhL�NIʶU�Եl��6�t[���\k�Ö9�����N��dm�9��b�B����������Cj��y�5r���h��S�rN ��u
�*�1���G't�B����z�p��%����&K�ma�F��FE�eJ2�SBdIz@���t�ìv��dKCf�������>����:�R��������$ӯ2V��P�,!�SwE�]�u��d��s�zY4>d������,����ܯ����!v.@�"v
^��z�^"�6Y�=&�=k�%"����)y�	�������%X�g��/�Z0�I:�����Sfh�z JM'��I��>��?�߻(2�8�m*{L�q�z��<�DFf Qpb�ǅ��L?��7&�}�G�Z�X����~x��=]�8K�e �me���v�*�}�4kP�"gGW��.�������c4J�b��[[um��E�0������v0:����)�V�-'�Eͼ�_5U�c�-��_|���H��B�����f�H;d��l��kW8NlN��0�ޔMYT2�����/��ܷ�w)s�͞jlf� �l�b���6�Ҍ;i@�5o*.s:U�����K��cYm	���o��+�<Fn�b��Q�`W����/�/���'���ǶhXTV�Nϰ�Rlޜib����������)�6����ș&���3�k  �Gaq�N�d���3���qo�PG�p
#�|�a�(�/6��t�mʋb�Y1��VR�������Ɩ��7_>~���-�G��^����R��_��ZG.�"j��6�����Ú�<�ZZ�KRCdC�'��L'ΈpXx�E��[S�}N�!jJ"����Y��sPzf�j��h,5'�+�i07m��c�U@��j��ձ%�{�g�k��V\&��6��<��G��X��x����,�BYx�=����[��,�xadZ�7)�n�E�)n���Ӷx�N���ɮ��J:d.z����p��3?κ�8��q�k���C��ĳC�o�osN�V�q Qm�ՙ�tb���İb��n���e��A���BiH=�<����0�9���=�Q�2ް���z���"��������Ɣ(>mE��\)�O������i�Y	=��"0�(wZ��WO��S&d�<�pr+����
)=��\�w�%�Ԣ���=bjg����{��ؔfB0��}zŲ�R�E&��p�{ׁf,9��� ���e�g��ɕ�JJ�F�&��S�$�d�Jh����8S-}�i�A(!�����o7���>�i?¨Z�û�(�3�Y}^��I0�,�N���ۑ8�ϭ�:�
Y��vߧ�׏��hUUuj�/��xj�./Z�^��!_���p�)�������n1\A�/�
��F����,?���ј݂qk/_A��-W�G����%G�J���%�߮��i2�tqd���i>��/"�&3h�B.��j�GQ��9�u�`ݹ�K��ث�yY],�l�!�뚻���c��N-,�F6�r��@�z�bZ�.j�}F��.�?j���M�6��Ê>��c?��B��>�\��e嶬=���S�ڔ�绎PQ)=Jhǃ_�w&g����3�v/c��[TG�v�8+l�^
mtjZVzt$'��еV�����; kد�{*�a�8�� wx�v�uZ�k��#��y��c8��_P��vJ�����}p{�<!���fJ��ԉ����Q��Gi<��������=�#�/�e&������2�c?��֠_��ɏ��6Yݫ[xLq�(�z��ΌI��Ґ6�	�V�ͥޜ=�ؕn�^#��Ջm3����ͩ�),㍈� $����і�/lg�5��-�Qu��b�����"9��/��F�Զ^GS��v����?�=Y��� ���p�H�n�խgs�|��s3���eG{�������(OOA�8 v�ia���6{~~=ş�(�/I��D@�A��E�T��H�Y�0/7˜pZH<c�@o�z� @�5B����G��}�.��=�+�RE�ϣ��Խr�O/�!T{����~�8s>���Ŏ������ju.��'ڢx���~�1��X�5��`�fks�+=�>��I�;m��7X���C��a�lv�sBc��ބ3v~�Ο��O�E;���"azK���~>v����s���>Ľlt.��p{@�e�k9˅!B� �<382~'�y���ɂ�tϔ֤��:|�R��i_so!V��ܦ���Cf����8`���i��s�ԍE7po �G�b�"�f,��%��(g/j�ñ�16.EfZ�Ş�Jcܤ�9/�z���۹�]���=�Dh �،�*�\:�<���^S�����t�Q͎�)�אEs��2�y8Ҕ�Q~�(C���eIx(r�л
�ș�)�Z&^��(������.�AP��Q���G ���l����C	�N^p�F&�jӒ*(V�H[���eW�U��5�&y�U��P�q��"uf@���Q-'��/t�1�F�r:��N�|����\=�N����~z�!�j��TRQ��b;��m����3��!w���X@�2
�0-U��b�DX1R^�{>$�>�>�}�t��N�K�e��7.��e�F�>4��Lv�t%�Ӳ�i�oPX�,Ǜ�H{o��\y��B�C�M��0Uk���[P��Y�T8�k��[����f�θZ�>t������-��y�b�w~y���a��w�N<����c���Qu���?��qŮ����b5�o�	����J��+�����'�qp������pzM�R���ԭ��G���3��W��~����q״E 0�w_�I�w�$0廨Zd$�o�ju�6���.���F��-#���ڝw��g{�k(M��պ�j!/���������DfT�*��F=�?�з�.Wh4tU�XZn"�pW�̸ۗFW�+T�]8x��dd/],IXE��͵+�M��D4��@6��p����+0�V.F�=�������p���@����4�g�t���`e�GY��S���ˢ�O� �<iAJ[���@�vj�&�Cj�iDvt�P6��c�='<χ�1z��Y�|j?Z����0��w���,�jV��}le�֨��Nsl�X��j����6ڀ�Ε����_y��q.�Hڷ&�Ԛ�.�[�w��@Z$�c(phd�\D��6:Tݚ��`�/њ�����¾=��#�}} 9n7�֡G�1j�o�Si&f�qy*?�h��b��o0���p�r3d2w�=����n���f�9��QHR��{eZ�ӵ�x�����|�7�׺cYCf�7�ƭ���$�s�X$�|�'?q;�=u��}?|cKZ�[�}<"�C�*��pu��oZ��?d�j^Ŝ7!�|�������shp�0�Ng�P��ȳ�k:���)T�,��M�F)�=j:�3�(ᑦ�P��H\�X�e���!Y<�
�����|�/��r.etrn�e�ӝ�X����ޛBA��:�&��yْ��lھ��XT`���-�����#UkL��nJX��,"��>�\N�9?� ���Ԩ!3
?�me��}S޸���e�f*����6o��|�i�YOM;�e��kqKY�TI�z������#?��+�鵃X&(��\��6�G�d#'So|��'�x�wY�S��tN���4׿\�����0�W�� �b)@�W�:��f��}��¡�̂L׿F���!�V��P�)H�4g+*|]�Xj+� g}��޳^����ǒ?B��3�ΰ�\ǔ��%װ�c��DQ��3�=�����)Kw\ցA��-֚˿<�0t$�փ�CAI_Y��\:����潥"�8�I�: ��`�lu��6�2��D{��eՄ���<+�c~��>�öA����7Q�8�hⰈu-���/VIy��9���C,0v�U'ĥ~B�i�02�捫�q!�RI��>��>7��>�=��ʝ�N�z�T�g��~~�cb�!pa�'hZ.�b�uAl��M�b���
�r:ޜ���=QP�o��U�8������,�U��k���Ʉ��l�`L&5��|�����$�4+�I�u�7�@.���Xl����3����-ʤ=m������"�ƅ�ج5���5.@�@���ՔU`?e޿S�b�vp�������
�8�V�A�?֐�R�?�n�e���1�$.�,�w������w�P=�fx��Ӑv�U�`�P���IQ���ߢӤ�B�بG�T���δx�D�P�Y��B�8�S�u�\�yN���U�j9K�xȥVH��c'����R&�Y˂e�o�\��	^��S���az��E���.�EJ��ǫ�A�6E�W�ب���vA��T�
k��(ʀ�W%�Y����A	��Ymq9|��k�}�O�����V���Z������*�&Y�Fa��خ��r(!�v��oh��>��(mP���L��x��=�󣰵9��C�k ^�v52`����_d�d_�o��
s�8 \C�i�-�j�o�uOZu��@D�˓B�L���;*�ot�pa���A��@xB�7
�]J������0e����e2�o�Qj�Ik�����)ؗ\Z|�%�F}ſ�� !��r�k(7s��0�@�5��W,g��=�i�9�����#?�t�o?�'|�{9R;�����������/���v}�b�h�1#w�2��r�ܦ���є_K�o�M��ln#�t��u�Wk�:���/O��-��'mG��M\F�m�����M�^H�t�Az�ډ�R�D9�i��-jM--wo�G
C�{�J��A�K��:�X�S�Ic��fQ�ŝ�#�E���Jb���B�W	cI���Ws~�9��'ԓ7�V����T�Jʀ?�?���j"�o��G�s�̀G�'ٷ_�Gp)�['��OR%l�-���k���S���`���n�Ů]{����4ò���l���==�a|���U ���F�Dd�N��@�vz
��V����E���E#T��L��[1�S���]w"^r�q�9�ܵ�^p�wT5��B*5f/x�´� �>��w`�'xJT�X�M�ˊ��n'�}q���X���d��ɤk4�$�X"�H���|��s��a�:؎��:Ny ��*����V`�-��o����>.�Q|���td����_�^u��M2�X�b@]�ꨅ�m��q�4�g{�F��b����fTz���2�zt�M���Lnw��_��rWM&�s"�^���CǾ���C�WȆ$�\8��g�
o�������={{����)�+����n}�!�i�}�6\mR��p�6����]��~�_��p:��?�'WU�z�d ���d���B���d��[���h�GL+�ݲ,{LgY@���!�~g���]���!����%��Q�U��>�A��o�˃��W/��5{AN~0��.��e_��s��ϱ��P����x_EF$c�|�Kc�~���*|Ev�g������CV]��cR^6���X�nE�~��CE��}:>sW�
���`]#{��U����$�A@�%v�0U�dѠ�U9lb���r)01כ��E�� �K�vg@/�+��4�ySQ�����1r�&P^g�h�H�kX[��5io9Ҷ:f��qk�4��ﵦݻp�,�ؙ]���!�e��&J��v�o�����mLB�|}�T�<�'��
�`0j���r:����X[�Cx������$��4;�+tL������["��^�|�~��?v����>1F����2e��س2-/��ԍ-f2�J�vB��6�l���ʲw�(�{��������5l��|��hX��)$BS�w�<`pVt���$�3i��l)lG4-C�˂B-I 3�UD�&�㝨p� T� y�2����(��y�ֵ0�@�I��G��߈�	eH(u����dj� *��^�Ώ2����6K0��b��2I�V:p���U�	Q3G���~��,<�-P~������TZ%�kqCiu^�D��|9�0�#u6o¬��c�s��EY���D�.�0�x�~�rV��}o<��>S�1�b�S �� m���BrPHLv3���UOM\�����)ǵ��� �V?:��ƙ��Y7�Ev�g�_���I��W��qo~��<�����i]��������)D9 ����q�<�0݉���oR��w�T
5^�VK��& a�9h�7��mNJETAC��h��h��I���v���4E���u���+i�RD��|:q�K>|�l�V[�y��i9�um�v�[����Bt;�[x�fS��rS�tޭyl��
��.v1lXN~a�i�N%��9qե+���2�;EByva|� Sܪ��J��6i��i�Թ�w��� V*�z_~�Rn�KVR��"�?H�컃�D[8�m"Iq�p�����#A���?B����ֻaO����$�|��>�R��A/�雔(�`��:��޼����O�?~��>�b���KP݂-���{�l1
;���\y}K�eE������`_-�>�߭�Kj~���@L҂���A���%���%��3��?WcM�Z����sV�̈���f^����L��q��K����0�h�v���KUaho�/e����o|K��f*q��S�S{A��b�ȸ�=	X��`C�0|��2�H�(~h��T������j{Ѥ�hE"1�L������Y����w�Y�J�]I�Q�q�k.�}Aư_���bڳm�[v���Y)K�q�'�n�^�\��P�l'RT=Y��p��q'����%���C�4��q{6����sy�NgZ綀˂�l��Dx�x��"X�.�a�J;�q�H�M�WsZCNfD�N�?$Ǯ﫥Z�y+WG���>��h�|��	b'k/x=<�Z������8<�i��|��U/�5�^�t�����:8e+�N.ϙIn�/A�{��$ڣ��7�ϧ|̷+���/NX��&������TR:���c��/B�ֱ���C� ��|�'�c�s즄`��vk���C(��c�{*�f9:�����z�����7�u^�բ����\��)�uߢ0=�_\[�ö�Ъ=v��rT�]l��ۭ֨��k�G
����݇�?�q��$���0RwvF�H�odZ2�:h�A�PL���`�ʵFi8�t�����O�D�'�"��o�r�ˀ0�`� �Q��2��<m$���0 �1��(!!d�i;�`�KA���͢���>2p'��KշV�-&���~$W�t��V,a�V[7:�ƈ��pڌ�mǰ�Ѻ��fIY�D��{��Ǹ%��-5���DӚ{� p���E��0@|_/�W�̤�������1������?h��
XLB�鮊�g~s����?�<��+Ń�&����Ε�u�=��	T�[�瞏���~to,��F��_j�0|�0[R�!���\���	�x�����]�k�H]�d�j�M�>�<�DEC����W�����_����'�ij��ca�?Tz!=�Wy���%��p=,�[�g������=���7��MfZ�o��/Υa��HY̱P�n?�Eck?�����A<dF�jrMm��$B�&¶/���[�8Ze��m%+� ޸���f��<+����P���3�p�c��b��P�2�;��"Գ�>�3�s֌��J�C��o>� �� �C�H|���ARɊ�U���N#!}����[��Dc��0t����Oi�9�fYy���(���,j3�7���f������bD���h
�%����yx+�؝$��s�Y�j�d��� �~�	���C��h���L�7�ڊ�<(8c��𤟟s}��'�S@ #��P]�_�?ljX�Pb���>�O#�id��.���*�X"�n�rK��bh��Y��Z�J���V��6��G)��&���IC��[�
�^�.��O�~��
�9��p�@7�c���/w�1����reC?&��n j��t
�����X��zqԔ;J��vu���̘X�^�-��|Y��Iea�i��\�]Vm�����q���iv�G�Q����6��d3�YXU��1>_�f/�*�Q��*9��׍�$,u�Fqn{s�X����R��8v�}<��Z�<����G<B�S	LS��� 	����Ivr�]B�����XJ�/z\���5�.�n��6�M�-E�) ���,8@�*ڼ3O*�6�a�sq������[N���v�.��-���r�%K{:,���D�.e� n� �?!%�)�(�wN�v��՛�P�8,'���������Ȳ�#
d�I]X������WaE�>Eǎ��Y�d��4��^ω��Z@h@����1g	Rp��^��9���vk��a4�=B�V6��6Su]j����!t:Pòd)g���@cgh�]�v����/�w��#1�L`~��(����� 1N�!3���GŨ솔�7#�h�����YN�?�y�ih�6|`����c?\���a{�����iqr�T��I�3�#|��>�i �F���|5pg���E֍��g\�o��'�u�!K:Ǥ�t/ �S�_�J1�E����p�ZW��cm�Þ�W2�07 =�m~-��⭔Sܓ[VF�Ŝ�IDG C�_iNE4W���N�Wb%���!��b4sڇ��.o��3�����x5y_}f���"��A��Y��<YD��k�S{  �y�� �eWxo�����[�M �x���!�Ta����K�6EG���a�L�1A�VJ8�7�E&�����	e�6Xq?%����W�V��F�U��#a�7�q@�?Q�̕Wg	U�����Ϗ���M����P��'=�dO<j��O��U+sQvO"O�6�������8�Sx9V�ӈ��{_��Ugo���U�h�-��7b7�)����Ȱ�e�WۅFG����A��uf�%]$|u�o�^�����	��N��.RxF*Aov'z���k���(�f~S!�9E�0���T�g�$q�S������n�j?]�`g����<�PIa��Z�����! B�����[�)��2)���(���� 9�V�ց`�icX��E�+c��*Y���F�BϬ시Q�?C5�&T��H��W�3n���{ˇ�p����[���S�!��^��:f���J�_��Բ�N:��1�D����kw�7�-$�L~4������~����!���7�'9y=t �h򃥾��'����)^%DI�Z��.�Dܓ���� �D�y��Rw��)2@�x[2��d��h�ʩ�漊����C_>Ku J��"��\����1v�y7�����4Ϳ�A�b������9H���՚5�*��DkN"�-���y�ˏ�1M$s�8�������(<*��D�B��
q��gI�'�4u�U+��j��.#���¾�Á
�q�ڐ��n�X�G�m#���m�o�c	Dw����b�ȇkP��=�JER�1�YDc|\�w5{��tO�3��p�'��� �-��ׂ�ذ�Nb�;UT<��q+y���3��܁���>�E�5_���)�5�h?0��)�]�i�lY��1�1��yn�>^�Z��0��ƍf0�؆
�8�[%�7�(�ڔ���.���^���,���3�V
��(�Bd��}�k��:�,,����7��u�F�G��bf
J	Z��2�MF�������a��$��gJ��E�s7���١uM����.�8�L��sĤq��Z8�r��Rb��쀂z� {?M|�<���HD��j*�8���|��b?���q}������<|�E6����J�F�h�`��Ի���3��E^���A}u4���ª�wAg����8 �͞�;��|���y�U��c��p�0$!�ˡ����nA��g�l �u��r7ϼg?X
Z������kV�W�9��?��߯$@0'��s����?:��0�C
����ɉ3�\����o�
��=he�x�U6&~4�!I1�M����5ai;�\l%�+�#�5Ů�ݲ��a�g)v\S�N��%wne{yp�^��7�ge9�?5���?�[.�Y��,�m���v��^+b�ҎHT֌i_`u-��{�ZBie%b�F�+v9�5�R�=2�:����S��n�y��yH��ܬ�U2�Һ��˜F'ȉc������yA��Ҕ�ou��D\������R�/팹h���=��� ;_��;������Ĥ�p6"~�	�漺�\�g�3�3�dF�k��S�((fN�<F8�6�A�3�ikVG0։jV�k���w=Z7
ʔ�6x<�������d�t�bK�g�9�V�mP�&�|,'�Ɣ��Q �p,XQ��G�(N_��T�Zv�f9��֦�❲ �Ɠ�7F�X����##|0'b�Z�������~�+��:+�q4��w��&�/�&\נ�7tw�v(�qħc���!��m$�i��)�̍��A�����y�UHT+�k������<�5����C#�`�V'�;ؼ'yг�ի�I�S���,5��J+���#�4fgn`>J�WxUc$k9�MS���A�W{\��*u`�_��jݣp��&���B~�u��Lc?�fҩ�χ�kkT�I-rI6�H�o�ƶ����O���J��0xWN�*ջ�fY0u��# EY���n�W�x}�$z��+�(I\öE�w������4
�}ԈJ�%e�Ze�G+��#,	��\�j$���]b�ϧ����qSo
TV��1��җ4�׿L���Q�Jm�m4D���ن#+�<�9�	������U�t�z��_ˈԪ	k���!E#U�
>�S�K���$�D|{o��Qpo��ū8�'U풔b�z餆c�{�!�&?h��v�.��f���&$�^�o��D��8�g��8��>��(�u�YB��y�[�M=hQ��CzFl����4�v�Vݲu�8�SQ2E��8đ�S0��:��޼X.�-����#s>L�Эr����ӛ�K��Ŀ����! ��孑���4�o���Bw�'�q/�����0B;�%8��eA����a�:�nG+�2��(M:� �z�����.�7+y.!4�_��vW����Sf\1�����%�4-/�x��Km�����u��)H�Y�7��o���e���Ζ�l��<D�40r���Z�ӑj���%���;/�-�IVĻ{���ޖ��J6��iG�q(�(]�P�F��<��� �	N���59��H�,]-O�D=�\(}�H����Yо1���\�B�]Jrx�����F�k�Q�(���ס��x��af�z��"c�S����vt'�����lu�q��,M�~a�l�v%���o���NL5�~��ػ;�!�h���|���Mn��s��%0��H=���(Ul��u�?*�}��|0�Ib6��n*C�����a�"('9E���r�mo"x��u�!�8�'��e�>xsr��amW��bڅ�o6�s������5q����]�DF���gj�w���>�x�d8�<���=k��ܸ�ǜz�[�Z0��� �c?�����z��_�z�l3���p��B�=��8
5Ukc8Hª�6|.8�w�-+�Dߗ�X\��v$��N��U�����H�&���M���$�b77�z?��S�	�s�BתC�i�=
78#3�yZ&@GR�1�B�"�I�k�\t�%��/�Z��"צ�S���ݿN�S=�"e�X�O�	 �=�FsZƈ:���盨jw��Sl���Ӵ�~���&�6�0������*�YSwlKĝ��w_¶�di��2�z�یFۥT���U>}�(�3!}O�����1��c_M�7���i�`QڙSa���MEO/g��(�А���f�Ǭ��'�1�W�0�Z�A.	M�Sp��}�B�^����b�7�b�'
�(/����"pR�U�N˾^�{�F�0u��k�����>�(o�04��� o��E���|�H#�``|��x7z�@�̅3"�̗��M�N�7C5��M���1�
RUgü�o]��>��#S��4��.� [;py(�AZ��&�Xz\�عi4<T]�o�|Y�f��^`$�ݞ7�F�4H7���..m��/��Z���i�q����Fu8�W��r2qܞ�mOY�{5f�Efd"��C�Y��F���1��8~��T��evp�^����_��ڕ�Q��	W����&�Gǥ��͏b���T�¹p� �t��f`��ZP]�74>�+�_���mr��>M��K��>\��~�w�P+��u�x�W��My*�Nl�fBh\ 8��;ϛ��ʷ�P��Ħ7-"�5��\SxO2z2*�x+�O�<ɽ�;l�!B�7��]u_2�e' ���hB���qۄ�� ���R���V���*!2xv譌�͕}��,2��:c0�8HDK7Vjk:Rح �싞�ؐ��ݐ[��78I&�F�KmӱW[���1(���bt����!ʺy�|����7�:� �9R)5��X_�i9!��j�������GY�65N�g%rj.Q��	���!v`n�^`̘�4a�N��o�q�|Hà��~��8� !�%r`�SF�*��h��oXN���̆��s}	�_/��7�x��0��͆e�H{�kJY�f- �l���[���#�L��;G��&'ݙ�Y��k�6���+L�-7p�t�JDA�^��$�<f�����P����嗗#��5t�{vCj2l�: ���k4/P���>�|"��#�v��Wq�7Or�n����C���z��F������<C
/�Oy��ٹ�����G�����j+���3wcP���<F��
�)�Ã���.-�L�CD�Y26�P��5�1�`_2~G�@+���>���ez�PJ�kR����-�!���Jk_e�*=���n��z����}T�v��E)C|Y�� �1��(�%P�9�xte�	�`�#g%"
fCw0�@�9����ȶp�܁bQo�U�k���r죠�k�PZ�K)s�N�{�F%��D��֍���ǬK�7O	Q��y`j�=�>�O���2���Q�K�]Y����k�đMe�������U�F>�2���,t��$��DR�z�Cx�"�r���g��Ȱ�9�'
��6kC���բ����b. ?%Z�-ϡ�x��+�j�p���^��R��uZ`��&�r �XQ�dp�����q�, t��U�fث��K���-���w6F}�W�*�Q�S;ړ�t<"�4{������]��ӗұ"W�7ܓ^�ߣrJ<�z�n��mV�_��*��w�7E���Ue��$R��-��@i/���䩛������F�^���g���j˗j�p��A�{���I>��AK�&���s�2�s�ΖK�Q 48"�>/;���2�2uا��XQM�5Ӣ'��#(M0��?hM�H�<���'��<,mpY�7����la䴣b-�0
2���۰y���H�2UH�'V�mgh{��dO��+�ȇ<;�dz�%�PDbF�'^��^�,�$�1]����}�Ơ1.��Hz�pB��K$���J�;y�ě&Lо�=�U.��=E� �gC�Xe�Sԝ��P��|�"H��U�IΟ��x�N�%�	u�N"�E��d(��5B�V�`;͝���W�Z �=�-���q�kf[Z	r�U�/Mj�����\%cfW�e!Ry��_�v���g�#I1~�'����Ү�W��ǈ��S��:�S򦏗�3�I���qޠ�7|r��o������X�*qX/����%��Nx��(��=H���t-iiEie����FWX2����	�-��(<�y;aX5檆J�t�@�h���\��k�s_�<T�"H�8�(g��Oh��(�� �Y��Jec�Q:��}��L��u��TY_�sCÇ���T����Wy��	W��˙ě�o�������D��k���n�y$-�S
D�})�&5K;��87�|�D�����/"�WFm�z_b~�g���:�s6����=��}�i�'��őbd^����'�(.�w5�t���/����7������/N��C�q��yBt�d�Ρ�1c谻 Fvo��B�"a���/���QP`H�E��X��`~�����,h�֐�M#�5�(���"tn�W�=8O!Zh���#�s��?*ho�7�>�ŗ��oܭ��9<L�1`=&�к@�?8?�yVp?hE�2x��;��w�,p�l�u�dgj��=0��hW�&`G��V�d�A>�%`�_i��@%���'�JgDc^w��ʷ�8��;�!b�g׹74)w�C
�UZ��틀S<t�i[@����5�~ L`�*F�W6�K��:fv2�>/���o%|�WE��K�����f\I�����!5w
ޖ1`�6��b��s,)"` �_���~�U�]��%,�S�FP��9}Ʋ��Ϳ��8|��@����1�e�Âҙ$,A�E���JZ�"J�B� �>�+n<Ѻ���/�G�����pujY�y��@ 2��
��(�HcI��N��s1����)���bf�+hy�D��$�]a�<�% ����8υ9=y�.Tu��r����A�!F�U�N�Y}j�f�/1ZcD*'+ƽooiт`��rjD˘�I�Z�s�X�S�1Kf�<%���q���8.d�$Nc�$���8Ix@i�
�b�b8��	����)H2�ܡA�#լ�ȓu݄|E/�P�
� v|���ÔG��,��^ �'�`9��'�c�|�XZ�3�؃���H���@��sc~_�Ue`I�YS����0<��:}��P�Z��E��z���F�ﻚ���*�ԭ��4���~�S�q�S��?��.�W|A�+k�#"��mN|����>Wi�0N_������Az�@���D��&���t��&]*�
��K��yBR�R �Ѫd'�Ru����+:u7�@B�uq��%:�2�!
�E�`��i[��@����Ko
�R
ܬUHa���X ���� ^t�(Q�6�QZT�4r�v��"�X{�����0�0��[�8l�B�K�-B�f{����-��h(*��ԸV@��N��T{Hg�OΧ�p�g���X�q��iSXۮQJ�:��!�T�z��S�*٘?_X�la$�U�
a�����.W1��k�\�$#�&��R���J_����R'�);�Qd��R��d�]�o(P�����g7�9`l�fb�{�!'�k�s�<�(	x�����\�Q6f%�o�B��i�ܿ=�4���w� `�X��M��&� +*����	��MQ42.�E�،�7����yf!�(}ёs螺�`K��4���U+D/�d�ȼ����p�XJ���.�97&8 ��9a�ykE~[W��CG�C	C��hj�o+I8�5?���/���"�ST��]wM���ʖ�(�7ѣ�"��3iP��3���_y[�(�8���s|�1[�$'l_����p6��>�����-���4iA���"�����rC���Z0�tba�=wD�ᙸ�7%ӱ~8�05���X��>]]Ify�e<��� �Ѻ��BfU��"�R���N��m^}�z��"�?�T{	�?���@}3P)2x�B]C�f�'��iI���3R� ;F��}8��yz�F����O/V}�����{.�:�#�=ݽas�0�_��[�D$���tsZ�pw��_�eW.���г�j%�4J�q�&e�f�i�(�$������U�ksr��dg�P�ډ�@�$C�Zȥ_�4⺛��I���R�X�k6f�����o�!��'�D5|hF�ht#<Q���Z~xڡ�a�`�G>���Iݝ�2�K�b[��UoW^�����N��T炇��d��N�k��c�|��Q(6ww�e�^��$I�r"a]�Ld�nIQt���@~hR?�<k�2$yʓ�H$ǘ�{E& $�����础���R�3dӡ.w�pƒй�V�94H��<�Ƃ�H�D���Il��:���E�H�o���>BT�&3	��ύ�b}�h՞J�#�>k��ʹ�E�vmg�ü6[=é,Q���K"`k-���K�i!��
�/3C�73�r�����Q�ȅ�.���C���$ώ6&�۲n�l5���%���[n`.�]���T�����}Ќ@�(~q���#Q��x*���ä���
s_��ʒt0���}��\��b}g@��i�������V\��,H��a%c㎹pH�c[���2g7�?a�)�a*�˸��[:�����$��y��.I�L
x��qj�`��Py9\F��حbz�
{���;������P&�M�osX:�?`^�k5#��j1��^G���,Y��%^搬������-��;�=�^�@�]�ά߉'=�%��<jIN$H�u*�LѬl\��ܥܙ�$�<�1���3�(�n=	W��.��u\mr���p�K�S	$���r߲�#����g0�OP߇b��M�����T������.(@�������{D3�����}c��%i�h��ta�)��C�3�O�r�V�����~4Y4��p	�ŷqi�Q��w���@'�U��7��Q:i��T��_TCWQ,�2�]�c� �̣1�`���Ё#��}���E�M%��O4=A��(���1�aJ֖�1_oG�u�1}���]kFjw$����5��6S�.�O
��+�l7�����+�kq�5t���;�=,�V�D>`�Ǐk�����V(�*����a��J�`{Q�G<��D���p����! ��Z�s���8�#r��(��J����EU�h�nUYC�:[N��DV�#U�>ѿ��ȼY�|�=�0��
��(��q�=��n2�hHmN`u崧|�oG)E���p�GN�JK�`�$7�)���f]+������A!ů�b�}"�w�Sg<�{�2LԃS�Q�!3����T�����L����\34���d��{��Z�\t�9�%fL�2�&8���<��x�k7Rt��	5�A��(��;�j>���
��y��c�����_+l��j�$�޿�h5��dXts�2�	Un���A�T�a�f֪�mXX��*���K���R3�]�E�N��$d��8�;p���kh�\3|Z2`�o +���_��m�z��?,m}�(��E��'����{:$��y1U[�#��7�E"��Ȇ�:�s��?��B�a�e"���p����gy�/��'z񳖂J>LE�a>��ѱ�K'�������VO�m?9��|(�i��!�d�	�:��g�H�t�H؆����b�3N�y쬳�_?4�X��]"� �o�k��${W
3X�c:�{	k(�3/t�Ĳ�K�)-���n�/ﬀDEʫ��E��c���'G�@� �U;`��5ݎ��F~��KN#u��
>�Ͱ��^���6���Ր�G��&���o�Ӌc�\�H�$o�,,x�$j?�[)�����8�o��Β@���
������y!�6�2"�c��C�49f���:ޡ���o�!����>�e��d`)p�7��[`�E��XB�!!Շ�$w��%r�S��͡�<�t����s\���lW��v��Pn	'��4"�y�,`iÑP�(T�@.���
�½�O��q>Ԇ&A+�tZ��ѳd\�����zd�|�)D���V��i��gx/���~i���6R�H5//&򓈀����ZjA�W�dDd�0�UgW��2���J��D�l�솷�F}�\�������W>cV s�IX��z�M�	FD0��mgN�ռ�����l˖*:���r��_ٻ��,�@4g�#�ғ��]�j{�˥w���Й�%E�L ٢�l��2LlT��m9�Y_��h��������-�T�WA�㐃����4-G��l���S��72K8�C/�[�����F�ꩯ�~J����_1W��~�7�:�]�*[���
N͟:UܸA��QQ5��lt`A.T�����gxK��꫖ �;��NU�_�H���t�%�P�y!
�o�տ�o�����d$�ʭw�ױ�e�J9�<wh�5����@�K�zH�����;�P&2鳭������!b!���M�ű#P���]2����Z#B����ND�
��YA� 1wA9������b�G� ���������瞋`�r�+n�;S�#�:@�@��vB�8�I/Bs/VWߥ������ʨ8�J�����9�z�H7>�eF�Yv�Rg.aj�t� �4���Q��j�yx3����Oc��5g��;�κ�Z�D2bd�;:X(�2Oi0g��]�u�~<Y�Y�dc���^���z���B�]���d�1��]a�W(~���mՙ
��t\��W�{�嶳��.vX[�fa>)��y��>��Nq>��W�b��'�XC��X8�ͭ*�{0�m�<�F���_�w�0Ze�y�T¨��(E�o�_�C'���M��z�
�����6��s�H�4:���L!=������h펯�`��P��Ja���׶��)LP�{m���H>u3$��)���#��~l��^Qx�u�p�J� ����H��eHvM��w����^ o<?��E��`�O3��,;�&+����2ʛ�X�����
��A[0�	Ak��B���Sh�`�N'S�@(���r�L�仙��vL-����TO��r�;���d$`u��r.զ�E/Ŭ̓3�m���8E4@���=�}p����a�΅�k�B�EGB�ǠR�aF=`b���lG0u� �x�k�zT��Hx�.�ZZ��<�t U�v[/(���&B��V��TP�94���/��A����#٣�tt�b뤃+����\��{e�M�p�B�����f�����˔h�aW����Ǩ���*ZL+��3���ʀ�e���1Q�j]*Ϫ.(��bȴJ{W9�T�{*�|��(("�<Mv�5K�&0�t�pfVo���;��bu�����~�=/��^_���}���	��/8'�5�3��1�js�B�)��*2���`��G!��-վ�Ctjfx��:�/��ŀW�}�d���f��u�:MA�b�^���q��Z�?D�v$&ﳛ*�2H�{���S��N��;��x�۹���c��"�p@pǈ������Ej�'���{�枱+���qM�I�� 9gu�Wr�l���`K��޸Uc�F0"n0f6�R����j�K0,�k ���ǣB��/���V|GY8��	p0���([���d����ϔ��R �l�l��z���dL�S��ں���(\��� >���-�w�U�ڪ.Й���_�Z�����M����'�Z�����n[3��y��15RDo�W�����z9�@Ϧy8$[�R�/���*�� =��v,}~��z�Ba���z0yՃ]
�j�2QjQ�*��N�J�렏i>ݱڋ���z��V��8�ey�6�?=�x���]X���{N4Mv�6G��1
���]YAo�';.
߽B6�lǶF�+y��U��M~�a޿F}�p�K��ҭV֤�T�Ϡ�p�r�X�OH��Ɂo��}���Q�`4��z�ms����DJ!�m��8<�O��j� d�NR1���^&Y�q�1v���87-�3k��I�|�K$W���}�fa�L����a|;��n�M@R�jk7]�����8���$g��S�b��_`!eX�s�`��%���Vb9q��(ekԚ���WfJ��M�I,v����:c�����
��}�k��7D��-ۑ��^�p0�LM�r7�1V�Nx%���'����za�v��u~"p�����+��dU�Ĥ���ע �`���H�^_��W����_�O+�#_$�/��%5��3�jE�4wB�us�bΒf����ɛ�l� ���X��n8�A�%z���|���蝷���3�"�$�_���',����`Z^!��pJ��Q-=̆Fz� �$�2#�Xਥ���P�ݞ;��&g τk�2��{�qVr���uF�D�_?p4òg�wH�]qf� ]���ҵ��P�!g��cU˜�FN�𩫘��}�6�6Ộ�)J��Ԙ�����7H��/�X��Ƨ��UI�;n�l׊���9��B�;l�>K���3�"�0�'SZ���I�8:ޫ���х�.�_�ag�Aѵl�ܫΕ�.����}⎇?k�$輴7A�ǡ��ZU������'�7����>ޅǅ�[kĮ8o�&#���� ��tR�h�9S��3R�W�$x�.�M��8`���4n��&�3F�%�n���n�è3�����m˞�/��H��g@vS+��G���!:�Ћ��B �����奞>�{&���'$?������b�O������6�5mp7��!�z3�u���1ն�r�m`{�dyȎ�+��3ʲi���'�^E���gSt*�Bj���V	����1��ἄdG�;"I�$����\��D��3�֫���}�?��R��YV�1�����L/d�J ��ϯ
�3rR�3�M��,o��	l���:=��̟Nr*O\��
W�u�s�Y�ħ���W7Yx�hH=�3d�&5���1�J��V����/��w�s�b���+S��9�ʌjGǧ: :��ǩ���V�¨M8���Rښ%�5}R����U��^A��G�ue��Tcɚ��y�C �q�4�I�]�E`�����K��+��X��o?�`����`��GrF�6C���;7rZ����_9���|�h�$9����"�/Kf��ś��V=v���W�I��?/�z}��@5f�G#��;�܄�=�)S���1.�Kݶ~��a���м�r�2Vܵwd9�F4��Y!��k��!�-�h�m�h@d�ZooT/�A���sb����x婆
�n_<����Rw$�UV�f��T�$T�0h��b�iRS:pֳI��$m��P���BO�NU�yT�^ڠ��`���^؝O{�/Ͻ��.�'��$¨yk��)�s��R,�����I��pO�?�)82{<��-ԇ��6ti���6��\uKc���@PE��g��R�P ����yVQ��;�9�d�������S�ptC��STմn�~H)[r���[�G�]�	Ʈ�J��m��X����-��� e#�Z3��T}XL�*/�ƪj��c<�F&\w�����9��-�悥E����蒈� �z݁�@��AS��ь�D�_�]}��{� �L�����K��}ud��d�v���H��Ci����y�>��Hy�_(���f�9��QS��Bi�/qZt*I�z��y xU�ڑ�3��o&8��qX�<s��U�QTI�ҁk���[0l@Ӓ�T��ķ�;�5��H�3'^��P8^�J�����fz�r�_#+ֻS�o�%����|�J��nr��v(,=�Pv4R�ty~=k���1�V�ۑ.��?��Y���᥎��/2�}�y���*E�xy�P5c���_џ����l'C��eRL�����kEގ��VXC噝�\pD����fSw��h<[�^zvz�z-�/̒�~ӰW���t�oԩs��"���"��� �}����U`u�D�]�j��o�ڰNp�0)�a��5���:�G?X�u��`1J�4�-Z��x�8�h���L��\3�H��g����\3i�)]��������;�?F̈́i�W`��0�u�H���(�g"���!M�X���߷j��7��{װ�`��H��"L�{�Fg���
��=��Aѩ�m�a��\�va�ۃ!3�jB�`^1|1+!�;U�+|B�+'ڤ��Z������<-�-�[�#��*�nw��0Z-�4����_ۑ��S�O��R��wd�@�ض�V����=��.�$#w\�%s���sBLe�1~q�Z�cR�H,�W�O>�T��ȃk���~�V�m�8��$hW%��P��m���Bu$-x�QAD:��v�+0�l��P06h�F����0)�z��V[<g��9�D|}����0${O"��hK^=��Zz�(u��˒�]�
��"=�d^���������º���a�t�4�»a��:.^��p�G)~S�÷⮟|-:~�?���6^$m"���o�F�^�iG��A��~y`�S����o֞.8��a�������)ğW0���-�s������� �n�o�xt�u*�_�?���G���ys�+-(;@�����QD!�����o���@�ܜxu-3�~%�A�}�
��=�f��t�'� a��E1g�w7#�,�P��~��F���]�4�|�/�F1��� �fK8��HQS @�����P���c��%��o�����:��\�@�	Y"�|�\���|v�:V�p����������J�W�RyB�iT��F /��z.Dq��ݿ��C�nƩY$΍�.�j�?�(�"�r�l ������]��oM���	g�3m����������Q
��[_h���sS��USNʍ���s�M�b�\��v����h�۴�~[��6���F%���8����A
�gحS��|���އ3;xҙ�<(��n
�����xd��D�T1�Q\Gp0�
Ѧ�2�|�yR���5ٶjc}�Iw��te3�I�?�4�vQ��J�BN�X��+05�to)no��������k�#����|�D���l�n�f.n�zЕ�7�˰g�[j�#�C�S�A� �|[��^,�������޺5T+i���c��>�o�#���7����䬨E樳?:�0��8���o[(`�p�4 �Z�U��(J*	k}l��.XNRA��o�z9�clW��O�Pi�U1?�t��k��}�!ۧ3���}j �ԯ��,���� ��� ��:R�l��u���M൰�n�i2��-�d�� Kڴ�/���u��/7=�������͠�,���) ���C����w�J4Dh�4��#��-�x�8�;�jJ�41�R��ky��y�Re�brL��N�%\�킫�� �5��S��pnm�м�l��t苐޺x,S!���뽜�����sI�O.D��%_��ȏd���]���S)$��b�SUrħ�mO����*�����[�2#*����*`z��_6���/_��Y�h/�5䗅r<����Ax��XI�E�C;\���E.���	�ڹ��,�ɫ��~��XLv��p@�`�<�a0��!���"F��٧��0a[�zﻫ|?��ˬ�V�O�U�X}-��i�W���Pjӌ^���E��LuFi�"�_>n�rMT�#���>ݭ�iR�/`���-yF��{p:~��al�z<�4���A阂�J����P1�7׍j���?ZMƺ��B��K7?��e2���]n�m7�KDް���w���4�DzA�����s����[����̉3i�%͇` 3'2*KN�����i�����,�	�1B:�iܟ�;iWe�ʟ!
'� �2���X��'/��q��U
LF��CG!��m��[�+��$^B
c�<� #��A`��H�(���dh�!e��	�'�����/_lb��d�&JP&P��
Y�{�kAG���û#���'Q4
(�pLƯ�e�F6�0���~���ĵ}dT`0,̵|�����i��������u�T|QuVwr}R��q��S�$	B���(��5��ͅ����p KYra�,Kt��.���Df�A�MD�J��W��/P���s�\��,5�E.s_'����ֹ�L)���)��WRR��`E_�>!�q���[�����x��=�-Fy�Z�M��f���jI�Y�s�����*f�t�K��L}������RoEL�����2׆6�dC<��뎩1J<RN@l�hE��F���JWt��_�t�<�L��4�	˺q�|�A��Ъ�˱Ě<�m��q�4�W4׀k4a�n��%|3��'c&ݚn4���~���+"4�m��_��Jg�m1��.���'K/3�j5�mԥ���	����Y��`e�<���s�QW鿲���h$y��z�P�l:J����4�m��Z����ީ�>�����Vd��_�C�I�M�'���d�b���fs��t�����Jp�Lt�3����n2�\-$\]���ЙAք*�*ڦ,�J��� �ĥ�N�ݓ�D)��:���~i��R{�����">��� �'߅Y�1lʚfg�(LmH�ERz�%��P���y�^��(��NߋZ, "������3ɏ쵬0	c�`��}r�Ғ\����.���_�{t��|�:�`�,��}���A���]vȏ��eN���/��>%���aH`L0��}	�V�i�$f�F�}x���=����m�/�J��1r<��Ӻ��L)�K���ä��?�U?����A���S�lB3�T���!��W�#��G������Y:�v7P`��co�i�Ϥ��ϡޣ���$�C��s�&��Z�@�H,���I��#Y6�yé�_�g�O!VA`r�7��y	Xi��J��2�\	A��hڎxoTU���44��	}e5�}rt)�<F<��^
}t����X�\�f��\���Z��3��+T�����CBQ�e z�VÞ!��Yf�`'o�_*��;Ar('���ʋ�������,��"x���!�3zU�HI�=����lFD@p0cdVF$!8����>q|�p��WyiY�64r��;�����Ǩ.��klB��"K�b�υ�1�+ �Gk�~ڡ�J����-�<�� )���<�'�k߷& ����`���dcJ;�go���Q�Lka�ɦ(n�Sy�~d���F�F�[Y+ٖB!��&bZi��{�Ւn��%4�q7z�氅�f�6��6�m|o�۸��ֻ��g�~�Bؕ��
]x��*��v���K��R	]+��\]�Z;�\�m��vӲ��{�:���MM�s'��OsH��k�7���o�׈�-⦱�|�������.�|It��rZx�z>��7�O����0�$2Vg\�6�������N�
x�\��i}� ]5_Z��Y����`0{_�(���!!�~(�ଳt8Ͼ;Y{(���hR���L;��XvA����N�6~r�-V���m�;/�𵬢��a��L�U����eu�����L�$�&{R�wo�9L�����A��\�/�WW��qҸ٤���HsM��ȓ>�D�!��GsX:� {��ťw����'P@#D�7?�7qT\��{¿)-��R�R���I�5����IiBtx��b	��p�Kt�����@�K��Z#mfwP��� f�������pP�+�c���C/d#��	Y�d~@�*)�'�
��G�����G`�kD����KU)$^Ō������7�f�{���d�jJ�N���n��[�e83��DM_��tQ��`�܄���6?Cm*/b�ˤ�_�nX���)�8��s��9Mp��/�����ܵ��*K;X�m�O�k�1}����e��M�/��w����S�X<Ɓn�Nm}|#7��&�����_1�rG\�W ��!�}"��ӚD\_�3U���pE9� �;:(�y~�Ł	a%/I	��$il/>g(N��jN=J�:!d���̬$ YmE?e-Z-���Lj��<��˼��J{J��g.����6�A��=cF���C��fE��VzRYf=�j`~0��ו�Ŧ'!��^D��C��"�F�$�HL�,=:E�w�4KN�����i�݁@���-%�f9��Lt��
D�d7�M�{��
Q�2� VC��j'�T�.
��5�*#`���`h��(7Q���x��8�p꜂ _��o�+t&�����#����tB:@�6�7�p���"�f��a���A2�x��g��M<R؃<L�u{����M*�;�Ǐ�φb3+�0(���o���n�ٯ��g[G���r{] ~�ho�N��� ����V<��J�<-\�0�gՑ`�+t��8~	��X//�6�9듼��*�o�2v�9��@Bfn�y7h9�Y�\b���^�n��q��#�|a��<`��R�`���:��y
=��� xyY��ǳr�{���Ɠ�['��6��`�(s��٬�u�I&�5V�B��jT�,����.p�������3��M�IIr�O��X嚟C���{K,٪�0�#�v�;3~)�K���4�7@�y-7�0�eyq��m_L��~�ׯ4 ��u��4o�?J����x|�<�O����Xk�AQ�u�s"ʤ�8R��n��&2<-�8�V{V�q�]�Cu��c�9�\��I'�����gf����Tb[���`�7B`_Jh���x_�~�V���M�V탾ڇ��.��x�Tp�����AnI�'p�\NN�kE��V�oq��v
�yIH�	�f�����a���p�o��Dj�u[�j�������j����5��^�7���.M�����Z�E�"�?Ek#�V�}��@M:�o�ul�8�z�@�eG�A!I���[�ިF��%k�w6Iݝ�k�̲v1l<�@�D˙k�uJ� \$�L}e�XM̣`��O�_�!�e�>[Ga�ڛ�sν@5��2
'�f�m�?<�r�n�]�D� ���W'?kz��w�}v��^i��B����9ȴ$Ɔ�o��3�Ƒ(bK�WM
nF�����'�e=T^�����!���~�u�i��-�1N4.B����t������G��ã��t�
�r��\�L����b��-dE8;l�#���Ռ?>�ɲŚ��g�o�u$I�([�H>mk�������	^��l�BU�.,O�v��&b`U�q��8��_Ѡ�{&R{�2��?��U��>�
�~�!kL����"��׆�����U��>�b1.Z�/��R���Z�g�.���Xd?f�.%9�)γ�
�$|d�~�z�=u�����d��-�bY̳bh�JZ�,�>BO�_��#���2�"�C$�^�8�>�B��y���Q~�Pv�[y��!���̪2��[�L��kǄǹ��"ef@�Z��A�Id�@f0��f�U�g_Kz튪���$���O�XZ�[���<�5Cܲ�����P
"%�����p�U�q)�489:F>V��C��v�]���m�Z[��s�yۙ�eq#)z	�Y<��!�i����\u@�!"��+\��FX�E,�Ќ&�Ҽf-'��b^��l�~E���E<bG�O~�+��(8�×gYjr<?/��*b��&Q�B��9o��;���h��ˠ��Ue[�������V�g��
C8%��h#fƞΖ�Y�m����ԜFXYTH/�1����ȓZ0�iD��|`p���B:���ģ?��H��1xL���䛸<�S.�H����H63Ȉ|�y�/m��b���n]e?������H��D������gͲ�7]#HP/��Hγ"�s/'�^r��j}�ĉW0C�.��@� �5�S���n� 56��'8㚔���q'�]f*�2g��)XH�����Lӣ��y�yR]�ڜ a�� ���7K�褧-�I���TE� �Ž��
�D�4������A���zC�%��9�j�fO!cEE�>����S��!�U��PVhz��<ÿj[Ŏ�Ѐ  MkYG�7�맣Ѻ ����St�를�A�:�$������;g��>�N�h�X�;d*ۋS���
(K\��~��>(���Y�5[��)P#k��c�Gg"��*��u��Uh�C1צ��:4c�+���U8PO�̄��Ń�i��1�#w6�n�s��i�
�Ad��`��'L(�sg��JT�z�����t�{|=��v�u��7����b|�9�ƈ?j-��&n9�c2��f�-kbu�9I��cY�g�ԚZ*J�R���&(��N3�.�E����N6��m�$v�<�S˫I�zku斀�f��UP�()^Ԇ�|q�-�� ����A���༂��l���͘vD�:�f�ߍ͠s��ӝ� ���y�ی`�b���t.k�6S���B��W�� A�e8��Y#�ɘ�j�7�i:��lܼ��R���{l���k�ܞ���g����˖�*WC��y�f��.�k��QzǮj ���ݡ5�e�S��an�G�d�f�o�F�Qn�o� �(%#��"�*�+��[��;0Y�im����x�0�Q;�� ���ȁ>��˦��9b_�_�k h�0�N�oو�g�fL@�F���h'�0<����R57-�d��4:�Y�⧏[�fY�Z�i��A�������G�M*o�啄�?7�]w3�8Q$��%�R�V{kxD������f�M,�w�&z�K!ክ�'"�`�A�/1H�k���2�șb'vF�j8ӂX�p$)�bi�8W��,ͩ>z�[�a�{�e6��� �w�)�'���z���i���*[�W�{J�9��>����N]g6�3��2��ᬼɍ�/����4D�\y�	�KM�5</ܢl���n���9�M�XL#�â���@gۊ����r�Iq4��l��e���(~�~
+-t}	��(p��{�(�d8��t��p�,�$q�a����vJE����N&�g�ʉ�߲�JKF�龝D؁#��v���my��*Q�����ڝB�ꢨ��p��������-��W��5m6�9Bc�\����Ң�DA��?��r�r
���*�v"�VF&�!�b �Tճ����_�7H��2 ����Y�a�����U�0mFR���^��ZT��l	;������%,��;�3G�TD}�GZ��y���˿=h|sD/�,sSI3�`�/�u�Mv��|���A���p���n�Q�m�9Y<J�ˮ�E÷>�(�7F�ؘeZ_DTTE���I�VUj��q�� �*I�c��N1�כ���	�'(W\g��{?i��#�H�Kŕ�%i�2��<y��G�%,cܧ��J*�f�!�y��)��{�l?��~N��q�g��S�lr'��HOli>��J[>Dp��e��g�̢cyDo��N����J�
��Q�Qmz�-����`�NIy�a$,�[!t�ب�!4��w�Um��ſQ�V0@�-

�J�x 2����[A��,��c�Jm��2�yEc����7�O�pJ!d�d�\I;0������膙�qv��I�����p��f~PS�o�:,)��k���l8�1�TzP�L���=j��0�s�3lذGKEj� ꦋS^3���ݮ��q=����n�%��>��+��cb�6���?��5�/c�9)|�޳6�R֩�٫�D��|<�7 N����7�b�T{��O�!X`}rRLGʆ�Iis�QY(��H4t�R��¶��;<ޠڧ�Л�!���"W��uaX�˭�{��rMM�d���X5��QZ�5�y!���v��̪'��>�O�n���� �ːx��Qo���ؿ��Ð�E��1qU)RVA��"��{��\�I�&����g���ύ�X?��q�/9>}O���pvU�p�ɛ�D������q̸H�����h�.�H��p1��(�.*�qX�_��
����(���T�����liu�������b� 95\xT$�������qt;j��Q��Q4b"d4Y)��'Q�2�_�����3�D	v_F���r������Qc��Ӯ�XCpU^C�P��2��v��nC.��&��qL�}�o�]Ӕ7qGx�+�ַ@Zm���_����Xq�.�!��j4��QM4���U���
�=�e���l8ݧw���Q��rk�f��@#�x��j:�R�FP�v�B��%f�ȓ��I$�}UX�[�Ft��hJ��:���YM��Zh7�xf޲�$pa���}v����t��m��B����1��xK��Ab��w�ʳ��~���p1�FV:�� u��>��~Wj��7G $&0���8��V���|��z�q�
���,Z��l���E��F��U;J1q�)Q�����}��;�,�V.��L�{(�Ro|��C\x��(������9������Z��X;א�.� ��[���~\��J�&#�_S#�m���CH�?Q������4�FX71�3�a����?/^��A��a��э�zI�	K�dm
gV%�I�6壒t^��HM�`�c�����m�Ў��,V���e}~;>�8���	��J��^��0���ž����C�3��/Io��~�\���^g�%��$(�;�tÎ�"xB��E��m>�q��P�4�#(�#���03u�"�0��UF��A�/�<�r��q�kh�����7Kc$b�3�Y̟�On���zA=�Waa��I1�a�,n]h�s�J���l9FK�5��1T�O�%���}+����.�w��^�o�q�R��[r����?@�ˆ�ߺ�r���ɴ�e6��	h�����ল��F��'�$��ؾ%�㜋&ߕ2�C�+Jq�k!���u� 7BNe��Oh	�dvL�qBL����O�x_���79�9FUR�������nŷ�ƌnx����Ύ��Vn�E_� 
8�%N��G�_�"h0k�v���3iI*	��(�=��$��<Zưnj�r�·�Y%�_������m���h�"wX�}{N�X1l�U�Tp�㵏S�i��+�-����w{M#p��BGL�dϋ�4x����K��v�jo8}���%��YS���o�q)F��ѱG��G���x�؊X鋴7��˂B'��4�ߊ3u�yx�@��^ʖ�U�W���-�,�r&N�K�W	��!-C��+C6"�o�<sb��#�wt3�~�1-&:ٺ�=���V3��J飥��}���Sh���N���'6Zd�,�H]幤�4�lA�D��X ��,�" 7�z|1��C%�K5"������A����YeI+ςN��M4t��,}�$�`���>4�6&��媂s�_E:��B�)��S�xH�G,j6���r[���a\���ᱰ��P���0a�����6��M|B�z#$�O�э?��{]�T�'әs��&kH_�û^�#�O�c�
gkX�
�E����&��kK�ռ�rFDw�U�u�΋�>�h��ңg?�n�0� ��&0<u++]/���J�!�f��3!N��_�87P.���y���hz�n
�����VW)Pw�x�"_y��B!!#p��Hqdn�ߟ+��~t�����K�~���`���5f�I9�v��RfʷK_�>(�3l=?x���b&�D�R\^���{C�Y��jEt�X���'���!��T���x孫���b�>[� �+N1�����b��w�bC^�w3G�-� ���E�Db̻s  * �����a��"b��ׄܭ���:܃6�#��}x~����і��y3y���,5id�ǿ>" %*���0Y�˶=��b�~c��Ƽ�[<<љ���J��g��{t�0�h��GI"�v��zMc����'ݜ�!�Zɫ;���x?��2�T�()F�c��[�xTƠe@jE0�����U�.]�8nf���en	r��*���˨��o���fj(������ј;p�J�����k���Һ�^���%Y��)^q�o��WH�CY"���x쯔��e�>�0���o��O�NR��mBK�-��� ��)aPK^�H��۽r��w��a���"�jG ~�I� e�H�Wt�j�t��S���]gtO�DX>6�FlTs����+��D�Y�-5@�,�Ҫ�l�a>��l='���.�T_���j��Tk���6���hzU���#�]N:��T-c�7r�:N��<��঱K�L�����?�f�jqJ�u��y9NoO.�ʢ2҅OL4�wp�M�<��a�]�l�b�opո8��Ǫ�j���:R֫�=DH�^��琨�&������8�]{T0�^m1���G]��8�����74�!�X�q��H��%��N��6eܦ�RP���i�)��5����g�=]X�Ŋ5N�I�e}~	Z~���?���v���7���"�uJm;.7�tj�CU���qOU��E���T���Q�E
D���)�+am�Z���\Xs��i�v��������Le@��#�,���9��."Cׄ��Zs帜I�cn���*���P��v;my;�6��(�D�H�'��a��[��F7N�#�5��x��P7��]��F1ڄ��!O�������Gwp_>0��}�}2r���m�{���V��ir�E��FRΫB��&��V3��s��u��g�����tjl�\������nĂ�Pr��Joz#��}�z�[2Ƚuᢃg��0��z��B8�'G���deA�IU��x�����g퇶�E�)-���`-��K#ӓ\Ɏ�%;��mM�Щ׮�*B�ĸ�߱���x�v�pa�ÿpk.��YJ��d�Va���T9���"_ �c_ƻT<)C0|�H]|�/5D�ݕ���y�q�3a��v��sW_0q��S�)ֿ�!5�m�^�2D@�O�{�[gΏ�p���w`�.�F�W�������C�\9_8߰�F��h��qn�n��R��M�����}#<�)JgZfi��S�@��ֳ����Q���(�������Hz��/�^N�샓5&���LS�b���'�6���Xfm	n�X�1����M�9(S�8��f>@��h6K�ܕ����4��~�A1�7o������+)Eǭb�g'Qk�ӑW�n"2��R�g�nL��f�	$�X�j3�|��s�~k�+Vù����V�ע@�p�7���ܟ@��{�q�aUe�C�Ac�7������\M6�/�H�a���~�����L �-B��[Z�u5�W��d�cQ���-�Xʪp�_y�"*�<��<u���_�УJ���)���iK'���AC>�+�fu�r7
�%6�p����慓�]�Ӥp��k�2�ϸM�����aW�#���Q9���X�~�r�l�~��npL�.9��\L�������	�S���A:OC>ÜM�����6�[�^��YE(�K�1<*���i�� �=.�P��PX�� %?������\ƿ�4��yR�πM(��sj�������yE�&D�1�ݸ�}�v��ʻ�<G�է� '7��T�}6��e	�����{�`��2�4��Ӄ+��c�w��Y�t�m��UtZ�UQ��G0��cX�@�e:"�ά�)J�	!VqO;��OK������ߜ������Ul��0;x.�ʦ"���.�p?���H&C�c^��ۂ��q���jm��l��Q�w�3O�j�]��! c�"g��5���G�yA
d'T�%R��D�����mo+
5 ��].J�؊8US:�.Q�)��s�o1�H3�88�m��\�^�����
>�N�Eg|�)W_�r�4^9���<S��ov p��7��O��Cy��վ<�@��/n������ǐc)�&K�Q'}��8��	E�(}N�i�� ?ε4��5�
�;i��:��)�Rd��j�u�u�7����u�x��>͵���K�C�
g���'�Pް�=i��9���%����C�ˍk��*Xv�dHd�Ŧ�#e���w����s�>����y��o�fUZ��v���ܦAQc �Sne�WY�M_�;�*eR%���g�����l���sư �`�1s��l�cb[^Hw@ّMi��A�����tV�����9�������>�M��1Lh߃��:�%d{9�[���T�[��O��i=׈����~����������b������-/d⭁�Q���]��`�s�x�D��-��sN��Pe��ʆ+�!ݘl�鿗� �oc-���]W�hH1�>�%�����M�a+"�
����ь�Uӿ�M�VQ0����A/GJ�� x��8����\A_�zNO۸�B���t/�o�C�"\�K�:n�ёr .�C�:����tV��i����W�p�М_�	8=�c3Yv��@�Ɩp�@n̡�@"�`�~�7^a��trA�J(��8fݓzA�ڼ�(�e2I����H����d���H�h�Ex����j����DsR)�d��W*A��^HTi��7��Rw��y�2���`��̱��!�C�rSN&~B^*:y��[!�����d��o�^�m"�ߺ��Irc|9�h͆M�c9L����F�0�ק��Ӆ�%�QF�>]Q���k1Z�uu~�:���n��Èt��d���*�A���PK	��B^�&%1���Eg�]�_%��=q����#�ʔ�}��O9:Q�XT�&*W�$/��Կ�5�N����eP+[��JsRJX��b 5�Wr��N��R�������Y}��C� �hJ�#�~�ܡ��d'�,jJ �[R+(��.(��f�s�(��a�t�4:�q���k��0U��8B�U�8� .�S)nb��3���ݱފ��l��o����3"O�Fa�Z�_?,b?�� a�˟�xy�\�@�'�3z�V2H����B,7����)D��#�fi�k����s��C@S���dC奏�D���$|]��v^�� v��Q�> S;𿺧�2h��ws����mj�:����P��FH�?�t��c�N\5 2;W��"�+���������c|1�r�p���������ٞ�a� ��B�sC���k.�58��\�Sl�U�|�Fm�1�W���A���љO�N����͵������m��n*����B~+�yUkj�fLR�a���&V�@�n����ʙu�T=�gec7��"�@����s��^�5�f]Jd��81�*�����j+�8D�����K��Rϓ�*2�Ռ>k�m�;YW���\�s*'�N�&\��N�F0,Wi����(�f��8�oȞ��\W��c���V���LO2{��e��ty�?���n2�X�$��q����㦰as��Ȩ}�E�)��������Z�Fm�ɈZ���т��LK@�D�=��ML��I��I�Ȍ �-/a��&E-H��w��'��H�@x��O�DQ#������(Mh���d��w׫C<�2;pR3��M�,ٛ��ˬ9q�P��OpVp�Li�8j�L;��L�~j^�H�0é)���Y�(�6F'{	#D�
�h�4ut��b(�~���:Z��՗���`�(y�pSIY�����
���ۉ���4� ����"8
P񪈐�Gi��439��$��Ƞ"��M=��a���3:�a��3�HB�(Pz��$m?�� n�؜0`�8�I
+�Q.Y�2�!��;e�:d�P{���ӕY��w�\�e�*�k�B�V��3��*=K�E����}Eۧ�ux1UT�2���,Pf%��:�:W��H���)BߡL�+̓����Z�ȅ�[ܼ1M+AU�T�d�N�kEm��3��EU\��ԑc�$㬹���}g�5�ڽ��d����AׁD�и	\�?�IC,��g=l:v���\N������p��)@����J�����0�<"H��`5�˺��*7����9p�4O5��=�HS i<mʲ�=�2�sY{Bf1Q��v>u$�>�s���ET�3!�6 ��<PR�ʶ��F���bj�j��(��Y=R� �0���JRt#b�1h4�Ԥ�������@E7��)��0��Wc���&/.��s\�ӝϻ�	���	�O�:�W,���������m\};��Rw1���'���ը���Ԋ�ë́$�K�80.Ŕ�=)�� )��_	ͱ���v��Q�U�����p�V{%�.t�����gx���!(;�Ѳ���$����w[�r��0���wh�����h��+�x�ئܺ�E���:��2�*�*�/y,جW��V��z�
N/՟����Q�6����v�ˎ���^Į���(RnrT�}~2<�j����
�7��I�;t3 n���.�1J��J����m5��,M��<����x$m�SJc{=�b�J��p.�"s�:n��:˝Jg�H��c��:3�����8P�g�	���H\
@k�t)fJ� �����;�n>��=�͑�t�֗g�^���pr��B]ǠQb?�E毊j~��O�&�{�8+6/��8s-�����x�ReT�~ݰ��A_��4ғ�sZ5)3�e�&�N�W"�׼��#��������3}-����G���DpR'�65��m�7�r��U�����3���c�;i��i���n�ȥ�372i�G{��i�	C�r�P;|4?>{�o;�?���}[ �Z�j{E�}ol�	�V�+�fS�����a�$��f��S��tA�7fÅkQ��W���5>��i�.�}S����#RYB���=��1ˊ'�t�����kmt�B�^�����-��9��H������	�(���Г|k"�����v��.�!���!�C:�x�����:�� ��I��^p�T��m�]��@�c+*�ݿ@7�B<*��u��?;����/c��3�3��-��Ĥ�1�F�@�s���?p��1a�k��lD�W�Z����r�.���n^�QC�O��
�CjXG���d��Z�/ ���5,`��ǽj�.���H�YJ5�-ۙ8�(��k��7��9R���W�+j�5b'ߙ�`��vA;�rt�J��vFtv�H��OR(	��ʆʵ��('���og��fME����_�?��f������A����P/�d�q�b?�KR��,��I��z�l �O�q����'�6j��l��g��X	&�Y���):�8������V٩V�� ��s��,sw��o�USb�\$a��|N{�Y�_��߻�2Z#�<:1B:�x�՚E�xv�o�T[��[�Jꬕ'�)�f�)�Jf�(��!�� X{���ܩ�[=x��2�G�7��aݓ����D(����ЫR�hTV����ݶP��YH�(݄5��朋��	f�[>TR
�K2*��W�������bdr�)�kHOj�Ʊ�죌�� �c�T�$̓�M����ţd�sbe�
���+p�2����O�S�0H�!�V�+�HW������i��Q>o�{w�!'d*�:F�e%)�6%>�Vm�/3��>foOl<�y5���z�T��Erc<w�'���ol��ZQ��f}.��$���xq��}�� ��͇,�Xeh}�!=�7_S��o�%��?�ǹ������w��:]�2���L��]Q�S���I�Fn�R�����?�;��A�7g%]ԯg;���,���9$w~��tC�r�;�Al��z�Nv�s��
U�T������bJ.k�=v�X�0�YF�5b)�s�J,|�R.��@YSj%8���1��ԏ�T��hED�C��y^+��e���Q���M�y<��k�}�*xU�{����P�y`��$n/��B�$ ��׫�y����&���J��Svc6�v�+���������1�<�u}�ɵ6��"�Y���àzhM�Ð@��S�������������A�C�hz����Ӏu�Kg�y*֏��^�4�R3Bq<0�V��@D����p�y�q��Q�Kx����e���6[��n�G�-	�Q�7�P��Ye���+�9�Yj!�zi�%њ>��4.y�"t��V����rA�m����nYwX��?�/:������?:K�x����V�z� ���S�H����\y�~F����r6�e�=���G�)�"��#�F)�*��rgi&�EL0��I8�غà��K�"�
�����"�1�u��d�ic^ �5��.8jB��.����X�,��a�t��!Qn��X��$J��^A!˚P|&�k���/�pqz��Ϝfy��� ���N�~���'z�u��z��¶(֐��{��:�Ƶ�y���@�p�6��s"p��怔��&q���C�ha�>�˔AU���Q�K��&x�_\�A���)��B�]h|�&܊�@e-j;��}����.�w�������"�+97S�d�X��-��� k}������n3ail�)�y�r��ǁ'%^G��d&V�=��*���y0�G�J�/֕�T�^H��w�EB�E�7�b�vZf��s�xB	��Y-7�m��F��גym��U��n��W��A�56c�		��q��1Qb�Ɨ=��`��:������ރ+0���C��p㒑�(��S^��y>�]�5-� �?��xj\o��5����6��-�����ƀ�c���C��\��%�q�;�Q�2F���O����C��
\�ds;���'�]��jK���G��r�=�������55�VǓh� Ǐ�Y��"��B&=�XC<쐲=�y�@�$�I�k��a�(2�_��^!s���-1���_P*N�6�B0�2w�#��C��o��{}��2I�͚���{O�F��i��Tu����PB��M!(}�X���U�����.��e
�FZ�-�P4�.l�Z�럼�*|��LC"�l��W�&��p��>>>=W�����Q;��!v�u%u��`ba��fo��Ù�/ֲgR1���@�������Q�B-!��%>�.�P�w���O�c�Gƅ>�-T��L��V�:S�η|��=^�Xt���(�D2
�c ����a��#,&�n�	.]� P��S%Dd�F3�2$�V�!pn�έŦ�k8�ú���a��G��Z7G
�玼W�nyd~�]d���s���6(i=�x
��F�JzG��"��)��s��#�;7 ,���m�F�TqM�|��H��rwk8�/�D�Cng�wI�U�ٹ4����W���Y��Ex��;�PH&�aX��r�(�6��P��%��Z`5*�:�d69\�ᐆ���'�+�1y�b�cӰ�"Ķ�,w�o�b8v��b\Y�M"��&R~{G��X?�"��9B�1�jFl�'d*�n�L�*U�4<}߯�ڭ�Fb6���hDcЦ��:�*7<9 mÿ��4���h<����&�\Ɂc��.4��� ���ޛ���З!	�A���1	ϝǗ��tj��(#����b*f���rpwc*�^�ͽK|��0�W��[�
�-�Q��T�l+{6&��|���ё�A�hD���.>��ݟ:�@���JM�ek��������/��:��ޯ�h�J
g����°�*��� ��`�T��`VvJ�(�%�(�"3��?���������|���:�/�,KEq]YU��@��՘"��Wu�_�����܁4d�5�x|oq��P?��y!::\���)��WU�g��#�sHе4�0�斿���$U�[h��v���%�*��1��
i��ɇ5�̗�Zb�-�o�!'��G��a��ymV��BG�"��#��Q��v����ꒁ�w�<Kl�*�%�1�1m;.MIxѫ�颳	j�@�Nѻ���T���d�̼օ��o#aP��!O7w����q��s�;������h���mC%=;!Z�\Ӓ&Am���xOΎ��<и��i�*�ǽ�	�(��� s#]|�c,N�4ʱ�{N�+1��$��oEX����o����{4#�����AEe#�7����ޗ�e3'a�!��
��f����<�Y�ޓ"]N}2��5޹���7�ﻡcݥ�B��|�Ƽ�$�N���حpAC͠�EU���8X}�k�6�M�!���0�{��Y�	�l�V'I��xl�I\�@dav=�Ț�4�S�NS��~�l9�:y�\䖧vn���*���5�j�H�g?$eO��%E�z�����ʑ�/��󮂠��h��a���֒\�������T��ȒYy��$h3[�����#�`VpH�ǬW�\�C��S&t��6�τ��7	�B�����7e��X��� 7��$�3f�W�9W8�� �P�C�R8E)��P��e�]&�~faȡ
�~��+be�K��+���zN�S *OVN�ad�!��9��U���i{_�E�Q"�IV2
��d�e:����0,f>Y苰vGd4����Xj}Q�*�n�����><J�-C����y)/!�Z�!����{�%��[�xUx̦�-�["�X�Ǣ.S�eC��i�5yG�;s�R0ƛ�G��d�a& )�F���~T��s�V�"8��|bx�L|���_�>�^7)�DI�2�dG�sv(������:�YO�9�Q����õ�Grb&��{#�=A�,p3������-�1���kMV�T
P��Wyj�/H�4�� ������h��� y�=����`��P�����Y�$�=�I穄�~��Y��̓WA�?�4�q�֋�<H�'L�K9�����+1�>�7���]�P\��n�������d�y=���m����B�F1Wԍp�=܄Q)n��r������1�S�2����gQ:���=�� QYr����!ߖ��Cnj�}}ؼ���{Ǩ	��09��
^��T�,���rLզPҫ�?m�Q�ѷX�xtƱ���vq�J��!E9�i�V�I�_��'+���?��@�in��9��\����&�Z�xd��Y@���z�t�@r6���.V�*����Šp�=�8���b}�6��q��ҽ^���$��>��|�FZ=���}�~����
N�X�W2��+K/;��s��u�S�w^�G>Ҿt��SW_�R@���mR'e'��7p�\��f"a��Q�b0x�%$�&
P���6��è�o����tIu~>x[۱D��
�S���(x�)��s��z����[��:L��B��$,S꥘�9��BW�.���'v���f��5.��q�v|�选Gmn�䱸�桶�V�7�ہ�e�Cb�p:�Qr�> �6������eqY��.N:t���y����	g�$��L�E�[����ti�s�Y0����d�/u;����HpP\K̤F��F����5��_?�﯊�Eo�0�ؒ��'k�R�[�i9��S
U_��oԛ�����6O�>n���f�f�:�&�`?s���O��L�9�H⿹i8�'7Y�t]������Э�~Yh(���0~<5�u�y/�p{�܊��_Ў��4���䁗��M�(���^��a��-�r�6