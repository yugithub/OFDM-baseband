��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6�0��a��جTEٔdYc�~�ˊ�+����'ڌtV����bT����+p�k�NȽ0���
��_��T��˂���ϙ�=�dFN1�T��j����0�I
W�*+![�܀���==�Z�#!π%~H�1���&Ev\����¤�$�����}��I�G(!���B��/����5�'{j��i|[n��,�m�����[Y`~٤�M��( 4NV�yZW�HK�a
�6����JpP�D�^�d���,,��H�&�E�H$����S�5-\?~�[#�����-J��B�o�!@���kI\�\����>$D���x�G�O��ו|�R;�I]�ٴ��u��嚏������I�7g�}���]̭���m���+l���|e�1%p�F/�uv}z3��c��E� D���I]Q�}�hh�"~)�b��r��2����eS�5�hdJ^�
��նd��k
��w9� ����Z��Y�0Ʒ�mഷHt�9�-�����n�a�eTf�����c�&>
%�O��UXIE��`r��K������>J̙F��M�,�Ӎ6��'ic��)����oOK؂~��"�<��#S"%ֹ#"(_���"�,њV�,�.�LY�d_������z 3�Ht�t<l���H��6֫8 ܼq��r Y�.?@2']ōk�z}罅�6Y�:;^�؀i1�2NN�-lN�x��z�r���}�L�]r"� ����O�E�q���9)�/��؁�t[�/U��W�N�>�t�ܸx�@��z&q�G���l90�#b'|�\���c����0b�_��U���9��f�2@��)�s�GZ��4S>)��P�Q�q�n G{]�ռ�%@���~���-Q�!&{K�(NǙ
�@�8�
[�5�^1@�v7�.71���������`e
x%���x3HP~�m�L5e���9�{�.�C���y�S�Y���B�/&�,�TC	*�$K��n}��yc�p�����~��9�0g�ݗkо��{�������ݑC�O�p3�a���Š�yٙ�52��]����Z
��"8+��pE�ܧO�c�jl����X�:�`��͑�|P����5���T��NnɖLD�6��̨��Ռ]m*�܄z[φ^/�;����Z�@�z�b����!�9'm���L�y�!�Iw�O�@b��<r�^�V7j��5����L6��#���`��d�坄T�H.�5>�3\���g���`>�LI��2��߷��b	������¼�Aa��*<�y[u�X��a1�{��2��z���`CښnƠM�~��" ������ yjJ��&I�����$X`�H�g�or����|}�3��g�PG����i>�F�^�a�m���$	�)HA�O��6G7����z^R ��g�h/a7��8��U`^=,/#�ռ��3�%��!���г�&5�N/��.�H�UIz���b����B�H"�V"���3�?�D�FjRYx��-Hw����}�7�g��̑*��VA-v5[X�Z�{�����Ջb0YR�3 ��������4$�5���k�1��:MQ�-�@5���Wv�4���@S�R߶�,��D}�^�S������'�Ŋ��c�	�K?�'.��4i*�����#�A�g���lT�A����v�d�v����"�uOt�5f��Qco
��]�,��6�U�Z>FoQ��]����ɤ����*i����K��Nw� �B ����'�1({�类�:[{_���%��~0��*\�r}c���� 
�Ӫ9���I�������YW��3S�=ufZ��Ղ�u��"��A��R�yr����q=���o���=�hD��x��G��},,�|���^�9Z�ެ���t̫]4�E�K�z���=$@��q6���W	�O( qick�Ж8��9$=�u�I6l/t&��l�F?"i%��8��7�qkfh��\�甬�o^ֻ�5�N�e��f�7��[����`%s�P3tQ���dZwKnV� �R�A0���Kc������YQ�y���ܯE��#�C��}-#Ֆ�	�-n� �Ѿ�}�s�乘74Y0�`*����%�'�A��5�}�4�u�}�m@���I��h�E�fǽ�J'��(��oF҆(�ܶ�cS�(z�>�$n�]Η�=V�<-2��n ^/�x��^p���Y^�'1�_���8��(h�d��ܑ1'j��]���$yA��Y1	�;�1�k��[ڙ���h3������z�Ȼد�(���]Zv�,^�k^�\�[�oQt��%#>�H�*�M�J�Y��6W���N�L�\�Q�ڈ�H��޶�=cQm�;6�fw�7�j�y]��U /[�zsP�W��gS���V) R)�����H���,�Bn�7ܕDE����\Fސ��
\a}�_<5��QO(���}��%��|�QV<��\S�-Ѝ�ϥN������dI_��4�0A-p�kdͮym�6��b�*����l|7����Y8��a�߼/L����e���F���O�(E�d���T]�:=��d�bs��n3��@a2<�KvB;������ŧ���)��i9����j�m�I2��f?IٲB9H����S�Nm�zP�4��q�%|B��A���bfJ�E�ڮB	����3���'�#R/������nG�� )�p �A"s��g�� ��k�%�ã�RW?V��aL:ܯ�w�q0b\t��7��P�Y��]��oO��1�z�7��PG�L�4!��3 iy�J� +���VX�V��&��v���� &�R��>
V�����|X4�����\..8��&cO�����:����}����xઉ����>&��|o������]�T����D"Y����ߓaD0=\��N�̝���AV�|��.�cdu��j����LF�	�d�E}���m��_����>��^a��X�Z�;�+#m������b���&�prpr����
]|u�7��ti�du�RB����ӎ�O��f��&�`�m1�D��+{�L�,�X��|6MW�����6�zM�6v��&}O<�y�9�Xu��}\WNa���{8	+��/����*���Ӏ��
��*�'�ZqU?�!���MhG6�=8�����C�m֍����0����x6�V�a	���6����8���}�r�e� �m�L4�<
�&����9�
�C��¸0�GZ8v�p���R�H�4  !e����D��ٶ�����:O�������N�=Lҋ���{Hv���T���fL�Z1�'�� ��~8��+k�ݮv�q�x�2��Z�h���̪��t�.0�ѡ��+���%��{>�q�gmp5�
p��QL7�b�q���`,�kaz2FMG�]i%���uH2�����N���+P�?��z9dWXx�8A݆�+�I�H�k�)n~,�*��#�,Ӫb�d����F�=��2�)5��n����O)�ۯ�6!`���o2=����/7hPX0�Q��k�������-yj�*o6U���dH3g�� fIqd��L�V�K����d^yhi#�{JK�<���x�:2:�>��15�����ܜ� �^2���4Dz ֻ�X���0ev�s�Y�'���Y"0/���f���@�x������g1v�ܭ�����1Ρ���y�H%�c�ge��Y�8�q)	}o�ψ�I.R�~N�@����=����;���_n�x � ��}e�#PN��o���?{_��%@+@�g�B��� ��8�
��3�t�=������i ���S��H9y��ltT^V��g�i笔�'�kq��9УD?�j�u��mM$���sb���i6(L�%�ho�(O;�]����/�A���s�"%o\	�6���}6 L��V���XV��zA��U��&�	�׮Ny��D���ΊoWHf�K� �/�v>`d�Z5��Ԭ�-do9����'p����;��7�R|�K�#%�G�~��Ȭ0�������>�2N6�s���M=�5�bu�?&����r��`�S����l�e-�W��o�w���=�L��_>*�^�Tŗ��������`�Oa��<�1`��׆,{l��W�xP��H)T��8�om!=�ԟ﫼Y�i6�*l�p
�vO��1N�CPi��#���������vS���H=}	��=X��q�h�%pKr �8J1"ԘE�b�}C�Z[�S�[uum��ж}b�@�YF(�b��b�$���?XA[SEɡ���e�!��	�Q������y��+{'1`8�8做��L�1��PT�h�{V̨�z|���|q��u�_1�����q\v1Z"h�H����mG�s�V�5��
ZTf={M��_ʹ�W��åIGT�W��)�լ� &�4߿�]�Y��F������Ds���b�ix�o�6��)Ҍ��J>\�\q?�ބ���ߊM.�v��z��U��q�X�U�u�;��0k�讀b�ڋ�z�IhI��!6q�ä���#+�=��t������m|�_�X����A��}���n|'�=�"�b�y�k����FI�ʶ��{�e�,l����2�~�e�^�O�Jw��ҍ� J_�J��i�dq�K��)�CLJ^ppRw���&�"��l�7|�nhE7<�3���C�b�a�n��40{V�w�jQ{�"�Cz�԰��T�'�~KklaM���eH{`��\>�r9����<�ޝnu'L�#�7<6�����;�t;GG��M} ����?D��Ekd�yE���	��=
2]O��l��L�E�-�H��`{�[�"H	�!�3/�ux�ou�Ӂ�'�,mX�J�4�wD����v*D0~�z�<oo#�L�"JG���[�Xh�tp@[7BD�K�Gڳx�]
Y��{A�<jX�����K�,����Q	~�����!���/�Aj}@��嗀۵��F��ԛ�܊�L�M,�'F��fJ�����rڌ�����C;_C����`�x�r�;x�`��Y	��^Հ]�7_��c#�J�D�
���,<{������'�L��� Zdͤ�v��?C���f�,64Go�D������:���^ �?գ�E�].���>`�� �����i1�_�:C�!F�L5�N0�i�>ð��}�� Lԏl�4���������<�f͹�+ 뀜���ks�����j�/N���1�D������B(i�y,��^��,�\�TN���=X3�/��=��ͤ6�7Y�@��;��kL]7\��X�:dc�����r���-"UԹ�B��2�<�s��3�����r�F��v�V݉��h�m��Z���H%dy��k�d����w1��iێ�6��f�|�����ud���	�H��8��DU�(%2m�c�7��h��i��i�Rk���ܶ~U6���9UN�O ��\N��^ф�P�J!%f��_c$I���֞�DB|�2���]@1�sM$��}v	ƋL�GK����Ge�ir@7����L��D���><���SCS�x����T�.n����x��P����,<�S����S}$$��ҙg)ٍʐ)��eX�Cqgᬃ��n^Q�N�Y���Wg	6��õS����i�y�c/]����|o`8/�%ÓB�>������}���麁��P�8�<\1�0��s�_I^��ګf��/~|D��O�H�����1������� (}�c�<sD�x��9���}��ښ[�nI �3�N$�m�\��w��Ae<�"�`��~P%*�#��١_�\��'�o�	�t�ܐ'���+�]\~��h�8ݽ[������38�c

�s�%�n`'�r[]��ݝ$������'�Df�"�n�Q%x�� �f��{J��ـ0l{#��̆�H�q���������0�����]���6�?�����T�'�*ܼ��nb���cF�sB� ��w��4fh���;H�9���cY��LD���8:9]�U�@{ + =��R_���X`�N���q��0�5�6�S�z��M���=�)�N�CE�������T��	��t���{�����HBET�*�')�G��q��A]g��m�m�Aw�Pl�x�=4�2RH�7���U�_dP)#f)v��A�U�}T��O
'ZB�Z�1&�*��S�Cٿ���Dc���˵�譫x|�faw���Y{4|��Ӭa  G�ہE~�� u|}Y5!��Vo/�t�r��mvS�\ָC&��J��Ԓ�w�8��Rz�N�_�V�ȹ�C�Y본|��F:�s�.�����FyoQ-��7��N�!C󷞗^���)>��͵�F��&��;,����{�p�N�Q��aZ�G�V*�9�T�U�Y��v4R�w)�8��,T��V2B5�-Jk*�cEY��1$��t�=�����j���D�PȻ��3��;�r�s�k\p
�v��dUqL�9����q�Y�f�.�)�ԧ�o���U��ߥ�(EJ��q�n6,I���'����k����l�b$�>}��+�Xk��W�~<��c����%!�S��h����r�N�E�xn/K=�i�E���_�r��{OO5��A��_8�v�#T��4���1%J{�ȳ�E �JCl�:������i@�H6����]7�Q��^�r�pv�+�V<@W�и�r�/�وp�ޫ�T]%� !of||,'N;4��Wԍ�'�Y����T�	�k��M�Hm˦#"�
�Y��Hc;;?����"C���y���Ԏ�}M��>�u
��ǿ�ϗ+������V5��i���Vʆ2(2:��&�
��n��<��6�;�@~�%�������j���w�{9os��)�L�`2y+�l�7������{��c���@�E���zF"�P�bEi٥]�2��/v����/����.����Z���G@�B��}��`9��Zf�G�dbo=
��ܪ�5B�G�0��&�eu!�?=��gC�%Ow5�����}�?��R�j��[{V�nHjݞ���Lpe�j!>��l�d\޷�C�~��ڋ7�}�]ZG��D[�s��CҤ�XD5�m�=�f&B�W� �D��dnm�g�=WG��5�����DO�F�D=5se�V�X��՘}�h��ԯ������/���D}�V�L����C]�(λ��ؐa����|~ܲ�.��u��T�� ���i�n跍B�P�M�lھz��J��5q%H*~�/h��.$m��g��g�,��a'�^�^���=+/��Aw�=q���Pv�d'��D��bR����z��O��^���I��bT���������ݾXį�|<Ȗ%�K�y����GH��M�ۋ���.�	�3"뺗f*Ӣhh�����DJ��-I4@p���;��h!�i��G�TcH ��n'�̀
���,���mX?);��ݖ_%�c7G?#u�����E[�i<����A�q�x���v�߬���p0��U�P�_Fѧ�3��'�Y[��'���o�x;�@7���޼�cZ	����s���x�.ֲ�·�(��Nghӆ��|E����%��`YQ����gU��4t\�ܓ�DBd�jߗ>�~rq�ƪ?D��X����_�p�����D��:M��Kii�9=��!Y���k� �`W��-�bAA�R�E�㩞@�=źd}�by:j�7>R�-V��&���p��կxQELveH�-wA*�3�fZG��&@&�y��V[}��}��s��䄮�>%��m�d8:�\/�3�3P�+�u�%��&X��B\�]	��l�B��2�"��X _l�kf��P��N1~2%���|B~�Z�׷�Sņ������U�\<��Н��Ҝt� ��������b�`��ǈ_Ǆ�C������cTA4�/\��ȭ�n*��`��<3��)�mz���TN.�$h�O4��i�Fݷ�g]�?5$��D�<]T4���c�O�����K<�\��-����;���BOu^2���*ˮ�Q�˕��x@� ;p�w�H�vC'��L31����	��jb��5�w�԰/k��ş�T?�ѹ�
8��-,Z-��6��{_x߅�@\ ��u#_��r����V��H��PC��Fo�Bv/�ƘA���Gy����&��dۇd%�����SY���b�K��P��!f�����r�L#�������W����?>P:�z�G���N��C$�7�����[H�b�>HP�h�A_��J�!���"�)�N\e�Oy"�����E�HeI0���>^n���q��'�9�YDHQ��$v����c���_�B�������;Gw�F-�|�
f�þ��H`Iu,+�!rwhm�IW�;��2�jd���W���uY��;������Lt�Pm�ʲY�Y(z�w<�Ԍ���� y��R����~�zI��?�3Su͇�����AN@���4��T��0�P�����N��
�	O5�h\�k�=�p*~2�g� ?������Th��C��Tf�!��Ɇ'tF�:�sS�}%��Oi��o�e�N��dQ$`�R�"g�����yh4ğ��h�Ҵ�w{��)]1�ꅹ�(F���iK�q�C����!��A�������9����s�d��/�(�5آ7�F��3�m)qΟ]Ώ�m�sn���#G��J敨n<+GP��)��)a�P���I��<ŒQ�{�F�l�lN^�V�\�O��S���79�6�c�JW> �D�v�W�[�/)��
{��)�7Ȝx��a��R��*��/�qBY�g.�x��|і
t\��R���w��ӋR�L�Ƣ�X,���4N��������2��Wl78}(%)\}t$���I�\�są��ϠKf�Z'zT|"Ln����U�]@/�a�2'�f�
��y��ᔅ@�Q{|I�*�0آk�j��h�zY"���
S�H�c1��3$"R��눾z���:au���7��À������B�0*3-��!����hj(`��$k�×�b�|>.[6��e��]��bm���<-�|��n�!P�	9U�ݞ���@U"�:�<������M͇�gS��5��s+iTif�V1@lڂܤ�QK�8&	��rհ�,-v��ؖ��(�a�'CԘ]:d@����>wz@�T5��T!��q޵u��p�x��!ʤ#z�TK"#�������v���<^�i��$k��
^e\�u����Iya8�ŝ���!9�[&%JN�ė�.9��6�х3���%�8�f�O}����)�K��S5���Y(>Ū��ߜ��τ+H�i��?3���� tw�"ՠ	�M`���9J�O�n�WI��@8"o�9�ݞ��^����);ig4����,��ՏybnΗ/���+W�>���j�8
��)B�,~�]�L�̥w��E�H�U I���!%��9�7f�f���q���%*�@�(�=��̌��qfQ?�"��n��CrIZ��Q/�RNs�z����k7��l�U��*��P��
���ja�s�*�h��N�O�p�.F
?��e�0+�L�=�i��x*}i�*	�Ϩ��cIs�@���M{�K�2g���1����L����0q6tĠT�j�V{��v#�{lvrՖ�ƍ�����@BƸ�J�h>HJ�/\6;%4�LwJ�ң[8��a���
�/����L��x1c'(�fӱ>}��QH�%p2�l��p݂'�LD�`jq�T�2��\�l���������D����-`������!��d�B�ڰ��g=]�����T偝����E�=����A �S\2xnfX���Eث~s����3Ӷ�enݙ���p����x���Z-�{�Ca�R5SD��BZv��Aj%v[B�p�8P|$����T��=y#m�S3�q8c,h0y LJE��w���
b��W�`҇5D�����h�j\��}<�Y��RT'ՠx�?�&�+��e�B�U_�[-E"J�B�w��8n��a���Ų��
�)�y,�Q�&S%?o�a�PT�b���Λ��3⛫�����-�v��`!�#��n�M<2wwA������O��2>�����;%vb�X�D�d�Ѹ�Z���Fҁ��h��Kۖl�2��/!�"F�����;nƎ��}�w��V{�����Ց�Zmd�����w��'T��SH��M�|�j:���\	ϼ����w����#yu�6n���L�̸i��u0�.d,�Zk�>�̵ZjM�������p���`�;��c��q���p4"��3�J��+�8 �/�D����`R�+��Al�c�Jl�t����M�9����mM#��&qn��
C4�Ysi�ũ�qJ�p��D��3*��X0��&���7��语~9V�M+���M+}'l���h��;1�'���!�~��P8�E�pK��ӂI6����%�\eC�e4 �↪ĥ�h3�HA�J��Bx�
c�tF�_)�E�0Rn�#6?�����������<r�H'��g
f��(����BM��I�SC��?d�� �������i|^��A3�X�(߽��_v��!.����v�겔7K�5䰈ͣ�k����!9𓶽]�y�H�׆ h���H^�� ����pO�WL�i ���0�HiSx�5	�A��Z�t0u�[���-�.� .5Q�u��l�m~'�n�n�s��ߚ9ϝ��������ȡr�NEΧZ<�K*�K�5^2.�-�n@�u1�"���Am�E����CFeU�`����--͈l���ﵕ踰2\b�h{������>��f��t��1XU@\�ekWE�ap|q�@��J�B���go��Kק�����O��w��Cq7|�)�?U
� ��@_<�L�{�¯Q�@K��+d�@@��q�[a�1�0ܢ�=��x9������[�|iкuXL�?���ծ� ���
��?8`�ߊ�#��=�$-o�{�w�������%K���JX���$����1������ʲ�H�,��
�/(��x��YJJ���������=�R��
=H���X�0-8=�~����N���x�\l�٩m�ʆ�+�C��*hU(����xP�q\kJ�!}��߽�ӯ��*x�S(��@@>��_H�3zt��ps�"<2���R;�� ���D�t�(��>��h�W�2\J�g�,:<V1�Ec������{oS;Q29�����m�X��ٙA�_������j�'���m&�"��Hc,���>p�d�IX?��S��h���>���PQ�l�hF:R����le��g�}+k"����n-tN���*v{l�ef���d��lH�өޚ|*k���{����r��Q'g���J����� 0������-��J0�8b�@���[*L3�F��r��*����L�G�7����MA�b���O�G�5�`�f�5�?�'��GT��'�mS5���I�.�m;�;��;M@��ѓ�;��@^��Vu��(�`:��6���}pn+�B�ju�9�;H�Y2Fo� VlBq����Log���:ru�'��*G��2^xuR�:O��W��vL��h����T�"j:�VP��G$t+�6O��1����gx�Hp
J�4�����3v��ϱ��,3����I��4c� �d��� �W#< 5�~e[�D7��LGS7�
�^��Z%�`��R��bA{�Z5�yO��������v�8��3���~Ck��v�6�q;&�p}��1˵+�lQ���"������s�=Į��^�a�5�Uv��ٹ}����R<�����?�{��#�U�/��c�0a5-��g��2H� �R'��\#l���E,��Y����?G�Î�^�� ���6ُ�w����펦��h�G��k��Aa�9��B�o�4�-#�n.�A'Z���}���ҍ7���|�aW�2��=ne�"c�6Ĕ� ��
�z@�G���ig ��Ȧ��0 8a�ز��im��������U�{s��l�������QG�Ƨ@+v� �rP�WI�6�7�8rQ��l �pL�se��+Ai�(r�&��%�X�h������(
�AH8���͟�o��F�;;��pѣ:Z|>g�&܌�5�����(�8��sf��AʃC��/������:T��9h�ȯHx�8�W⏔�(P�sqE���
�����U.{|�Z��
�)������0N/hb!q�����ߊ�������N@o��Aa���l�D��YV�Rز���x����S=��1ݵ��@��P�U��ۤ�^�o�}j���!���J�/OfG�p'̇3��Y��{�4�:���
����c�V���3̣ �_����,y~
����Ep�z䜸(�o�dԄgn��5}lv[�h�l��m�/�>��sse`���8��Tbբ��SW48��/I�A�k3�=0����G�B��h�з]�k��7��.[ʇ��ȩ�ꉇ����qƞ^Yg�s W~M�����(�r�������ԇED��p��-|[Ҹ�3q�~�rk'�i��@��i3JPs���+P����±*�}��{���[�Q�&��#S���C��;nTk��z?Q�X&s#��o�k�ӟ�\��&�:|Z�����Zo�ou�s����d�j6���:t�4��_��.8�_⪡Ϩؘd.���*�8�7R��Pv�Ґ&;����n�CC�P_Ҕ4�>��h[Jdw��p��Lfp��}=����	%ъ�lTA����Ā��"��ǆ�k�"ڍ�,�r�8�����V���?	�<	���?h����;w��q��� �4��q:kL��LMS��8[�8�uT�
�-�F�a�NՏ*��pC�{�r�fC�&� �V���zz;,>7�|1�.a�t�ղ���׌�(�b
�;t��иCaZ-&}�
��r�}�&���BW��G#�����ĳ�h�[���@�u�M�d��kz�4�������bJ|ir5	=�ןf�������J�Q$(���L��#�U��S���M�%4��4�ڭ�����N�\���l�H�@��MBe�b�e�s��y5���>W�'i�g��nK\D��³B�g�7��$�\>g�j��#��յ, $'�D�@���Zz��׭\����c�Q&Ծ���K��p�(�2�l3k�..<�+@R2( ,/��a��ɬd��<}
sJi�Ӈ;{���P��s!��h�����F(n�tݑ�"Z���%cP� E�TS1�z���~��\��m�4A��(xK�!�Ӹ菦�����ҝ���<Ҫ`�h�z�&�!���-��ŧjlF��'V2��\L=t*vxm,����~��W���+��#9>*baA��
����-�.�M����Ad�~�0^#�*�4�Y��5���\��}��6MI�؍��wٌ�u����)K������/��ڪ��|��?-E��h�#�����0�B�A2�-�=1/o�&8��ԑ0�zJ���i���DYshR)�S�aXA㻮y�(�d@�Q��R�������Yw42�
����:��>�3�~�F����pB>S�4F���I�/�l
L#�|�]�i�>V��.�Ҋ�8xH�,����P5�wQ�;�/7���m��j��//���\3u���T�3G˨��p��ѭ:C�x�%�wg۬����Rv8�=� 3f���?({HU����(��/a\�'~����bސ_9��T�x*��>-����ؤH�g���& Ps�����.~�N���`ߚ�/��,[a�5|�;�";��Vӱ�ByIb����������o�y�"�;��3�X?�Ӄ[��������X�9�x�и������R��B��C0YW�X���k��v��m�@��V�bԇ*J_���ۭ���-C �峘��f�qa�����l��'v��\|g��ަ��-���VgSd�TY��~bڽ�އ- ��f�F��5&��>��X��MF��_�SNk0#��3 ,�%����&F�p0����Q+z����1M
��qu��r�}'�&d�Ű:,�+WD���l��8~�E9�ϱHEP(h��v��GghU�6
i��a�_6�+!�tM�8�!�@pm.�˸J��J���מO[c_0/�;$0,_$�ޱKlç�h�\w�Oa�h����T�\��~��tq�=���)��'�I��īn6�
@����3O��nc���l
�5(k�x#S_ҖwrJ$�_���gQlى��%���o�csv��^)�����d��柼Ѐ�E�Y�כW6��g��D�#�nЮ�i�\�db�w
]Q�e�̛+� V����K^g��Ui�}�b�nz� o����[Ķ�He��hܙ?J�p��3>�7��1n�w��"��tu��G�8�a��Iiِr����s� Jy:m'�R��P1�c��tG=�C3��� G�������1 ���5�;��_�����X��������L�Y�]�C��3�Z)7A5��IOY�̤9��������#����4�*Y)�>$҉?mSDϢ}��W-����:,�+�Ԕ��P���ӎ�:6a=�	ϹI����m��|c�]�tD�ɍR��U'�V���	�H��lF};!mKc;�Xe~L��@��]��[w� �g}0�V~iA�@]6�Yֺ�WE�G�E�NKy�N|��'����c"	IjMpQhJ^���I��M������*��E�9a�!졏}��lN�~s#K.��7ſl�8D�����2� k�Et?G�&��((�n�w����C}��Y�9�u��O��PD�D�N���Ehih�*:�V%]��	���βa�+=�"m��d�k<z\�q����Z�^FN*J;B���7�1j��0�gr+��ȴ���n����@�щ;7_� �'�E�>�?E�����,ܢ �NO�������q��?޵�?#�7	Wak��R� Ɏ/ \��򗽽B��p\��DgS���Z�)�ǽ+q6]7���,^�Y�[�z��+�11�.�ʿ�!�Aaˠ����׹Aw��R7�%pSʇy,5ha�<~G�jm�_4:o$.i0%�@#᮹t[��r�P���^ �vM���u�	Ē�8j�l$47X�|���1z�� �Eg�s����"�tbv�E�ˆb8QϬ��њ��]��*��3`�}"�檆C{M���hѠW-�+���'�����]��h�,�)�dA}og𬢁�&��5߶�T�Ȼ�"��r����}$k�S�w����J�6g/�at4t��]<1"piuY�T-�դ�T�*�KZ�N7��*v<��.RWBx'�ȸ:K.x�Bb*
jn�);���WHأ{��K�`�hɆU��H�[��e'S�E&�P�9�Kc���k�p��Sѽ�Vv>3��د���%=����i%�� p�EM>��E+���͌��K�AQtX����v��D}C�����e�E�(G����"����D|al�7�N��+~�J��w�n��m"���D\|��su�t��D�F�]��_$n�\�/��4��;�?�Ѭr0�OJ���H���b��>j���8��G4��-�M�n�	`}�m�d �P�����t>�#	o(��U�c��J:�KO�� �V3�U+��U�o�ǯ�[�m2ߵ��Y�*���b��\+�U9����x�CL�q���?r��NcV�t�ŏ�{y��wkG@:3����A�HGx�Tڇ)�,��CA��`����#ı��$w��@Մ��� �s�{��9/N�����Y���~�l�{<`?�a3���3w葫*_H�Th�-��"M�S�G�n���Y����Rc����\��7e#�+ʏgL�w�4�.&��7b۷��P����9MN��GY�u�N�,��F>ߕ�>BA�Mt5{�7�o6��r8�/�o1e���Ir�I����'J��C"`��f2l�@������9�.�z�߬9R�����z��+�l�� �kI�S��Ֆr�Gj�? ~�z4S��կw��Ϝ��n=^��K���\$�z4�jf�	��@�c�bG���`7���ԄEe�RO��6��Bw?E���#�,�)6B�{�x��B��`R�H�݋�\'��y���O^���#8���"��NȘ/��;X��.f������l�9��^��sfro��};����Ч�}�4 ���MW>D���z'��2��}���/�L�z#�� �Z3�B_n����A�V,�G�Ο.�
�~�nr�P��'' �(Q��hE��u�,`��R7g���ff&'G�=Ε�����`����[���&��������$,�y��A0~�$�	�'�b�v%�} ��B;��.e+q��������K�+R^��J�W�
���e$S�R���Sm(���D�cw02��%�2���^z�{��7U��Я!U�} Qs��x�~egr"o�f��Fރ���D{	��������m|w�[O����Rw6kb�w�Mȳ7o)n#��*��g޵�;�gz�Me��ߞ%�ҿ�㱱_D��i=�� �{gI*ISQ_6�Q������$�4#Mw��U���Wy�J�����"�["�o����*��ݭ���$����CUH�1�ϦG!�Q�h����8;�h�h�=�cy�M]�K	����iq���ƌba�ז�	�!]��y��h�PLWm����M�oA͍
�u����v��tHd�-z:QԌmyW��R�A�lmX���"��U0�w� J�Xф��?=R+*\ň�v	ab���@�<mOʊ��:�"9u;�X��Nim[�"<r�:rɍ���xp٬��i�0�KB�4�(���.����^����@��8��@e�0����9�uM�4Q-(���Z"d�{0v�e#�b�;��$�n����/�gU���mJw�cV�"���a�!��'e�̱o��72�h��>}7?a&C�A^}�W�?co��P�����QdP	+ݠ������+&��sW`�]��=AA3�:��L6�3i�@��×ǛF��ZBᨮW� W~0_H����qἍB˩x�7�`�~�Kf��~_TwQ݊R�Ð�'[��X���G���H�-��t���ҭ�Q�����2���p8�z�C�x���ڹ����?�>.+�>U��k���}�x[���&�K��U�$�aϳ/�6�'b
�x��$C���K[�n���ɢ&�3R^���
8w9_���{X��Vd�W�ZԦb�s ���X�z�h��"�o�8~�����#j�)�\*뷗����q���OR~� �X�5�.�m���t�!��rM13B���|�	�(S�HHcC���w� ��#��]d/:�g��D ��$�M�A3j��'���X9�L_WU����W����lkǍt��z|&+[�#["퐰���9ٶ��dez�\iQ8��u��=g�fm�����GO�����@p:����jɷ��}�ڴ�� ���[���5�8��Ŷu�>�b1qll��r���D��s0Ț�E���u�-����z�VHM\}$0[��N�  �|1����*a.h*3�;��a�Ў�-��G��0xw����Q��������jv^���1�����f���~	�����7V�f���ܫ�H���KL�F�˯���4�a皱���.h�(ۈ�ҩٱ-��=x��AP,������n�VD���1#˘?4__z%�<�O
��|v��1P5�j� �TA%��ڣJ�s��3��`\ݐ]���\����YfG�5H�km��D~(�{$��(\M`Z��
m�~;��]���D�ڪtL�Φe�U��U�#��_�|�!Ͼ{����kk�����=��9fA@:Z)�7��f۩k�t�*Js�6���U���/��h
֯��]U�&�)X���ݏ���U����&ܐ<����l�
�?�~H.Z=�K�LbĿV6j�P����R�? /~<�VA,gt��П�86	�?���>о)���֕��O;k�oȮ�s�����B%�(-U���r<�"7$��5�Kd���~�Z���7zB���{�!��!i�:��і��o��8w���H�H�R(��>+�D��6��Z
�K�}n�{�϶��7;RF:�QƄŢ<�k��A/��6u���$��˯'.��6���`�SP�)��0?e���G-�4�-�<���[8'rZ�&y�乿qC�A�';ηx������]��R ��>����غ{_{����Vr	N��T��J^�#w�]���Y��bQF�^��:N| 9ã*�Y#e�ϡ�_P��R����'�{��N m���=t���^G4IKW]I����o�o�ʦ1\ڤ�6��G��2h6m���?��XhY=ѤYO�0/��#R���ܹ)0�H`IN��<�$}�qfo��sH���䶡����PShw����?m�ʣ1h-�A��#���Xr���<�]
���G�ԓ7��l  �ϠY%<#�`�*�'���ջ��s�L1�Zwy�	`;�Ͷ�ay&&%CC�-x�>�D=��,��1�C��EO�=ڹ3R���A�:��% �A'nIU�ì����ȚCa��s�d��k�Ɋb�'�(nT���ӣ�'x����B܀[G�z�⯁����^�o�&4���H5�2Ï��"�9b\��;�*O�PA�����j)i���~f Д��a�i�+�RuMY��4G#U
8���@��LCD�v����g�����`�9�eD�����@x�nđ��8��EZ#����C���H*!H�G��|YƺWY�`�+qI��_��5ޗ�ψaAi9Q��y���.���^�m~q@
�$�2��Y;��U��f�G�Һ��P3���݆�����*Dx�d(~EL՞1��5��_�*}�l�Av�5j�Ju0�ld����R"�B�\ښF7>.{bd���1
x�D�ΓӺ�{2)lI�::c��p�#��p�Ւ���+�`8�A�`�rI'��m忭=fǏ!��`u�H4ҷ��RCuX��֢F�� �A�=]�e[�e���b�z2#+e� d5F*q��bt���l5�� ����e]��AmvC��i.:�?��6��%F�\nx��˶8��
�n�78�� h���Lƫ�"B?P��I�x(�?GX<
���Q�Yy��;�'؉9i�F��lǭ�ٻ<zc<|s�!�5.	����m
��c:�8����k��75���HԈ����)�f�	WAD*�e0S�F��{JP�-��!Q����f{�h���=�t2_��C��b	C$���h�b[>zK����V+J�[Ʌ�z�@������H��)�Q?`����%��a�PSo��Ү�x�ޏ�������C�3!�P�jnXI�>;tQ�JLq���/���Le��G���2��\�.��Pm��V
�!_��_�R-�4�t�أzm�}����͛�T�k�����#$�x(���f�m�����z!������̙��cK�L�5A@ #������{uJ3�c��.V�R���I<��t̓�U^�Ý�-��i�Me�F���2�sm�,:C�{��������	C�J��씆����I���NƦ�������*�����c���U���7i��^(4I�t���z/��j�+�ʼv�ܩ��~�l�6��(j���O��|s���y��{_���Q��J �Er#�2O,�)v=�I�)��W9 Č8��')�@��9�:LE|��[6�7�Q�;���g�q%��y�<x�M�=�-��G+��Ġo�qkB��ם��g��= �`�^�)�I��ۧ��G�u-"o	d��������Jju`��p��y����]��ƽ�B^V �����q�L�nA੿���Ѵ��1
��.S����x
�B��Tf#*&�
�Jo;�VD�)��j�˶0�7K��T/�K��D�k!�5�5��NN��d�qzf˃BH��@�@��I^՘�(۪����A ��D��A3Ë� m�ˈ����[;�]_�sc7���kDf�d��w)��	$��a�ٔ��!��;��Ģ
�MȽZh�g���'�V�#�H�£>}Y�R0�)� �_�s ��T�*�VJ0#�ݳj�ߊ�_�Sd���� R��K�;W�c�U�$Eߍ�<I�x�Ë�L�^}{pF@���`i�T����ϜvL`Mt�=+8�)��}�B^D},�ɱ��Q��u���)��c�r��˰<2��GX@1�b�'����|Y�.�L4k�V�b;�·�6ߧH½�_N#�i��(͏�Z��۟HQ�x:R�F���%��#ěKrX?��1���L���֭c�U9��Z8���Qo����Km�+�˫A2o�4]���H���@G�T�¸����4O�P�,��ܣ��Ou�9������1'W�����\.��I8�RE��k�So�S�W��L�3�0wժ�,��XVY��QZt?���"���0|�B���R�wil��l �s����V�`58�������3��ǖ寯X"�D�e�T�m:�_���#<KÜT��S��n��Mߞ!! �I�?ceD"b���5�s����FR6�^aCŚ1ˇ;�d�1_�wj��|�)���2Еʚ+Y��ZC�&�?���E��>mqg�t+W����:�|�Fm�*<�ն��·V��Ĭ���i���N-QN��>�!(qKoM~��T��4�|�T������(�f��A`Q�񙖬�vV]X+���;'يk���qۆ˷�5��x{�� ��̹`ҪJ�	y�]��c�A�
��6"�v�o�)Ԧn��A	'�BX�v^VEF��@�O��Ď��O0ՙ5��x3��bf���1N��C����Y�"�k��W H\�o���\��r�=�PA����1���C�=���o�=����6
��x^b0�@E��5��c仟j���:�l9\2�>�̆��s�V�q�=��%W�'��5�5!�3�N}���� ��IV���B�s��L�����8}���R^�6�A�����i�/�B�9���Ò8���N���J�P.[Y�ʱ�xY��2�.�zX��Qݔd,mk�e�D�z�z������C��GY��qxy�V�nJ�ѧ\�[)��� R+�A&k��*j���^Kّ%vU�a!��u��j�}��'>/t�|u� }�_B׈g���Jȉ�k���pA�7"-�$	�s���c�h<yjYAm�V�i�r$�j<������O��C'e/��Gʚ���w�<���碪�x��k��a�c9�$e���%��=��M5�H}&@���vŝrO�m}���ww�0�lB��#L#������Q�_�B�ܗ���p��2.~�=�.�k6�%p��T�� �����A�)�:�`%��9�V�L�!�LE]�G�K��O	��zJ�����Of>� �6�M�l��_�69ؑ��>�!��JCԁS���_�AW��%��8���Z��$H&�+k��%���͆O��J�<fq�ӂHL5��W�����>|y\��+fE�ox�}�����O��f�RGn�����d�>�'i���>B��½_'���?��J3;��Fb���Jl����f�5�F�&�� �z:�Q��[��92�s8�$�n����SCrpoBm��}%��A�Y���E1;k.����ݺ����N�k��9�ƹ��t=VB��2kJ��K�N	�([�0j��T�ZUR�D~,C����Mw!w�*����CMꍐ���|�31��}�;�g�+'r�{궶�n��<	��R��{O�a2�Hm�igs��[��䶚�����d̫����u�3HX���]\��N�A<u���$I�7Ӟ��h�}x��.�&�c�T+�?X��#N2�C�-�5��1�"(�#��r��j '1c��:|��s����+��؁�u��M�vN����_D@P� C�5��o�m>�'Of�M����_��	p/"���K8jD*��2z�}�I�dvS9~�PR���䢎*����3m���W: n�!w��!c�ONmG[��X�����G#�`�XO;є#{�p�����4�!�o�N���mP� ڵ�5	=�WuV3�Yxv#��g� )�[�{lI�Rz��U��ǘ��cW�W{�ز�y	�o�xP�X95�z� A��űV匞��N�ZdvK�,����U��f�e?n�V�}�I'�/	����Q��b� w<W�,��n�ʽ2������U����y:�Ӫ@z��?�ǧx��ܓ�15��t��Ĺ���OP��;�"�
����p��A��{��Cy����&�o����}=���9uʻ#G�c����SEs��ͅoW]#�g6S}�G>7�`�c��s|�^󖻄!���H��Rt��G�81���ՑcJYq��p��_��+����f���с�;�ޣ�L�O������-L�r{�%��v�����3v�<��9����<d�*�7N�������?��ZqL�ҟ.�7�\�Y0ـ�}f[�J���=�.�L�;;�1jђ������_vEf%�%���[.��y�+��1/>C�Qy�R��m_���Vq�%'����U�"\��?�c��hyʞ�0Yt?Ρ
�����$�0����Tw�Z��rs�^����� n���<�4��s���5Ӑ�瀡	��h�����Hة>ɞ6k  �N���ym����H�{���#F�;]J�`���b�S
��Y���:���'h3��'�Ybمw\���>"䘌Q�5��y�s��;������*M��he�ԝ��jo~eo0g�컵�=��i�H����pK�A;)�;�IH�c.}�u�h�>��G�A�p0'�˓|CMav2YG��=l����G~��
�Yߌڶ��:Ԧ�
R�f�zL��ؘF�4�\����24%�Y��0˭��6��l�yQvHH��
$�ۼ�p���:������f�#�,�M����,!�����H��	�>G-9�����.�a9<���mg������t�n�Õ`���$�����G��nE��u�T��Bš�c��`&�X�J��@�����������;U��j�ܿ���4�CZ�0���ϙ��&���l$����Wu���/OYc�b�Qu�2ax-�N�Z�j���a}Ҡx���ϞL��*@A��[,쁖��pA��M
�;"ʯ�(�<qW����Ӊ�h�WyRf�n����<���[zR)�����>q��`9�����x����N~�w+ P!��.�O�~-Z������Zz�\C3ެHl�_YGO�w!�"�����Eĵ��G�p�^�Aه/[<�-�Ӕ�/u���xI�k�G@΋΂�ș�R�	 ?}�
657B;��#��{����Z�g(�ss5J����͍��;�},9yCX���YJ�4�A��[�w$����ߧ��[O<ue��n�,���L�2T�*ӡ@�$n
�-,��؈V�
�[����\F:kt�2	u~Z�(Ҍ�1y�4J�~jM���V�vN��,ź��{��_�1u�� s�':��>�h|\��@�ӌ�xJ0�McN����6f����ƛ���WP��[�#t0��Q9�`�z_��L��կ^�DkԳΰ�9�\���K��S�Y�Bi�mp�ӹ+�?�.<۷xj���L������č�;����x���ЋG
���Ÿ�F��r����n��Q%��,�+��31c���%+�t����7
�z ����5�Ŧqƨ*��l�诫��k4�&K(J���m96q����T�ݭR�Pk=O߹�H]J6v� �/�̑r?tu7nM&�{|�Z��6���n	��J\Ү��c\�S�nf[(!�c3�l%�3Dcۜi�o淐�����A}s��r�90���(%+h�i�e�Mu�an�ȇ��;��Ib��zL�+\���A�8�IyC+��=�
�oK�X�xa�\���>�׍ӛ��@=r�;A�O��ͤG���0�O��~�O�5�k�x�Ő�Aۺ�p���6v%ASC��t�s3~�A-p���H�C4��5��P���R��jh=����:N����/G�$���K�&F�'zS l�y��Ԟ�$��۲��ӱz��\�N<~��1FPq���݂����"���;��s�x�9a��c��Tè7��G��}ݸ�?��3@�}�����~���ZeI���]�ҚM�Sr��J�g�'#6�z�5%/�f-�r�1������j�Q���p�}�o����C�}����Թ����L��k�8#��8��Y]���|JXha6�<v��?!$�&6�%O��A��I%������ӥ�旀�\�S�4��P�>���c��M*��C
Tʍ`�q��̀/��~�{��/��{��9S/soHr<R��ifz�)I��I.u�;�*���m32��Zl\���Mm�Y��K/�;�>�^#�	d+y)��6��6@��5-�QL5`�_t�S�T��Q��L4Q�sB��m�YV�+v^عCMU�j���z���תJ�޽��MX�/�#y��7+�( gջ�+�0# ���7����d9ZX��~�"�����kv	�;0�ܯ�6#�꟟���ݭpƓ�nÚn���K)o<���a�.׾q��G���
cg�$K�A����c��h)�:��W��S�+����WM��k/��N�lP��'B`,�!�w�(�
YE^|Q:��T�O�ȬF�O�0��y�.�qei�F��@��v�:n�3V�>��*u�~[�u�z�vkK��>�<~M�|���1���$ʩ�/.wIyE�����uvJg$��l�����'-�L
�rHT�'��q��.�����`|r92��M��}���n�o�O[QN�kx�n�*>��dŶ�(�I?���KZn$���o�\ղj��̭�r�|�ZnT����K�>.YV�y��R��@��7p[��;�{��#�&��]��i�? ����-���LsT��a�;����~�9@}Y���,hRq�E@�+>9ݨ��p?b��J �ö��Lf�6g������tk�z��=�u'�=)VU)�}�9�S7C�ZHr���x�tw��˖r֩�^�1�Ʊm��w�%�?< f�q\����f�E#���$k,����i��<��+- F���w��S���A\��ތ�)��ȳ�;;�����P�7�t�|�0�y	�āe������{�Bc�f(Z�ݕ�x.w����ͯ#l��l�<	��x��#�U�?�֖i`��WD��c��;_:�I�w��r#��?��,��k��:���:�ϪU��)�6�a�)�buo%c��(�kd����@��# ��b�oȎqg4 1���5�J�	�dHNő��+�I�v�[�8�g��,:��&BY~O�a 8B��m�n]/+"�cZ�wG�f�&r̕��x�XXЉ.�����(� �R�Z^��]�O����zބ[z�7�R
p3�V�k<cA݈�	q��R��*7���6�ݺ��$}��)��eiT�;S�[F�-�T�V.�� ^E��>lm��T�O���;$��gm� ��\����Q��?���
3�9s[7�[@ZhH��"~�nŵ�9m]��7%(����Z�-�P%_�!@E-S�u_i�\�����2*P����)L~ }(����i觼����'�؊p��H�*��%|]�'�r_q@��GQ�Ϊ�6�9���b�����+)���7�����XK_}�h��<��m��!���e;���u9ATQp��!����`7ii���y�yv�l���E�tβƇ<���ab{����~� n�Σx�F�� Ea��_+a�Ik�,�a8�k�_7��'']0�$d;���@5��;b�'x��������K���y[o��S�iR4�M�M�����]V8��fwy�S�wN(A�~M3}��ǟ��yF�NM�Pw����f�� �ܛ�׽\�P�))S��ɰWTѲH������J���lc~�7f�o�Jܴ,T@Fp���D�DUJib#�˵�U���0��ݻ���1u9AB�Yќ�)U�;��y6ҝ��(u�-	�l��Ly��ґ=� qQ�z
�]jynz�8�̀,��ڽ?����1��͖6#Ÿ�(3���Ѹn!�/z�u�_��3��A�{6N���n����������fY��\ꪼ�36�@o�p4����ƃ�vg�O=�a+�1��}|�Wy���k��|���;�g�@�C�6�L��wDU��=�&�r��G�@�Y�,|�>Aɕu�_Byݺ�n!k�{p]l�ߟ��nvWtHS%�HO|��5���>,�y.�U�3��9����'������ϡ"���YG�^L\5� f'Ed�����������Kf�Η��Sq�6�
��J��M�W�Ņ��W�Yi���S_���h.h���3 ��>�)@��3�Bs0UHoT.gY�O�I�0">^qK"W�$7�>�?���EF�r�&]��E��!����%�(4p�7PƫҺWq��d��Q�p�<�$+�@�0�ik�ݶ(B�S����gZ��/@�H����^ʹBW���X�G�}}&}�#�G������OhQ��ֹWG/Q�*��sM���,J��>˷A?ݵ�ɚ�l6�5���[�!Ǟ�W�� X�j�J���M�gs# ?�`DQ�l���;�����cM�M%�K[�l�*��`�}2�o���F�*M������AK�)���?WB��Kz��md�4HȊ���l�j�{�0VMVג�C����/P��$�X��pg`���QY�+��}�^~��;��vg�m�Ĳsa^�@� �1�s �u����&�bU�����c8�-T��^��?�m#�]��Av�@g߲#��v��=)���u�V�%����PT��+�h���Y���`��X~��jdO�I�&)��$4�Lk��:�-���/�:����܈�3�^$iY�&�:�u���'Ў��a ��ۅqz&�n�H����/�ɐ�	����H5�tM�Nip����z-���D>˥���>��5���og¢z+IL$Z���:8�����[s�89�{�/=�����I4M
�|్��_����Ay�ĭm�Lo�b}�������l���6�	��<�tK���̓U �f�n�عx'�s�=<4$[��"��Vc ���T���Z�h��{tǔ׷����!ϭ��l3���K��O0�!��_��Db{���?j"aMg���a��}!�e�c\ʎwd��o���H��zp�cQ�sz�,o������'cew����nO��#�p��$N[)�'7�C=++&w����5���9
B�b6J�e�� ~���	ha'��T�cMl���?�t"��r��\�P}ln� =x����,��W��u���/v+��J^$�/Q�eƑ��2/Ca�Y� �Qw����_�ԑ�e4
�m�J��iZ�z�C�گ�i�I]�����><c5�'I��:r:<${��\Ou@���ņ��.�B̾�&:�#����^nLN`���/�����;�q_�$������q�A�{�O#!Nm��
��T�)�i���u�M�7t�n���s˰�&���7i�!�}MD���j�!��lMPY=A��f�~!Ё�q��cjpa{�U��2�E8��ô�6�;"����}$����W�������~�!0=W9�O[-L�ߓ�MJ:~���/e{m�B�[k!�|
�5V��#dmW&�Ϧ��J�����D�r����Hy��M���(;m����l�uk��X��rڅ�֠����jV!����$�Xr�#�#��\�K�5E����w�]�[��q.B����FƋ�u����yyS?��
Y��ȁ�8J�aI0�hB�A�i�FTD.�HLY&�3�����?�C����!;�Qs^�Zk_.����j�	;������u� 0+��p$���V�\����P��̱��3q��;�/v���t�v�<�pK�0D4���jD`�U��U"�79��W�,1��s��'�ks';c6��3��ˤ��/�;_�^� ��-�}�ux�{N^�2G�'ϊ�$.=ߙ�B+�]Oq޶bb"�{G��|�ȑ�sNtK��cG6-;�����Y�VZm1��r��Q�����R�1�D�/���x�뵑��DchQ�3��GҌ���5р��f�����T/gD_O�1�.4��>�yˊAO�R����2�F<w��Y���̴�C?� ��2d\t��L���A�҆dni7҇�QP��"�  ����_��ymOɀ�F�Q�R���
�|S+�u˯��o���NM{Q6�"1�#$� oH0+��/�B�����u�]����z��O-��G	A�,�� XF�>�[�v�-��@|���	�.����ZJ@�3��Eg`�Q�����6�'��f�ᐎŤz��a-&������lc��B�}�ļ$�I�ۧdj<��1�6�m��s)O�X��T�r� ���ؑ�Q�����0l$M���s��1���24�G����N�sS�;�XQ�|X�.�I������9�z˿m�����?4l���d"��xD2�P�O_��Wk.(]���ƞP��o���$���|)�Oi����6���6�錑�s�,G|����q�ݐ#�4%b��,5X�@�po�V8v�e.$��C(>;�S���&K�#�փ-R��5�b��ї:n.�A* ���d7[X��`	�����'�ݸ��¿H̴-�X�z������%%ߕ��@�YR#��ik�ר%W"ח/|6�st}��s��E��W�7po�E[�f	'�p�ɮ�O3ԩ��<�0��W��/�0Z���!�m���0�����[X��������� �� ��4ݾ���o�ԳD���v�1���|�7�i�07����_�ٸ�|�6Zq�F�(ÖiV�<�=|J��k�����?2�6Fp$]��'����QNH/�gϲl�t��꾳۝=)�j�)x�ea6!���j����5A��t�V%f�R�Ʌ��[;�(2�{Ql��?�lޚ�S���a*[�Խhh����g�{�(�5Yʀ�½�(���W�"��-W"ʝ�	 ���R(�F�_@�{o�`��~�I��ԥ�<q_��7r^ߏVJ>�U����HO���Q�Ƕ�	'�7R)2�|uk��:񌛥G�u�0��	�Y�)w�DI
��J�O\�O�z[5uts|��P�P�Ʊ4[.ٓ��ㅎ�DFBt�'�}���VR�F�-��l�O{�anQ�\F��+� �/7�-P>���uo�ƞW2�+IմiJ�!�Ʋ�"~s��V!��T���+�݋?�.<�O��Z�ZU�����7P�c�	+T��ȭ���Ѽ�D�v�<D�_F\���^�����l8�	�)A�sg�}�Q��֒usnfx��=���f?uOa;/���[o�$_��|����hبވ�g�2�����F)e8�y�}!�c�ݟm%�S߄8D1@B�2��,�+��0u�N$#4D{#��)�}��:�3��P�gE�U��àj��Y&!�3�8g�,�c�j��6��?���G/>���`>I�-�U#� �·E��y)U�>H��m&�悒�(m
$���*�T��g�PA�P�@�{�|���?��oqb�/�t"B�R��@��wΓ$�zb�+m�a	&Z�B�f��G{�XP�P��p꧝I��ܶ#���,@z��Dq��!���-7WO�M�@]��ܱr�ط]�ď!}�L� �C*c�Ωl7�U��J���A���AB��0H��������OɊ�:%����1������O�����
B].<7�l�ƺ��J�i�R�HÔm2���yVF�J7q�Up)�9=�=��/ʿ���|eίE�M�7��?��'�uz��3� u'3si�C�s�(	�<~Q�0O�e�I���8�q%��z�ݹ�v�P��M�ĝ��ƙ�Z��0��Z��7�~�̸�&z �g��v�眘�{�|�Y�D�&7-�ub�c�Ha]�����3g���6�ϣ���q����2d�6�}-C3묘��}8ǻ���f��A�b7�c�%��)%dD~��/ �F8�BgZ^Ҽl�G�"3��T��nf%Ї���󸮀2����ݨM�O}���j� Np^ A�D�:֍�B��z���3��F�x�O����.у�eY,��|*�������qI$P\fʃ�H �g͡6�|�L�R�^�� ��%	��"��S<�Btu�(��	$bT�)�������"q-��]1������A�&��*4���Uډ�>R�${j���i�H��c�����q��7���
ኤ������w���%bB��V�1c�$Z�M�2��ZgD��I�uީ�	?�M�86r��i;?�3E�D�84�\��G���9��6A7�[��ŏO�́,��L�.J9#�Kp[����������0A�8��4���sï3�e��l�ܪ����Q�z�ό
�u������NGzY�[!�P(����{�.��j:
*��҃⓼�91����~&��23F��M�B2Տw�l�H���Z=�<*�LVу&�G�i*����~�:f}�B�<v\���e�����k�ߒc�:�O�)\��E���a��%����am�\S!�7pWn��2��[���}���84�f��.	���ѶR� �8S~/��	"��'�Qw��H�7a})^�z�.!Ӫ�.�J:�&������Z�C-:?0g�^����{�gj;
��M�4���5�Az�p;(�RI6�k�������&9�3Yw)��S3�ݏ��3=}8P��z�:i��
��:x.b�a٤�F��דww����ڄj����~���<?lt���[�Mm	�{ǼO�.��������������Дz<��?�1��H��9o�-B�qlLD�O�����w�鵍��=kb�d��7޿�,�����D2�	)gʸ��1Ӣ�~ht�� �C�Y�u	��R��C���zq"O��H::�d�^0x���y�q�HF%���F'ӯx��TO�0e �D��Y_rMl�O��@�Jl�yfp&��ڰ6�_�/p�R�%�:���W+��Qcn��Bp_8��K�I�A��]�Yٓ�
��$ӒP}W�I�䤒jl�!2����������X0=Af���a|�:χM�M��eʡwS������Y��8r�$�h=��B��J!�dS+dM.۵��?����'���g}>u��t1:|D��	�A��l�-�R�t1�^:K����\�.�b��z5�D�p��5��]�ݱQ��};����9���͑�����d
���j5��۽=c�̯']�J�K�hz�`��ec�$S3�?�΢������h�Q���mkAs((��v�K���4%�P*_�� � h������r�ص�y���ǨtQ�O0����$&9"x�⎳����
��'�y�w��I�X�ō'đ*�.�G$�܌
XL/���S�y��N6���a����'�ˍ_��%�
u)�k��_8},iy���l�P���E]���X��n�"�;���ݨ�ݑ�ã��[,2�Zw�Gt�#���5v�<�\�&՞�8w�B���1�YP�'��:�\�qw��Q� ���;)]�V�7������V%�"3�
�L�N�}��F@�S|�	����.���୐<����p���=2��e��б�@¨�vV��I�nl{�uSޟpAD�M�����#o�Z_Mצ��O������ѱC��He�cɛ`�N�WK�
}����:{�=����/��08�{�J��h�!��P�ҝ��i�It���l�z����e.�� c4+g�kq/��`X�z��'"R^] ��c���Y��uB�����X�-5���CYH���-��
��v���}o�����壙v8�b�_�u�>/��jcv�Zݥ�#��z�(���q����@�#��۴fy��^"��m|24�L���S��h6˗E�Co�u!�kI��	��u��]�6��5�k��L�㷤P�@m�=��FN�0]V�Nn���l���M�q��.��CǺ��H�Oy�����!�F+7�-�Y�{�֥�}6��]�p���J3�6���Ж\���;�� k�tA9���-
�#�����7�'�>��SC
�I��gMvP>�c/��i	��S�@�~%���}���H� �c��>p������O�G8�	���+�q
F�+Z���vl�JG�4"H@�z��틯T0Zkb���P�I!�Y� 2'�����f�
��OH,GA�����N���!te+S�e ϙ�u��P��@\+�^�l�\m�����婸j�XR:-.-�t7|��g �
�w`&{�@���/��	�c����Q~r�������X��qB;��X>X|".�L�#��'5ؿj�fV���QĻ<�:�����w�_c�B��4�W@s�s���������*�x�o֛m�#��;F�r`30���mNNkĎ�3l���˨UĚ�c�#)wC"���ǽE��D�8�U��plϔQq˥:�4�:��.^�1��=oM�����	dx��M�;G��x����¥/��eR�eJ�='�1 ��0O�`�x�6/&:[��"���do��ю��6,��2�S,���s%6#t�,Z�G΍	v����fA�9U�A�X)%�henj��8�9�����(.�N"��R�H�_}��<�_�2�z\��*S���C�U�9�V�-N�T��-�l���N~�U����dӘ1�j;Q�{��/��j��T»M��WE�҃0�g�k������]�3�Wb��$xa�B��#ě95_�2��ޯ��q���ۯJl%�>�1-�q�3�\	����h���3�u���ܟ��V���Ɖ(�oY$2)`o
����^�4�u-3f4�y�q�2��s.��WL�}1!
;ck������A��c�oZ��.�yb�ŷ!����0@�9�δ�������RՄ�	�����V�I�qե�Cs0S���w��&/���30�s�s_߷/�=��>���W��h;�ϫ]�)�@�AR�(���</�&Qu�d��',��B����־^-�rh�,���>]ls����2�K�F�S��SP(<ɩ��|�}ې�J�M����,l�T2��D�E���pik���f.��EQ�}�� ��v���	��g����C��u�/�(Y$�����i\������vD\��.��Δ�R��_|7�Tj�À�Ed�Giq�x��o�)8�E�a��@
���f��J;�Υ��6G���1��r�1���|���]�f�x�M�/-`Aj4���5 ncy���Kɢ�2Pv��	���`��X�۶������J��p.ɴ�U$D'�A�@�ג���c)������$��4�	\�s��|EX8�I0E~�]��W�� /}���~��i�����ק�ϣ����x�������W�/(ݡ���4��M��a�����7aƨ����e޳�rL���<qp�z{�"GX��4�F�Y�����cP�q
� ���7U���	��Q�5M����I٠��;�L��R�iY7��kļ ��8�j�y�'i/}g��.GNt�2�Z
E
���OpfTl�H���S�;I�\,b�/N�="��ʷq�$~�J��z ���v2]ԩLD�r�c�d$g���+A=���$����9~�'�`�q�ѭ���A��]+�tI��t�0w�7k�;�dC}���x��u��O�Bx����q���*�]Y������LVUeq�r���	:���q��y=�o2�k�6�Z�=qy��I�rN������pO��kLf̧c���`����!�`� u���C$��U�����rŕ�_��څ��Z�LK�A����K"��v�99 u/��*|>]hN ���E��91L�\0�}�$�2g8X� �A|�I+�^���O�*���!�W���W�=��*��)�\D��{S[�t$*��=���-��.�P4��ٿ�����
��=�ҩԜ@d�"Aו�Xw�
��h+��|.cK�@��-�6��'!=��s6fZ�B/�̕@mTw~������s�Ov����:�%���	j��e1��-b�ڂ��j������݉��ތ���Ш���r⭣��U����CG�����#@�����a�x�[�S4w+�(i̓��f-#)�~���ה7�Ƽ�]���x��U_Wh�i�/��a�>(�3n>QjAW�8������O�7,n��x�����m��5$^��*/+��T�)pOE��\�kbp�@t�Vߊ�8�z�Ha;��6粬x�NeeXN(&��)sg�;�j����e��-��/C�~���.87�Xp���Hy�����.���DJK�1b���=��@`�g��O<ɸv�(�ճJ+��h�q�b����k����q�Ա�2vS�w�y�I�|��g}q� �OG�С���Y!��o��M�&s�.icz���g����L��U�Pͯ���\�	/��)��y���D��2���}��x�g�r��j��]�X�9��m&��M뢞˰�yn�`A1.)9lm�)}�W�3�A���'�-�"Z�e��6N(���R���G��n3>�G�Uq��jK�qibV�o�.@�Č����dѵЏS`n�ir$��~����ܞ"�Y��h�q2�Cy�%��%:A�1x�(���077E���M��l[~�#����3TR0*Ai`�H�C7�i|4磼g���R��(ӟ�Vnd˅��I�ș�\��l�;�48|ܽiվ/�}ԁ+�燦�殜te42;�SI�"�)?��h^�!�o���	胉�H ��>g�?X�D��j�ֽWіB�:��H]�����Vy� ��t�ݟ��v��+��凃�����P�#_�َ[���r�����\��f�*;��DG⭇�1�J*���
o�l)=�ӝ���mG����6G�e4t���踙��0w��"Emv�r6�K͆�P&濞eB�|"3L\?��UP*;@| ���@c�h��T`���4������1�,�~Eq�B��a�Í>4>3�����V9Ůr�8b�Q�:wfͳ�f�\�ʇ� ���'RM��E���M(}�3�_p��-��=��ڱ~����|$���S�|�ArN^� E�K��f%�;�s{-)��a�����a��a+̹��]��U�~6H�R��F~(W���8^8u9(�6ۖ�0!]�#=��Y�2ȅڎM���&S8�5;&<!(۬�I\��]n�,}>�Z���[T�:7q~(OK��UNJ�\mv��<�/�w$,z���
<�w�*
���Omy�;����u��2���{ ۼ�P�nc��M�0�/T-�SQ��R���R� 7��af��v%-���wf�u��O2z��f��M�ݯ�#R�p�Y�%��i�5����ȗ[H��mŇ�K,�gs�}hv������x*:~�v�ӐZ#eo����w9C��x�M����I��1�Rk'���H���&���{2Q���r5A{�gT� y�tblm7�\�ɓfD�1����b�����IO E�G&����9"�D��$��sp%�{�ڋ����B����M�+Ga����g�6q\���G�1u��[#��`������`M��i0��g�\���sbA.���Q�zQ#���J�5�������2L��G��W���9�;�L�h�Ĉ�hơ�$�1>������K|��ʛ ��P��5�Th�h0��J�a�V%&�	i���Ծt;%n*��8U��Fﲌ.�޶bE�͉���;t����с�xO�J�O4������ӫ��n��y�4�L�� ������s�j��Bq����P �13l]z����w��O*��	��[&�\� �Yw��5��~ �N"=��#"l�ϣ��Jf����`��%�i���M�x��̰�-b���	��'���:��H
 YKM��~K�$�k��n.����[��k�n�0�_�a�ҫ�3�T��tUQk�4��(������3��P���{Bd�~l 9��̆H���ƔJ�uh�w����z6�U������~��	>��v��+�F]�9D����&�Y�#�Zq�۱}�B�{���ج�&�峪P���|���_�YF~J!*�%�7�����tÃvhѽu�1I�����ӄ�'J��"ac�G|�����!�9���lZ�J�(ن�6mѰ}��G4���DF�Ƃ���[��}��QW�"cL����
3��>}�"~N}��}�XO�ס�2ۮ|��d"�U�yd�N\��g"�_��|��[I�L@�*���{�d��Z�s�"QwkH���h�{w��� 9�d�J����Н������mj�k�nDG���I臹Ta��7� }r�����/�؂�x��_��c�z�)�U Yl��z�9�z��S�jU�+q`5�*��_�"%I>��Ys� +��$$��i�{���I��F��GR����n9&�Ր��+#����]��M�o���
��-���Vy��X>�_g�G�@c��E� ��h�h���o�����:�-@�ud�E3�=]��C汙}��޻乥����I�t��-B�u
���T`[OX4�s����O��f���Ԟ��R��O4�����)(�DT�b���%��gp[V�]-�Y���#�(�V�l]� B�<��M�����?�_jV�%ݖk%�˫�����&O�8��#���m�x��YJ�T\4���Hs�K�E]��<Ѣ)S�y5g=W' �qT���)��,]h�ً���m;0���K�XM�t�+�w�a����s�kOe	���ǰ�3����r�D�1��u��t�g�2k�ER���3ӝ\���A^4��5�Y�����E�&�`�����{���}��ڹI%��j�A���')�'8�P�U��ڹ���;?�+lѵ+���:�F '�~ߞ[�zRq\:R�Wk�b����T�R[�4�o�L����P�=&��Mm=&�~ߕ���7����	[�C��!�é��U��{8��}%]S;ӳaʸ���ą����>~�L8 ��9��D�D�<�e4����ґ��tWc�6��#��딁�6� �OdC���Z$*C�ƍ����� b�w�D@l�Nrㅁ��ֈ�W���_ƭ"�
d�0��i�����T����)�Ռ���$��YLB������%��o�΂�I��8��kV����%h��:Z5��!$��A�.�*�{�mȶ��2���Ӂ�)�b;&�I]ܫ"d�����[t��x�j�������p��=�e?��.�\k��vW5Q�ؓ-����k�{cB[�����R=�0&�@;��_U��Q���%V��	��U�z#tU�J��neA��a���M* e!�/�ߘ��A��ݟ�⯐(g4,�*�~g!�3�|iR��X�B��T)��N
��O<�G#`��̷�.�;K'I,�!���� �H�ݙZ�)پ�n���؝���\��̫�/'~H��oq����HO�ZU�KC��������-q �+8b͞L�=��1*'xtPAg��pF�0����g���.�	{z0A�rv�t���A������l�M�먮%�v �#8������S�Võ�k{n�R;�f����q'�^H��l���Aj`@{�4�Ϭ�.�ym�Q�7�o�$R���[M��	�|������P(l�޴���޸$�ڳ#]H �ƽ5�T�\��ڄm�5�7A��u��.'
���"`�;�.�&2\�Ĥ�Đ���qrs��G/BU��ak��6�3�.��%��;b{f�/� c�k��)�/�z1�Lq�����U�j���-
���O�K�4~�����{���^�}?��[?vA z4 ~��hu���G��wd�I荎Erf,56��9r���EM��W�Fc\"J듹��Rn�Uf��Zq��+,���g�n� kʴ�M�w?��������"O[�J������7L3����\xk|>����Y4\,9=���MG=�����m0=6��ٶ��-�S�X4"�K�
��bE���z[[��JH�?�Sގ_�M`U�/�
Kۗ+l�)�BڹU"-L�\���r��	����^��4m��__~����.OY��~W�I���x�K:�r�F���ڬs��;� ���;�N��Ie�m̿r���q�k������G�K�����W�S7c��&�-�I���r�!/;��zn�(���Ȕ���?3��LU<k�!�2lSZ�j3��Ps�Rv?������p�
I�6��L�T��w���0j��Ȑ�u�|Yh�F�kXj���>��l�D�m.Fy����AQ��O<qJj�^�U�9�:�~ܭ	���+������F��TC:�v_z�hJ�ѽ�W�Ҕ�
�V�o�������!L�D�CE8���A@�N���I���l�2~�9�X�v������S������R[!X� B��$�*yd�͉��u�Z�ܢ@a��S�Q��7uyt�ԍ����4��E�������o��.D�c~q@���2H�3��]�vn{F�U�o&"�H��k3Y�9V]�/��n����jI!m� �Q�O�KIe�̵:�Íe�V�:����?�)fCc{�<��n0����ڌ,2X����X(�ʭc� ��_�D}4��~8��ŁT��D{��5&�- � �S�|z:���(�Qe��]��(��(E�.��+I�E��+1��* ��Γ�8�a�:$��&&Om�C*���96u�+ևǵ��3����u�I����5��[�pF��#r����C�j�X���_�F_�U���S�O+H x�56t��x��o��4?0�6*������(�#ɿ;YW=�-�u|����]��e�C��|x��,���&O:}�w'�X�Rh�̋�#����e��r_L����<�����'��^5����~o��9���ڛ���)b���>�ʜ'�x����5�=3�.��cL��0Ac����숷�=-r�D��E/XCf��L�;�Y��V�!��Á����1�j{R�kB̭��P�y�Tılk��s�,�Gj�$����RL���ԩ��7����Р��q��m����s�\�J �WQ���'�)/y��C�Ǒժd���Ƅ|��V�f.����L۠����"炫=�F���I����o� ���J�N�N*NEX�]���Y�&j�,�?AC:Oۂ�p���b\���h�}x�>z��f��m`��J�r*��Y��vs�p��YP��'��/�p�e�R���X��J�Pt{0�~G���ֳb�H����t�%rCݶ%��	��J�&��B�=~ֿ�!����K��݀�����%�t_Ή�3T����G��e�|V  ��L��L6��!�8���*���^Ał��׸]�r)h�o9��Pd�6a#���{ڢ����P��A�w�-�#�]o��f����ͱ���8�\s=+흾GL�����YL��nw�UB���C37�w�F�9�=;@�O&'���N�l�h9)����Y�H��FS�5�\h��~QY�-B�h�/I���R�O'�4���`d�}����Ga�ui��*5EQ!X]E��Co<�d���:��a�H�0$,�+�L5x�� Ep���� �bIaǴF:�ǹ��j�/�8�ցk�*�������������__�"m@h�%�h<��@�6H��D��B<�"����kU�O)�����}�Gbv��X�!�)���y�S��%�W�P�.�u�|#J�?�� ������P#?�L����}2-9w�H�b�Elm�nl~O��!�9B��~.�T���^I�<��?0A�<	�W�DcͼЕ+)����"���@B0<J/�S�����1�]e�:�U�?�l���6��-�oxe��`/1��-�z`SK����qֲ�ݷ�A�0�ٺ�Eb�ޏ�`:b�(�"���K���Y��׵��`���[��H(�t��U�u 1��29�r������93�d�9>"�����~؍K����hV{f'ʍ*�˲4R��2]�S�|��?���e���/[s�tB��	�Ὸ^ʹ�n�Q�m ה}^q���w�m�a�T	����^A]���G�9:���gfʩ)��X���
����s�����(�Ϳ�|��0�|-�/#Q~E�"Y�������A��О�7�=�U�'M�Z<ܱqJ߿��,X��!�e���w$o.X ���B�i���䐈�~x���9�����~J(/�dJ�LLu�.�Ĉt��<���������7w`]�i�~�ѵH��)s'9�F��	Inp�����3}�����:A�� ��m�T����س���3Gt�M��' 逄iܣ�}��r5�U��K7p�LU����c`;k�9��~��w`?f��)���!'�t���IV�s	�y躗�)rɟ�P9�]�L����t�T�eR��I�6q7��ѓD����@֝0�LDe�N|�(�e�:G"_��iu5��%�����x���t3�q�<�}�<��`6��i6%�I����a��tG�7��,�*#ӯ+$n�XpAŔ�Vp4��sj�qsɘ�E\)��T7�H����*�g�Ӓ<���癔(�=NXs<�L��C��ⷬ͐��G�f"�)1�Eҫ�ka1bR�K:�����ڻħ Mk;�[�����5	�`R��]��U��"��P@�n��F���f�Π�U"*"}��J�`:���8/�j��8�wd΂�#���N"��>�R�E�+((�_��V� ��!�t�S�
�:��h~ZӳV��JC����;�g�J2ajs�\�ql����r2��UW��r7�n"�NQ=�*���i�w�X�y��s	X�5k*�����ʐ�jP�=�WĪ=&��}���Ñ���.�T�
vQmE(�MU�`�����~���p0��ֈDZ�l&��<��c��(|�4"��E��o��LԐk�jAuv%�v16��e�2��M��
2��q�T3��l�cB,(֏�T"��y��t&$���k�����b|/jb�e�����-��|�c[ɥ���.��k���g~_�y|�����t��rϦ��T�H����Vע_�0���{��4�e!��p��8�Z�J�V8��9�tio�d�O�wQ��Ď�в-���J��ZL#�k���&�"�ڪS4C��^���R�O+/�w�_5��%K��O�Yjw|jނ�wD�zR�	2[	����,a[���}�����5!k�=w��[�~�hجfn�~,����jMu�����8b(�L��I*�<i�tFp@M���K dyD�Y��brn�d��t\h�hM� �!A����ͦd_b3�1�!QV�	�{b�'ﻞ���%�s��I����Ò�,�e�k}��F�����ܩAe�B �x�~p����g�N]��׹�ˁz��:��G�s0F<��9R�y�Qv�lT�
9�v�fOz����Y*�q�� p�����V�Z���D��pݯ�'�8(�%ι���+��4H#'&�늕g�h']/f����Ϥ>-N���%V��~Ke��wf6�!حO�������6v���PBu��W�Eu�t9{i]8K���n����y���f�я�n�a�uBR h��]���h�5ܕ��Ό�%X1඗x��������� �-6��_��rʚ��qI��[b�4H�.K`�`D��9���.\ �j��n��g���$y{S߈iu�DӨF��\i��:����� �d���S����X�5ʛ��W�ϛL���+:��C��wR/c�A����]����ȩ5*���R�l���G��@T�E�]3�pN�13���;?�{��;��-���42�>JS�(h���1<o�|���w5��0e^gt���= 	�y�H������ǐ�8�-\f�U�O�Z`�������,��((b�K�d�*�%e�pW��k.�N�i��P�C0Y�M2?Tt�����U&����8���`�KA����hFj�o���p�O�)&&2t�|�2H-zH�Xy|��Ժ�Zu��?m��R�0�c����~hp�@�hP;�S���	��\/� K,���B&g�&�9��2�sw#�,f�ȃ�o3�ف����R<9"�U�wQ3�����V'�f{(E��}iO�&��|q�]��˻I����ǚgQ �c�	q>��7��a�P�
�;/:9���HNj��nM2��ΓU����ڤu�9�E��sV��M<Q�h}i$���g�9mĘ��#��ݸ�7i���5z�	���VM�7^y�2)���S��b؜��Z�Q0#����Y6O�5�&h�>���e�[p�`j�zS98��5��v��	�8u�l����+�]LB�j0=�Ɖ�}��8�=_�U`6��WsT����cCW�R�7��T�JH]���k����Cyw�.j���C�>��ӟa#ڝ�`t��U.y֚ �#��k)l��e|k����FuK�m&�(N'���c	T?nN^q�Zi�R�
P�>������qC	_y�*�-��̖fӮX�R���j+p���i�P7i�"���qz]�J�V�9HD�zͫ}2W��!�b��F,¨ٛ>�y�V^�'s�_k�^7�jt�K ���6�В��G��</�A�+�,o(��^c��x�*h�{�����֝�3�$�b��Ro�S�0�7���[HGe�&,!^-����bY��G ���䦄	���B�:�a$c�dRx�mѱ�TRX�w��f^6���b�Y������̥�?m:VL��?]ؙ2q%��>iPG�8��>�����=�U'ɿ����/8W���ݼ��st����*�S����-U��i�a5�_�Y�I�iS��|���h�୿�bC�p~l�䦚������^L�7b���	�2"�!z��·�6)�+�C�v�����_&��Q�G7�����gv(]!����l�����p�R��=�,��a���2J!���}xyJ�9���u�1��3����c�D�#r��G(�RiX��߈OХ�L\�w�Ӗ�n��d]r�_�x����«����+�V��P@(�s�Qx�(\A ��nR����K�g��x��� ����H�	��V��.�`��2��z���s�#n� 
G��ߗP<�g"QT�����;�Y�w�Ő3	����"Pƪ),˟�b(g)��]��36h�|ũ9������&;I�����ll��l���,�����uI��Y��g��e��0Ɓ��YbL�H~s+E��ԢUo�_bp�kPN'��pg��[G��Yy�a
��,3{Ŧ�grW#��,x�}�8S�H��D߬Z= gc��A�S�a`&4�{���o�j�c�kc�ps�_%���1�F���{2��׸�^��Y�����uu�w/c���N�z�ƟOSt��S��4Ѳ��6���[�&w�ig3!��N����e����$�WT����U�8q������'Ӯ�"�+�o��s��El������>�'�H�[�!8O��<N��c���-�A�dA��&f������B�eײ^�3�7���"[��)X��MX�Ɨ2�盾��rD���x�hjt�'1���>(�(tc�.
l��ʵ8T��~��䋌Z���Ħ�1	!E&�徆��7�I�gq�� ��s/�F�:ZD��z�~gD\��z߬�I��5'+ ���W���z�4�)TǔA��	���n���|�A����5��0���J�>��I��7�-/�V����<�؝0 b4��V�f��z�}xab�'E��j��ȑ�{2r�a��<��Xa����첌�as�ȷ�U��o�#h��EPX��A��72������Gr��e=o8���)8h��??q�̵�L�{}�[<G�O2�q��e�̤ҮpO��Q�6ܾ���\Hs��ڥhb~�"_W4H,Յ&E��ڭ��д�(']�s� ���Y��x�}�0m���=�	�(QD�u���͞lXj�O�9��S֜�p�Re;���,�PU�+�2T�k���"ACH!�<t	z��Y��IE��{�O�=Ȼ|IǾ�����֡�u�x��9.�Ia��x��W�,��.��h�4&ޮ���Dk��a��\oH��U�d������9E��@�@ �7�H5�R���1Q�<Bn�J�͸',#�3��&>]=u�75b�:�Y���Pv,	y�	�)��qR&�6��M��eoNw��8�1��6^���)���fl�l�n��KF��w8�~{L��?�?>e�zȗ���A�F������1�֝'Gޚ���h޳}	nN�B����ʿU�NG5�R&���sD�5��U��TFc�ܠ�g�H���~�H��ߛ��/�}V�&���/{ r��ORzp��c%����a��K�k�U-.�������F�������B�?�[@۩fg�IH�(�-���`��� T���{�.�R�3̄�.��4����,˭�v�\���|jWSa����7��n��]-m�)&��٩;��^3!�`��@��������4��]i�8�u�#ʝ�^A,��&�eU6�'�I�	Cđ>��,ǿ=���"�H��!9a(��xR�$��ǯ:)��g%�lV�C/�B�+Z每=�=�4�O�"Hv�����He�_����{�Q'rJЮ�z^��@�]jd9��m�����ƽ�$:_����]%�p���3;8���rd0Ӥ�$'��D���5�H��B��o���1S"���7�xHG�L��f�˥��S�	����Unnb���G��n�����x���l赗�����0mD�i�f$���ؼ�i3��J<��oͬ�gJ��q^��|��=��~jYIͿsҪ]�	�н�|��*z�&75P�<�8*9���&�>�I�e�r��XG�s@1��4����U�2�E�s0Ww�c��^cL��9ʦ�<i���C�v٫ρ�ߜ3�C��]U�ŰNS�^��E�?�urw6>L���r�]�Ĵ<� a���/���y>����#��!�!���d�m%1M��n0J��Vi2��mS�6�y*��`��(䯗I������%UTh���dA��zg�E|_\W����Y=�mI��HF?�ڶ#L���g����\��"ѵ�K�ܞug�%}��ZW�!��F�΁�9���Fs��Wz]	��L-C��e#_�V�˝D�8.�\.�|65c|5�%��{̬�k�/dpw�bK���>l��A��YJ�0x�H��mb�+��Od(Un�5R9�7��h�,�������ZUM��
�f�\���@�O:E3��r�6�?��l�"�3��i�$�
O���g�U�^��Z��E�~�*��׍2�(�/n�[+�q�d���4��T#��޹o.&b����z���%��@���׍o���ۥ�^��Ju�*k����5>��e�o���#N���R]mDת�aﲳЛ�m0a��e�=l=}����mc�=�o�v�A4!�����<n��n����J� ?��?��C���3�1�N-�u4�o����
=W<e�I�j�3�N�s���g]'5ܿ�U��$��peM���pc�Y�(�	��j^[͂:�j��x��8����'ƊߵgQ���3�D�������K�ePF�]��t��Ǜ�U%BJL��_���V�o_�e�	u?���=�L�P�S����O�/�%��1g�P�����3���Cs�\�sF͑��nҹ�R};μ��v�%k�5�LM �t�XvJp��B�f��6��D�P�k��J����}g�=�|��Ǳ���M���UD���t������e�TR�	�������TA
�4p�A�gU�<A�xe�������,'���"\���В ��x�=�(0������>���W�d��&�̿�V�C�;�� ��D����j�jμ�J��O��p�ݰ�0��`Sv��¦��o3��WvY�+��ܷ�d]iSD��@o ���텪 �^�+��QlZ����	���qֶÆ�R�ۓX)�B���;~�P6M��:>�Fߟ
��M��s�7�W��g!<�� �AB�jV��Oiԃ+s9%��c�	s�	�T��`���}�$0Э0��=JGh��L:���E��R��/i|�ٲh!0tdn2$�b2ݰ�%c�â� �:�(4����2�g���ݳmK��
ƍG�����d��.�
���U�{�,n�
��೗��؞D���W,7h\����8��8�Õ�79��XEE�b���Vzix3��t�O�+��N�']DUĦI��@L����:g�3�6s��I.��������M��)�<_���>�Xǲ�����*���Iܗ�=1���XN��[�t�^��i������R����=k�3Т:B�+��G8@<��QBb�:.���\B+~�/N~�S�S<-G�Y8�*�b?���<2�Y����X=���G����J^�N�O�<�D(���C�}�j�WX���Ǌcc���G�����>�z�Ѻ
NJ�w�TKNi��]$h+�U�6#	>�<�=�>�Ԗ��uz
��uR3'LB�>刲�h;J�d�x�Y$��Kz����!�JukEj�\,9���C2�ll@?���Z�x�J�Η��XA�CJ����Z��9����E�sk�`�?!��g�EV�o�Q��*k�|a�D%�NoF��I:N"^@���u�D7�U�-'�뀩����Ӑ��^h����K�<��	��y��7�<%SCmuK6�B�my�����%_IV��2;R�!(��y��l�q3�E�g�05g�E�+�P"*�-]���,��u*][@�@Uߢ�8���k�{�8c���s�9)v�D�,�⅘#CAr7�G/oZIR@7^�3ee�g� n��[ t��#MZu7kA�o�W=�z8(�B���B������\��&�9��CN��ҲηD��&f�5�9s�k#?��#~(ɠ_�W��Eb>�J���cX~ѓU��;�HNCC	�ʃ�:aV��T�r���{��
R䟨v��T�O?���_\�>��{ҁ��m�.-i<�1>�w�������9��^�@u�A%��f����4���Wׁ�l≺ô����ѐ,��
D���Ҁ�go�v��L�g�R}�ѭ[�G�sZ��@
������� pkؓ��ШU�e��sJ�5��r
Lwp����ozN��:M@nX6�ݕ�̆Q�N{,)��ڈ����;E�����.8X��GOf��<��>�Unq���U)�s,(:v�)���''Z�>Y-��NJ����:��s7�c�w��[d�t�
ۛ30�)�h3瞊�z�Bn�'r�����L� ��>rULy��䫻��%s��!qz�	���f�I�Y5ª�q�vGB����ou��F������e�W �>��)t�6�<��,2��{��Lj��{k�@ 
��� ��=�w����Fr��[7Ao�.�o��"��a�aZ&�&H�>)�pƿ��% �pKѡ8���R�ᛤX���� V�%���l"�M7�B����s�j�o@OT�m����1��RC�H ��ajC��D���C�~o]�	�-�),"�����Tz��[��ڧ'))L!��ȹy�Ըpv�x��)V1��&lt{��jNZ3B�W��v�ƒ�k�K���@�5������M��p�a�d����BVU��8�x0&�:xik��$2'>��/cB\xE��O/X�\�%{Qb�j]�E����%�n$[U�vG��x�a�X�v1�×6�CW�6��{k�#
�H,[�Iy	!O�0䍎��3`�0{J�{?�h,����w�����/rh�[;�/�t���v�-ZS�=��}'g�x�����XR�fqA��r�������(ۯ�C��d���J��3��J�N���#������8զU�^2���S��� M*���>`+#p(���xL�`_�YbR�u��ͽN�P�I't-%�B�qB P�J̪���Ґ��&�'�����i+��U@�Bz�E�K1��A��張>�ԅ�h�	]�54^DR�K�N����W�Q9jX��3_����7r�	�P��KV"Ơ�7��TI�cY�zx�`�vO@[;�|>ɇ���c{��~�~~F�G�D�E�d�B���d�N��!����
Ə���-�]�w2��-��&�}����C��w���H���]b�N��݉c������yn�<�V9v_�:�sW����fB�QߐN��1�!��A\y�'�Y���8�P�_]8Gl�J�Qq')s1�l�k�N*b&py~��۞P�8��eը��IC��-��.�>g�ÃYP_�%��4�U�V>T������y��\�k�t���1�mɞ�Bm94��G�c;�&�GǤ�@^���m���x¹��}�j�\�nFe�kɡB���h-����ye��_�8�W�OB~����Ԑ%=������-���4��p����՜qy��і����Q"*��!�V+�i��'��a�V_�Aʜå9:�k�G�6>O�»��,�=R�F	��aX�+�,<�0�i.H=|���e���7��p�3R�<*uR��6��OQ0�m��,�A�՝������e_��6��HH��K��
7�u�N����_g����h؂�Pk��k�!��ӊ�,�2�A�ߔO5u��Y����/W���Y�t���Ҹ��ձG1��r5��d�@�mIMW⤋��G���t��c��ٜx@�!�/I�{R[-�$Aɏ]�[oizr�
?��O�$��q9$@,��
j�6��&��᪑�9a��|�'��=�z�b�����o7H]F�Y���+CU����D�[{�ԁH$'f�l�?&�>,���J�§\t@���X岒��T}��N�(4�vQѢbQ��t5��U�n�0�T��̀ޚ���,<��J�aX6����-��io�Q�[��e�����#�@lKPr#Ÿ"��.�~k��TKf�N�T@��~���:Nk_�����@	aG��_T�ḑ�
yV�Y�!�/�ewd>;�mlv��FYB6l����HjAo
F�'ؔ�z���m��ӳ��9x[a+��Q���v\2��V|җg�>k��q{����ݪ)0O|��6���@H�YJ)�۝.[��yo�6J����`fp��UTdq?Vn��L������4����ۓ%�;ʃ���[��py�T��wW�f����<y�j[�T�)Z�W����L����*���5���8���#�I5e�b+�SC�����ݩ��z"�$��L��;��MmT��r]�2�α9�d)��/?�e��M;�"�K�iRe(Q�J�*�
?��d߷	yi��8	�	cE�j��Wj��(�r��8�D"m�d��· ��,��6Qv�@�j��[z?;��}N*)��OvNN!����y�C�׿?��A�5�	L��+rE��.��n��^~H�X��Z���=��� @�����I����,��T�l🢮XY�0p)I�:�M1�CR��%�KXu�����P�`~t�;5h����wdX�ٹϒ����iIY��G\�<H�L!>�� �`�aA�#e�߉.�/Cyx��g\e<����B#߀L�p����)��F:���9n#�@؛�#p"6ȑ�����V��<�o���xz����]�h��mQ��V�0D�����֕�c|�'���N������M���b����5Y�/��|X�.�;���+�q�E%��ݷ8�P^F��.t�����F�I���]��&�ˤ������|$k�LOgD���"v�Kn�|��lOl�e-."T�>#u�7����7K���:���׋�������y��!�ӌ�ǎ)`ͪ��
���Z@#vn�ڃ�w!P <j��U@J��|�jtL�w�a��������u:��0W��J��3�������$�e�)n:�"Fe�]�N��NŎm�2��A	�Ų&�K�^���_q�E���x�x�O2)`O:�������cN��y�s�%؆1l����FE�&3C�pʻ��X�{��@l����s� *���veD���R�w�/E2�fϏ���"ט�e�r_��>�|�t�%t)AD�A��<��H��lU�TCd�
h<]�dTi~xR~��N�N���VE�X�v�g�0��z�R�+e�c���'��9~�T��M?o7Yl횤v$"�E�Rw�[��/%���F��8�K��#n;��"�=.UF�5��2��/9y~i�J��!�k�>o=
o5�qB�aQ�	�-'����$���)O�hXM���ڹ���s�J����13�Ǫ�w������[�F�:Ϡ�3)�Fc�Aų��RtD�sFx�;���Hc̜�9���A����[*�) ɪ�8���<�n�{]�^g򢺨��4�~�)M���5+_�ʱ㝅Qm^�V#�O@9�*�L�ʛ�5��ω�4._x��m���K�oG@m(~�_b*�]V]rXd]��z�6ã%�ܾۗ���z
_��;v�Cr�&��W�k}�V�CD���
Z^��T�	[Ax�ёw�G�[���$��0�o_칠��w���I'�@5cya�{���� �z��z�@v����&����S�` if�f.�x�o���!������* � �F�-�v�5f�v?�;�N�O��&@yu�a�@�z������5�]���q�K�]����g���\X��{�:��mcѸ�O�1\;E´{��Z�Z�������5���Hs$ī�M��Es?�%A}ĳ����M^��џ���n������uo����[ o#��ȓ(����6�)�_>�lZ��fE~<��R��$��A��:�^�f2:ԁԜ��A�T��un2p�N�E���Ჟ��P(��ixef�l��E��+��~�����C�j(�������sL6�7f~*䝶�v��̋�.h��IMD��hT�����<-Q+4��X��:�;�rۃ#uSY�'�9�غr5w���6WM�`h&=��]����*e��}9��w��2I�ʲ��cכ���ҒL�u4�=��<�	F|oW���'Qlt!5�����	[X��4�'�i���F}/��~0&�
E�T�g��-���<�wW�DP�}`V�so�9�=���؋��3�'i�> S�;�*}�$ǥ� �@�6������3u�����N����l}\r���6�I�7{,�rv�����7���D�b�,a����@}i�W�F�8̮Ĕ~�BY�cG�[v4SJ���b�w���p��uG�8鼔��1��cڸq}�~��w�r��ࠦNt[�,�z#7>[�U�S�ؔ���W�u���.f$��s�}O�������I�X3��kP��eB� _Ic�]��pl�����P Zγ���u�=H�t��k�+�Aj�)��V���A��̕v7^`7"P����,����T�S,y�u�)��w�6���]jX��'���K�]�@r����!������*(��q�>���G 艬?%����=K��-]����%/	n��(�!hW��
� &x��[����q������U)g� ���e�����z�#q����qI�����ޏ�Ì/�Lc��������F�t�ˬ�J���8᠏3�5�����Jp�cPIs>[蛝��4I�lHônڢ�.-0���xe���@l����o�{�O���Iʝ��K�"�)�Z1���k������k����+M�\�ҙ֚�Sr��^B����I�esf��Ȑ�1d�H��x�{i��N���ц��醺bx���_Zoj��-���-Hؒ'­��i��G�����9���V��|���i��؆c���m��?$e�"R�L���Fo�;�C�\�v56���W���!���R�⨡�C�K�E�<d�|��k���BL ��X��~G�m�aYz�c��\�����\��N�-��;�Ea�EH.����DZ/��6ө�Z��؇W�uӊL�埑?�y���LȧaX7��I�l^ݹ�l�v� a"]iQ=��M�-ѣ֠�}���-���e�@"��Y�ϯÖ2*���"9���A�A��#bg��f3����6�\��H_���B�`��N�-O�V%{����T<x$ג���e_����`��Y�H �b�R[�M���.E���l.:vM�A�TA}�e�)կmஉQ2ah��TX՝%u���ۋqZ�|� ���kGD���lt�V�w���Y'X���ÒA�n����e���L����{���m˳��!G���IJ�G�P��u��9h����j��3;p��}8�E�"@�����ӹ]QJdp���psN����')�����Q�����K+�z��&��z��`�>G��1W]�õ�V�G0���@s��p�S�����m�̫�*�����p�֦с�r��4	�2�^����ML�|�GR�-�n�<H�lڶ�yo;_���@n�4FS��]�rx�<jAɀ�-�㝼���j�7��1Zc��b�~�t��u����zOhN��(��qXC�&w�~ħ��4��a��,������K[vr���(��2^��=_��W~�S?�Gn��<U�����o	�Da�Z�J��Q>�a����Hu�?����-�oqQ�[0�w}� �{�*�|�+&�.�E-���|gpkKU�0}�}��\��h)QΨ�����MAWSatF&��)2Lu�<���@��j{���*��T��^�i�4|!H����t"l�l��#xǍ\I�Q@Y�Gu�}D�����L	z�3_�{��!������d�]�Z�+�����8#�"]�e��>r#1�X��BO��PWb�WX?ؿ���~���֓��Pd��G��6k�Z��>�NƂ�7 ����X�qax���s��S�:2c�Ya��1;�;�<�Vh��Q�����/d^��&8�(&K�fB'{�%M�Aq�!��c���DT�`k�[b�t������k�]!���!y5�
�m�M�8KkŻf�'�G7vw�GF:s�rjH�F�
k<�IM.��lЁG�k���Ǒt#=ֱ���ߓ�_�v��C�����ŉQG��l��`m���z�@F��Ұ�P�`O-TQ��]E�͹�@m��r6��&����.u3f����$�Ŷ?;A�.�+����N�#7��m����$Q(�A�U����ݻ{# g��P|��斗E���x���s❚�.��?\�2��x� �MR4��R��G�yd����vC�ɎV�hgi�Jޏ�6�;袖�
�ԝ���-�ַ�O��|�7��wZB"?��X�_���W�����֥/���\k���EA�<������V���v���������m�T�����t�|��k�|���	�L1��H�|l0�O_yuVA���ܮ�	t�F1�#���t���Cȹ�yNQ!9�1���\ lP�hC�NQc��C-��%�����: �B�LC�o�&�$��֬9X#~���c�fR+2�	)�A��C���p��gL�p��\�U���7d���!~2��������宦s��L����t-dO\�WVb�DMX��Ug�r'AW�*����/
�����q�z�w�mG���\<0���3�)�{A����E�)v�" 4��S�vK���n�L��o��&vעD7j[���er}��y~�E�P��8��gM��z<s2���a��=)��9'�&d�˕7�t���\]w��R�C�e�nЃ#z}Y�5Vp�g��щ��a3q��:P=/�]��:���҉hғ��3�U��~kЅR���/6���H�e� �����=_H1�F�}Ld�c���h��ĕX���f8gc>�u�h���근�D�inZAt�n�JyI��`���:�0
/1�ۤ����M�+�[EA���6�Օ�qv���I�RV���C�|:8-%�Kdo�R<�{�DN�PDUW�{E�P�8� �L�m.d�.���_#Ҋ�����V��v~}r��"��A���w�֢r���H��nE�L.��vf!�J�&fl��Zdg5���=�~��y�)�p�	}�=3����93���C"�^4��8��g�ې��	�(7��X���7A�vq[o��h,�-�8���ʲ�����Y��1q%`�zi�i��a�l�"2�E��#| ֟�5���.�M':+�qU/A��~n�zH�q�k������2��t*g�"���5�@���H.�FUznV��NGe$�s�}�w����R՘�D�>�ͱ��w���F*9T}y��a0r�?G�R`�p�4.���$b<(��r쟎��o!�l��nr#h��W�5���ca��NLɹ�V��;�6���IP^E�<\c�P��gUDKt�C�>����f�K�FX�
%	�ej~�SDmL�]�����,�����.;�����'؂��m��Ɠ����u�քW�
`��k1������n����Jf[*�7�U��F��P��8v�����gN�K��x��z
�����}�u�_:,&㮛�9ǒ���[[�.�UQ_q-۱�)�*�Y�����N��U�p;]ߗfPk��ڄ7�^�-��Ֆ��U�fk q��א,8�hUl�P�����p��7��D�q��e�/j������]:�*m!e��7�	��[����a�c�2�^&�Ž/�D���{w�4�M��&�n� :�C0n����H�gS�;Wz�'� �:���w�BAK���E����O�.�2A�c�~� �'~��'�7k$+4ҙ��]o繊_ �	��Y�����Tek�l��+6�®B�sMd)�b�A2�6QB�"l�{�E~a�ٝ.���bZ�~��!�s�Û�#?i5,�7ƪYy킭ǒf�����ޖE�sB�������N};�H�#)})��^��r{�%q������W�9p��b�l��� �F�D�5��h�mV���vRcŰ�WVXPk)�*˼SBh�q�V|2A�o�ȭ�d���������|{�3P �e	|a�
�Њ��^`H���zu��|�l�#J4��*�j�0ߟ���Y7$���K��F����˨<J���g������M���h�=�F��wti����Μ"�Դ��������1j,���sr0]�����~'�*���5\����o��_a/�+A����(�pA�ԥ�6ȑ+7�O�^���׭�cT��՛%Q.8w���/� <y�x�.0�'�F:�dp���`�/�V9+��E.7i�*k�iq��r3�D�͘��n�(Z�5 �s[,|�֓eO�� �6v>(אַ��w&?ba�e�>-x��oH�O��/dlw|�9>9�������9�)&���G�� c��ɖs���((�
U��RD��;
��!}�"*4��7��S�t�����x�YgP��t97k��.�h[�v�o��B˕��e�d�󡓞�����I�Ru�.�1�%�D+K5�|�����?���6�ƻ6��6t7�����W�l��zu76����Y_�A�ZҰ#/4I�L/t�����EE�Rں��\��H�Dp`;o(��N3ꀗ��8��?GR���䞶��;[�iS�������\�A�M���R�G`-}�|C�U����R^��V5��V	UO�D������kǿ�;T?��o�1���m4K�P����F��fi�c�	� �1U?v�b�_��Ɩ���5�W
fnh�Ŭ�!��c_�������G>Ō/�Br���S�A�W����ޢl3/�Ҍ2��<e�\��/�����l��H�m�î7��b� r��8Z�y��i"YXt�
���-Կʲ��^�}����/;	Z��5m&�
������C���*���y.��\e@�=�������
&MG�K#H�b�EP#-�kKqk�tr���b���n�;�g�BQ�a>FB�}=�W��Tu������(�­pl�_=~��$��!��Fzi3��u��6X������I�z�G6�|��K`�����E��y�;�A{1T�R��#�lzgZҿ�ZKÑQ٧��y��2��"�;��Ec`gtI���tN.�Tx��}�&S��?ZNh��vf��M���x�mV�	�\�G0�ig��;ov$�$������*"��� �R%� r^B3�c�U���/bӊ5ߧ����(y�J���3�����8`�tf�M�����`Je'1��7k����i��+Bz��'����?�@�k9�l�.$Le���y	����$ŀ������d�)�VYmbI���y��߉�t��9n���jᶔX��؉F�Ǳ��>+Z�r��J>'.�]�&�-��E'�|��ʦ����Vλ���A�1�w�&;}[��c3 ����W�cM֟�%H۩�Q;��;Äk֕7�D���p%\?�ZN�����M�>H����YC��+�.��;�wb�>�N�7b{�,c3i�8~��=EX�;�%7b~H�μ:��B�H_1�>#��_�Í��.V١B>>b�)���\S�[TG����`y}��ޔ�U�k��P�籅ɘ@��
�R�;:l�a� �lY����x�߷��D=8�gA]Y!��؇�fsωV�q�FN��t��;�*�X#$���	I߉�J �wc�aL�n*�&��]y�r����Q�>�Z������$�������9���#q��k@b���}	*t��􋩫_��CSS�_�=�"����n�3Lf-��f��k`|����b-ӿNǔ]�_������{��O��c�y����E��t�^�?r�׼���3f,�P(���nk�Wy�E
�\�%z�d�vT<�!P��ub�P���Q���T���<.��D_-�X_l��4��sں��\�'���9��H
@�y�7z�wў�3Q������싷!�@^5�a&��_��)�ߺ���	��C��a��C�E{��� Q-����Թ���=�̫J���>:z2�� k��_;��YPǄ��u��JSh��=�"���*�@Ui�4v��aҼ2��2:��%q�����dW��%��݇�q�� g9�H��*�?���G,XJ�y~�_�]>��?J���p�2���	�+>��3K��� ]iOI'��Ȧَ�6O���Gl�=)fȔ�<{�T�l�rѺp���@՞�ė�)�/�Ȟ��"ہ8{�w}���wH_�8;,�0�_�?���j.C��ɭ��>�CC��љşأ�ҡy����	�}#R��¢�gֹكg�-��'��l̲�Q"�M��l;5~D�o�@0MS�OD�BfHZ����č�'�-`4et��c��.5�T�L^F���j��.~�1UVۍ܆&�s*ʼ��q�e�a��}@�f{�446���~��HB�gӏ��{�.�,�?�#l�4'�c������d�k��p��<R]���2m�����X�͕b�E������cÇ�Ƶ6��Ky�d��U0f���%�>�����I�8�'��L2��4�F�!9����̉_���xs�2��T\S��v��4>",Lg��l�$��v��ͨ+%?�zf���X����K�A'��z(H�P��n�Yy���%�3�姊k�F�dƌ�].R��9e��Ơ�6Y~|~��tn�Vhc��("�eo�%X_L+Ǣ�	y[���
-3V!�"bA'7h��嚼���J�ჩ%���e�� ߙ�8�	\��ʓ��j^2�&��B�L�$�����Q�$�Z=�V��_s�_(�r=ɇQ�;�v[F�&#!-�A^����0E)-����D��m�+ç����]G��9.��8�gCQ�Ǒ�M����)�n�q����H��3����P��㘷,�]Zr�9��H#'͂��~��,w��s;Ư|�7@I�9Z�����&���
K�&�o��N"�>\O�=*����M�FeS�J��۹�n#�N�Sj�2u	�n���@�]aU^FB�ߒu}���d�5��U$-����xIYěO�v��]�O�p��r`��ݔ�-j;����8��-�gv�&H�O��0d�0���o=�o9rt�Z�Z�w�=,�U�pA{����08�iC����t��b#`��nT��k(U3"9;|�+3�5�O��*�,�@������ݬ�,斶�A���dKw���j��k�b0��P8D������}��G�gT�F�%������&{��/\�gb)Z~|F��<�dt�Q/��X��X��tj���$�O���{_�*wo2�������Df�Ɓ¶���bѐ8�`{� ����L��;�"�u���*�6�y�-���>$6WnN�x�Z�� w�L���n�_��'�D�uJ��-��&P��1�P|�_ռ���(cV*:�S���f�w��T�6��.��������N��ƣa8W֏����������Jw[���h�?��������GƏ����Z�(�#�C�塘um4��Jj�:eO��:��:wƊ��gK?�{�w�?^"C �W���7Ô��<�ʆ_���"��`�j%���ʷ��x5�"�T7Ņ�GP��C)��~�9�N_-�R�w�BE�D�I��?JF�<�������\F ~�`B�.f�]��zb�AA������MJ)�9 ����#Wp�:�C��;l���UP#�"�1T��K�&O ��74�9j����-U�ј&����^�k4~��;:ק��s�Ҏ�����Q���e=1�w�+��G2�ѭ���*Z��:@��c΀�7�T�ʺ�)N�]��hӎ���o���gNۑ!�%N�P��s�;jh$<�|D�[b<��0?K�Mݦ�r�4-���}"�Ža�.�Q���hol"�O֩����U��I;V A�>�2P�"����F�x����W�kUI�ͤ�������i5�L
��=r�(���lm��ϛ�㪡D�&^�0��c����d�y��>�~����ףr͸�L&�'{L#���X����w`��Ɇ�Hx��pj�g6a��8չ�}|b������0����a�2f������P�,A ��U�	�Q�1����`�SP�?a2��h�jZ��>�vb��\B�buq2f��`8@�s����v���"��Y��; 6ޮM�tq�>�y����as���c�1j>�x��&�m�H�|����~�2֊���=� ���'}��S4��o���=�[4*a�4��:Ѯz�͋k�y��b䢥7H����0$^����^���%�f(��[�s�-���E��q�lB4ݮ͕��񺛌E��`f�����-Q�B�MIq���n뀱���;���e��bc��ʈQ�f�&\v�F���q����ɊQ�+�r`#1m<�����e�]�Y��TN}s��`�[��:�}D���kW�kP�b�*�Ifи��} �}���<4s���j)�M�n<����=��r��O�^��9]�a1[�@�X��(�,Wbhs�8��i��!�(eP����(��9X"N��� $k?��C�+(<���.�<�_�0qj��V�ƪ�Q��KQ���biD3`�rG��{�~4z"Gh,p%��S*�=�%�/x�DӬF��E��#\|.g���b��y�A�(�Y��A��J���s�mp���tqs>�\"�`�/�/����KD�}��E�MϭՅ��F�Q�Ü��]�9R��Z��A �u����[��Pvk1R>[w������	<n	[�RE)�b�o��҅<Ո_�'�/�E��T��7�G��Q�'hD��81�_�D��Cpi����w.�#��l��Æ�/f2Eh���w9��y�7��iL��5���b��{b�R����6�6����:۶�}Iz.�5}�\;������m��<  sￚ�7�b�rآc�|s}��uEX���ۈ	�^8��`TZ�O��r�J��2�@�f�%��C��.𩶈��`z0��^-U�U��w~��TsyyhSC"���(O���2�`�pY>�>�(#L(��}ƫu�q�ž�9j�z5�`L�ڟY�tO�y<���z�a��kp�^	W���2��{�۪��[�yUD���y�yi~��uS����AΟ�M�#d���JnƐ���B~B(A4��i7��1�`�Ο�[��-@;��^�E�%�6��5B�(3$J��٨�u8K�0랿U��U}?��	֩xƫ���jZ��<x�4x&���4#{�"�B�جq�¶6��*ٗ8&s5��f��&��r.��qD�lj��a��ގ9�C�{C�V+F-
]��`{e�Ejg}x	��S����4��kn���'��Q����Y�p����D��Z\���r���T�K��fЩ��x ^�o��DE	��Σ5��|�'��_x�d�����߆jG�6ɝ��m$A�p
��i:�T��Y�L&:a���O��Q��8���ug�[�ΰ~h�Q�OB���|��t�QID�h�}Y��'���@&|�Z<�\��E�W#�SL��c�&@6��ȲE_��ڂ�.6�7�!h}����)�zbծ�nQ}���uW��,�����R�`�nC����"��`��wP���K�����ئ��k�=����Ǻ	k�0���+-?WdvCE��lZ��_%�n�'���|��������Ļ���!L�d�fe'�>r&]3�4���z�����.z�i��An�^;؃�؇�(�h��t����2/�b�e�cӪ��.|��VNC�!��Pd�Y�~c$I��O�\��nH�
M;~��X-֜����(����GI�V��ԷI��P����zN���eqa��H���c#~���A3����b?p-Y��A߻e�Z��/|�n�g/N�����Ti�>�~Hε�C������e���q�s2X����ŵdOpc���WwU���n�u;ęP� �k�
���C�q�����j
Jb:��j�T����s�G�g4��e�jm��(��ʘ<�TE��_U	�gRI��jl������V���i�������v7�����n�"%$�����2V&��fiqC�j��?�n1�TF��@5Ո�h��5X���ۊ���xA�2�$�w�P��c"��7�S�"S�y��Ձ���z-,[�w=		
�R� �|#�Ȑ4o����T��R!�	���s���f�ͿB^_����� sQ�!����pS�G�g'ȵ�j�%2W1��"c�~�:���_M�ʫC�@9��?� ��T����o���R�+j,\~���l��+��M
��:�+ʆ �ЦCx]�|�GTu<��B�b�U\_�aZU�+pۡ�����m���Ә���q�7R�!�05�C:l,�r��y��m�R�7�/Jt���2 �"�M�G|��g���FL�_�1�a8{sPE����,
�BV�����]h����ɡM�TC�ⱸ߀N��H ���q�+~/Uh�N2��lKEc��Ѻ�=�sM2~p��2���4���2��M��h"F@ujm�^�����ۦ2�*��Hf����bq��i!)��zT�W~[���t(�Jǩx�	$qp?�k�[bE֋�Bl0�R��}�xU���./��K�=����b�V�d���.F#��ii{�<R	5�g�V{�](���|�2КHj܇inn�X�-�{�DZ�5e�%� F9u�:Z$0��l���N��ԍ��A�m<Uyk���^�t^p%�\�!��L�l1��lx'�v�P,���o�!Yx��n�9��$�P��ʍ�W�w���q�<?�?�c��\�P6�[2��?�}�M�6���3y,��s�8���fpPfI�A��ߔ�_�8����6�ݩ%��A-4�������^T���2@�j�N[�u�p~���G��8��9��4�L� /��0��kV(����F��D���"�4'j��?:zv���Cs{5�g̠�5i��L�$�@PG���bC-�/d4c�&����.�B��̅w��e喋оi%��O��`j�����b�����U�enT􄘟ReO��5s�G��Il�&RC'9���{'����p�-�]#�]���`	�.�(� _�p+S��
^4��x[��ý��"�LpVV?�W��^�L��}�����Vp,�7/�L�%pస_m,�;�����3T��.�Lc��"�$��b\��?�a�����\��?�`�.��i�,娜^�b�愒y�{��|g >&��V졾X����@�-f��P�N	��}�K��o]<qC��P�%n����9��a�o%�s%�} :��$��h�-��j�8�T�5F]:�Q.]T?��P�nAPċ�����(��e\���hĤ2�%UPq3AF��m�o�>@�ݞi���P��P��p��Vr����U�Iu,4��<V��U:;��k�p���J��5Z�H�]OX~��v�[� �.T)���ZT`>=Imd�Z�!h��$��I}���	3��3\
~��_�Qߴ�#}�yR�}Z B}W|J�4H����{;^�Q�"� �#�R��#h�w���� L^�G��V���c=wx6�y$����Va�.�|ǎ�&��`�ɚ��8��Pf��h�����I$#P� � �PeO#�7K��qM���
2B�@a)�HV��Dx�v�Ho���}�޲:.\��zSE�}d_�i�-R�K���꿽M�ad����}�m8�=xI��s���eA!�-�I�����up�Tk#w���+��ud�0�cx[p�ɥo\���c9\��u��\���5��K/�L.��%�e鍓��G�輊qx�ɷ�B��hW�N��0�a. �c�(wj��LK���9�%���i�[��^�ƣA|R�(�h� G�TW�8��;�0����y�E�
Rd⃓����75a`�j���l��
]�ks��^3�?�|+�4 �n�=���kᢦ#$����j�����Ǳ�Y)ig�%"�
�j�o�;��!���Tb��f��b�I�J0I5�R�*P�.�
��7]��r|�(5Ys�'>��?�E��*є����:#9��;,>y���n����@ʻۭA�Y�6��](5'@{(���5ɥԡ���� 0�_cA�|�Gu:*��0^�F+�tf#�aJ �+�@_�s[E,6��#�������u�[@ܪSSf^��n��Z˹l��N������5�݄�����x����g~\Aoײ��-Ȏ��?|�zH�|u��Б��1�#0�4_�}a�N�y��y��*]�>��van-��P�v[�U��ॢR�sp[�N,{�FT��<�yyQ�M���f���Z����T2Q���K�rs9z��6��� ɧ�!�Y�d��&{5��ڮ��6�;xK%(%�ڲ�����.Fi�a�%K[锋�8����Xfx��9�Y�XL����%#þίR9�
ra� ��s#4B ��vdJ�>ݍ��T0���:�do`�X*mύ�SJ|(=�^���Iڧ��1�Ӏ� p$�/D�[�f�-(B�����<OO?�n4�3���\�[���g��2���� �^-\�N��e�������s��J�׽�=��)�"$܋�� #�w�A�D�a��rkk9mf�SD�Y�e������(�c<{��n2��rFj�Qw��5rZ� @�sM!��I�0�B�����������>ʕ��miNi`�&���Pg)�j���)wa��ޫC��T�}�x��߮v���=�~�N�W�+lD���@���0�eq�Ĵ-Ӳ,ё�m���p�놳���M����T���l�o�7i}������"O!>�N�e��V���3������J'_&���W����w�tj�7�|��;�kg����ʉ���N1�;C��� w�<�V�6���¥)@"?��b�4��2/U��z�M]Z��y)�~Ӽ�S���&:��ϛ-�g�-����߉. �y������q��|��o���ΛY��Y6{�u[�byv��eLT�2�6���)�8�q:�P���_B[ݒڙ��RD/䐄��_�a��=�A�ЧA2B�R���IȍF������.��5�<�"�E�&�=qoΑ)�!����[���LwQ���z���VV�]]Ve!����8��#�Rq�]r���׭�8K/cpÂJz=��z4�Q�y�FR�mȆʥz���%O{�o�	A��3Z���}�_�&�*du��cmѝ�t�.�� ��@���z��p�Be���ˍ�xYHҀ#��t5�>��/�2��F)bD�${�E,5t��\ӄ(���|cn)%׎����.E-|�t�_���s4�z?dS����%�"e}�W�� �^���F/@l�qd�X;܇���g·Q.���Ha|��a\�D
�}�М		&�u�D�e��|h,��dct2@�O�S��s�֋`0 ��饴;�
R5hogQ#�o��}�ϕ(P�c�+��4�KX�T�3�l��Zg�zy)y��}���+�Di<l��T*U�	cXN�q��9�az�����K�#�����Z>�CB�5�[�w��0��q}�V�� �;���F�C)��b1�Y�QV;=c9�V���N�����L�Te���̚�a�W�Y7�����X셵�4�����Y�smC���$^F���f��H���l4���)Mv������ju�� ��;9���e���:���j�G0<@�O��`�M^N��[u��^`�D���u�~
л����#�10M,좀�ah�xL�K��r~�#u���V��|$Pݹ�A�u�G1�QC��ⵙ���')�T�(.Y>��Ya%h�>/��w]w�$�E���|�2F��*��RO<"hLۄ�K�ݵ�
�?\�u���ַ~�Z�� lO��U��"EJ�E�<�o�Ím �� ���_���e?KU�f�t�����������Ba@�g{�2!��4K�Y*�B'<.L�;d�'�34Xc6i�9��~�Fu�$�s���CHbu{!Lm�ү�f�K�`�:���6G`�#Yܷ0<z�(�:8��9&�4�����xd�|���7I��+Wz}ы"���ozͼ�ɶQ3��+G�=��B�y�:������e�F3�f~�W1��+��$�g�t�R�B ���8gq�t Q<l�w����qb�i�o����Td���[�_��DhG���`ۖ��wH��В��3�;�߇� /�#��:�q V<�#T����bJ���ֹVI��y���28����ȝZ�Ӽ���s�A4��Y��U�7wi�
>#�+յ��<�ݍN��q�� ��`�؇_7?/��"͚�>�g��"�ۛZ����!WF�Z2�9�{���c�I񪠨{KHj�j�.O�Ο��[Id��Z��Ÿ�-����E��ʅ���^���V��D�h4����F�3�����3�͆��_ӭÄ
,�l�1[g�4a#d䰴�?H��N}Y��p%8JX^�J��r�W%�}�o`W'�rlj�,x��$M�Mb���-������p����fU��0��c��".P�-̧����TM��f�<�	͟�<�թ`�0Ԑ�\��%g���t:m�t��^��g&1m�����DC[�L����`B�������9L�j�Ս[��?��8��)�N&�u����0����&��B��
1bO?I�dp/	>���^[OP�W�qU��ԓ"j��#� bo$%O"���2q���;�g��Z���A�*���1X7��Bdlhm��^B��G e�ggL
U����m"��R�f����$TZ4Y���ƶ&�b˵5\���t�oJ�Z��n�"u�,�a�s�0�?�q=�Pq���ߍ�Y�T����֠���{z�R�A?�y�-��u�t�e��`�����/j�F��4#�A�SV�������Ň��h�Jx2SL��h`0��lo^��f����l���5�xAߏ���5��c硓j�����VX|'|�*[1���ČTwO�AQe��q�i���Lb�M��C�@�Q�<���ڎ�u�2�[�9��,�_ �j�DC��U�d�����5���h�-"_�M+��o��8�1���4c;	�c�*-�Tl^�-Y3�s�}��2��)q��>[�\���Dۖyʼ$ϪÛf��)@E۹�ԭ[H��*A���4zs�+�γ�*Z��7�J�{��x�?2�j�ܠt�(��%j��^��U_�*	��W/s��Z��= '�:~l���"]���^�J�����r��N���Pb;ߢo2l��l��˿,J=̱]C2��=�h�5��9���=�]?�z��Uz��6��eXE�N+�f������k�U�t�\YY�Q�K����x�8�u-DL�-8+�S
i��,^G���bOj��.o؞�;�ֿ�+��]�Q�U(�E���Vee��2>y���)5;�N�˒؈+�+�
n�qH��w�F����V�ü^�=�E�����O����2��J1��SSw�ZY�-�U	��U��s�.���UQ���i!���¾s�z0�8kX�獸�Ll�+�u��L��^��[l��>u�`}B��V�?����lu��nk0m��{ �G�?��IL<�Z�	P���j���|�S���A��E*VW�����R}�ԥ��׫a��Ψ�P��c���(%g����(�~���%����f�i���1@1?ģ���m¿�������뷜�ɘ9x�El�*@��Ks�c5|kht���B�{�� ���oeړ���/%��t��0F�`��T&a%��.�Q}��T�#�J���+����v<�u\�������`QV�iČ�l��V'9b���0:�W��}�� �z�(�S�D��̯+����E�%��Y�pq��3IH�[b���Ll�ؾ+z ����bf�+��2�o5�<PA�W9��'F#M8d,�Iot�	Zm�]H�T�!��
�_�nk8�.� LH#~}V;�:jxq]���2���
낙 ���f�V<�S�ș)ù\�p��6Z�f�:ں{��,O��R�ZI��+�n�SQ.�g����	��I�]ؐ�Z����f�'�cw�Q���B���9/z�v,�OS-����7��U��$��[���� a��Ye�9�!�!}�h'����a7�V}��h �Ň�#˞���-m�	`��^�U��������o��<n\��6�?`����f��|ɏD�O0^��j6�4��)J���PN��{Ĭ�O��7%�"X0jp��l�㼤�!�P��s�J��D��f��:�K��q���2����)�j�/���-�"�_bؾ��7F�zo�"v��.��y��L}�i�+�Ky�ק�+=���fC�hX`h���FY��� �f��o�C*>{� �p��8�z���#Fg)�����՚>�\Ξ z��&�-)�(GNj�l<�q߾Vh�msX9(N�z.��r]��W{��k�=�ݕ�O
������
��-�&�p�׻�I��
�~���Os��Q�����:s ���v���R]h<�-[�&�p���g���d	O�oK�P��_}~�>��!�K�	f�x��ނ[�K�d*��L�L_�.ғ�d�o��LW2ߖ��4,�FmR��J(��J�nY^cB������X����}L�ќ�ЃD����D�+{�9J�m�5�nx#5ծ��K)O��-拀w�V�m�_�4Qu�x�6� �\�2�@c���������I)%j7��?,A��'f$L@��Pj9Q���y�P%*3\ݞ�A�;8��N�[��A�寮�˶�S1N�^c;�)�kZl 1^ [ f��]C;�~KWف,�у����D"#^���>Q'��~[0� }�3&(�o��֝4a]��s��Ͽ �x���R����{Q�ѷ���\U�I�Ö�N�?�����hj)~�EZ�Ҕ�4f})��N����Z�?0֟@�j��)�S�M鼩c�d�=�0C3��۰3�Z���~K��?���Q���R�M�7>�<{A�Y�#c�Sv��!q(�U�
�ֺ��g���׭E\�kur��(�+\EZ��e����n��1-�7L����H��ΐӮ�j�[{�l�`Ə�b�T+	�"!����!N�T^q��1@t����T��s�9��Q����_�dƅH�dI%�R}����5�K992L}�m�E�����-_檎��	��\���i�K��4?�w`t�:�s_	`��\�����h3yG�gj��S��2��$�U�
9���qy�!ǗN����33�6�(S��ì�T�,#���6yJ��}�!�E=�ٺ�By������tW�#m�j��iQ�et#��ݑ�X��4�I��c�"��Ҭ<��L���{���뱽dw�QW���Avo�F��#D�=���\�X�sE7���"�6��C7ݭ��:��FZ�*T�:K���W:Xf��=K�������B������5�lok-���:M�E|�i]T��眵�}�2�&�n�����Cۮ�r�M�`��x�.~V��F��X�֭��Z.J�ʆ]��Xc���w���7i�l|,������z���<��\z,Y`سʏ���M݁nę��o�>\�qd��@�^�V�A�qg�e|���b
S�r�E���F�=�Vb%�nl�F�3v�>%�ͮ}w��#��Z�0��U5V��A�a���/V�0�}�h�G�ں��y����l��y^'"�Gyp�U�qh��xl1�@a��VХ��+�;�"چ�K�����oZ�>
P�:��N����������?+��=O�ى�i�k�ٞ8����a����J��>��D�A�z�t�'���}WEa�
Ct�;.���R�}w�O�/V�>�sQx�o���w�{���UV��6~���ѷt��m����^�g���L5oI���zn��$����$��QJDbh�;���#^��9A��ƃ�$r��T�u� 6�����P� ���HYJ�^w%��D"a�\V&�����o��96�
|���k*J�Eȏ§V3��J6�����1D4V	��"�X�e\@*��V�_Q�a�ޛȣ'1�Dק/�=�|�Py6$���2��}�%_��V7N���^Y�3^|��V���6y�+�屲,�=�`����PK��k֔QĽ^�~�2..�`<��	n�'�UgK}P��Í�ZoE�0��Ӧ���[<V
A�W[��|�og�<��grW�
B���R>5�:�^<�>k�HQ��R�	J}_a{�"0�'ǆ��.'��~U��%��f蒟�sqfH�9SMc'�L|������Њ�j9�8^4�V��Dhh6x3πVgtqCؚ;(����
i)��e���h_R�/f��T�pl�hAj�5�\lUcI���P�F14H^J&T��/�v�K� c��Q�@���������c���R{��R�E+1����F�\�"�rYD�lc�Y��������wX��rp�:VN^2YJQ[�Rhd���ZNp��o�
�i���?Y��퟾[�M��+,�P���d��f)�ֱ�O��xi(0m���
Pz��_�I�i$}��>KY�h�s�8�ۈU��������O�� ���".?)H�o29�+��󂿦�P/�ޖF��S� ��3�W��B�j��^��E_�P��T͖�e)��E�ͥ	��P���i��u��^�b;�pL�kϴ'eq0v0�흢��x�n9��	�A��P�;jI���Y��#�CY�DOoWau6J��������;n���3��,�cЧ��Ǜ�Q��t>��s*��u���$>6�x]V���U̬�����R�Wl�̟28��� ��c���+�����<�;�q��-I�$ȴ��@`� Ib��+'`1�}��z��Q���K��m��P�C�i�J%�������'2��笖����gRRL����=L�Ke��q���7�!%lyrձp��A�n(�m��SԲb��x��l�8��Ԯ�I��-	�eb�*��V�U<�%���J����'?�ͦg�g�Mm�Uq[���y�Є��H%��/�܂'	�*�@\F�fSW��6V-�˟6ŉ���3.�6�5�z�Pj��*���"p�VEˆ/&���ƒ�F�}���ك�k����d���$��0���dZ���;��i��"�j����]@yأ���f�a����E��b��q�:wa!���Kc�)J-L/�8�`^�B��)�p�3�t ͒`r,�<fe�j�B�W+�Uvqjw�ާ����-<��)�_i�C.��l{EB�3��ՓP��Z6k'�ԾZ�3��DSq�
']lՄ�����h��%Ї��C{.k-���!C�v��q�����:����s=E#B��y>��A��h�k���=��X�{��g�('�O[le�S�ꜻ���a��ˀ��IAm(l�b���.?����_%�C�wV��X�<����H�q�R׃�~
��d*|֦5�6����c�b���8[��2p�?��&i��`L�}���_A�N�0��n�X;�Y��t���y����|��v��/������k��'v��Mn֙~�\�yop�]��G�j��"V���d>�f����j�5}�L���9m��{Εl]n�~��,�A��x�~0e�F"q�`�w�}�F=0����a���p(�j#���s���(Y��6��1��Xײ��3��"�sR���I���/G���և�\�-_Vi��� #�;��l�p�����6����xC�i���ov�,�C��/�}�1XF��$S�'��E"Qwna{�rt�H�����R�^({��ˀV m�!Q�'T�L�s�wAt4y�Z��Yl��a��,�ߝ���6]��9�s�F��>�/�J��y�+���Q���myfP��I��o�}iC�Y>��A�7^~���Nma��-7�S�[c"I�J��8�s���Zu�%�j��\������������F�n�4�6-,!*�ܟ�ͳ�`�C�'�U�����*�����T��U�.����K#�K��t�	�bS�5`Y�C�����:o����X�x���k3|�U|���mE��	������eiY�3�#}@�vD1�(�����O1i�I��!�z��Cp�~p�.Bo[)8QO�y���05��TL�$�c�Y���T����k���E44t[Ӹ ����0��2�%����y�OJ��	>9��y��$q�TBf����R�?�#�P���G�_����츉�9v�Hζ/����\S�a
ͥcH��	`9��	�~dPO���1�ZxGL��~Iw
����WI�eDwN��5/,f�Y��E��q��(g7��;	3Sq��ϕ�b6=3�:<��u\0����*��������t�����)��ex�jA���>�{s�秘��(��C_s����;�%��*X٫�0k�� �F�.�Z�����֞0}HhK�"���qT.,E^J��#_8���.��a���=v-IIj�����n�c=�<�����]97QIϬ8"�;YV��b�-��W�Z���Z'^՚�w<K/���'(�	��3![}Ā�Ų�Ep��R�Ka�պ[�O�H�^�x�(q��B݅��zκ�*����.�>���~ҡ��J%���|�a]r��D����������G�z�^2�WE:e��t�[6<]ln��U���|_�z�۟�i�J/��L���R�,�c�������e�	��`-j*OE�d!s]���^B)�F�Og�����C����>�_j�'tdɲk�A���s4��:�6�z�����M=qM�dB�����ʶ��$�F� a��JQ��X�N��'a�Y۳���M���C�+m  �Ċ���v��Z�	^�7�.��t��|�[���Q�I<;��z����C�9J~ϑ���7��G���*�h餴�8��|>�Mj����_h�?��Z;����)�=�Q�'�mA�!�G�Hڶ?�f)���@� �C��L,���7���2���=���d�>%fz>
2���*\�hx�C��Mk��.�.F�,�'E�5`������6W�]@'N�s5�6�_C��w�7��P0R��'w���ms��]��@��_���q�2;�gO[������|���φ>6Dt��+l'��'� �*��猥H�~jh䲨�8

0ێc{��% $�UPƂe70O����S�Y�Ѓ�������'���OU�h���Af��:�VK���� ��6�k��`A�i�������C������3n�{w��,W�u2Tv���>��\����'^�f��0^�U9b���>4W�r��X��u0��⨺�،*zrv��������G �Ϲ����G��\��!��C�A?�j-���T�V��"fcU�Ϗ�=>�r�=w�8�]cA�%3�"�O��ɣ��W@��W��l�:�w��+%���>�6�Z9}סpiR���]�O<�"^<|7.1�Cڌ���1Y��X}$�w�m�/&M��8!n����!0���-�#q�����QUcps]mF`�BI��>>�t
��w��w�$'��2��d~�H�0U�K�����p�"c��X�!���#ֵ��߯��f�qq���Ȳ��9vCiF�!�,��Q����~~l�mi����`�*�Umkz���~��gJ5�ǄQI4��(�2���T�����=��;θ"�@�$\vJ�@0�D+5�X�SC��4cZ�&�i��𦴂�NM��1ʀ�yl�B����!:�V%��C:7�j�z�3y��va��I��oq���:;
��*MR8�wF���[����t�2���):X��q��<j9R���="_}�P�����x��Rx�U�|`ac�rD��֊8�&k�
3��?;ʳ�G���?Փ w�U��R��kw
~������奀��h�=m�^t&苡(ҪS�z����#a7Y�ɜ �z�ѩ�YBX���\�^ۇ�MJ8A� ۀ�:���Ϧ�� sԋ���;d.sE�P��zE�	��|ۍ�u�<�V��z��c�sg�[!�@�H��X�MF>��Hl�d�6z��Z+"���S��!\9<Bu��鮉{d^�����X�)\�ݛ����QE�>"���y�ʪ���؟�P����O{A�f�Q$(�vym,�g	I\�y��N	?0l����>��~����Dxt��K"�ίK�Zg���K7�١��m���eݗs~�#`}�]��!��]���p���H��B)���G��۽�N�z��P�|���=�Z�f��ba�!���B��Q��푂�ė���a�y�~&�E����ƼV�Bx��L!�-9�7ML.��\gP���8R>��0��`�e3�1�[>V/"Gv� b#��n0ź�Y�I�'LR�v���Ş����SA�����0�=o�#� ��s�`y�3���~ej���2	��T{?��4���_������Iix��(G�$�߻&�����ŽnY*|9a�J]{1�&4��`��;�q#���B�
�1�V1~�@F-��Q���{f�B6��.B����N'YP�Ny�:S،>دE��o?�j�(M�x���
���ڵ�c/g���Gyև��c*;�U_��J�w�#�zj�.��c��Or �!m� g���;��|�?
�&��p�f(9~29�LDs�[�x�a�Hg�K�9Ȧ�<�&�h�Sd#��0�M;�D���W�t��_P��r⸤���VW��B2�Bț���3Lk��ØC̜��N_�9�{~�W�c���媦�å�*�(i�*%���7�Q}]����N�$�V�͜H2���qe�$K"���f�~�kj,�*;b[�}M��(:�?)3.ޥz{!��<g%�ӄ��*�U"ګV1�$C"|y!��5L��교�!u�q<���!�AH�yg&^���_׈�%w����`����SX�ˏ�9:ٕ��+wLӃ�L_��K`�\�<����[�gӶcZqܓ�0��П����v�������*w�3-X����������OnqG���h���~�gsq3��J�0L�܊�+�������}�'fgF���M�43'ki���Y�����8!�*���pt|	�����a���@\X/�k�?ꗄf�f�a��	����Ӛ�w����yH�	����|'ŋ��|SӦ�]8��4�/��+5jg�Eh���Q�(g�z\����� حG/����y��厨c�5d��|�����}Z��5�bP z�u(O�p��>�V�5i�����>,�b�y�O�)��9���>� �."���L�cZ���k�f������%�g���>��8�rq�t$Vi\h����8n��`�r���U8���������N�P��V������,@pΞ����,��}��+E�s'�����ٺ��.A�S7�#�^��ي���A,B�^���r�c0V��ǘ�MFB{�ǝ�ٕ�ԏ�o�&R�E��(�B���=�]��۴E0��4�Mx���W�䲿�=��� g��g���&.��M���q���6�V f�������FT�]�K��EU�I\b=�´�%�X�K�j�Lb>�`���<�
�gy7]9l-����r��SS�Z�(�l?b����L���^�-�m�SA+ ��S��d���3M��%YX� W���G"[v�:	?�ͩ��bH��s�1b��=tjw�vq��|[&G���+��tg�vi}��[-��w!(4�_`�aſ=�\B{/}�^�� ?��:�:��֋4إw��bi������-����
4#�kX`n��/���V|S��{ɾ��Xq~#>�j��@`=�����.���rSd%Mk�_��2Y#^�6���톋����+��P�6��О�a�����/�/�\o����t��>Cս-�H�))��ʒ����C���@�5�<s����@r�����D��0|-��;�{��9�����O���$};c����5'F�`��K��|�s4�q��tA�#p���M�<&uӼt�p�k�Ż��~��Af�����w���$��Y�,�
U�W����6tOa?�y�9�J�3k���%w�u�+�3��2zpl�q�����'���/��I�:��Ρry�|OU�r,|&	n�E��qHP���H���Nh_�2�6C�*��N�r�6�δ�L�U�oҦ���l�<%Qס]G��������JF��\��2)���)y��.��s��Zf��G�������,f�.�';�eF�0��_P�>U��D����@��n�A-�%�1�E�~�-S��zU6�P�^_��.�Y2�Hbp~e�n�)�����5��	�Ƅ'�PN��Cij����}�eH6��'U��' 0�.�>��X���ߝ$�F!�<�������È��=��R�}��G=����X�x��*���^�џ�)��ߌ�@#<��_c�;�<@�����ͣ�Z}��3���OuS��9z���Xr��̙�-�{�����>iN"L�Ld6k��b�7A�v�&���L�M~�6|��܌���n¢H��+�����yV�@���H��4F
vI��婳�a>�M|��P���[��C�'�p��l-�Ф�=���OW�!h�	Y9��\b�)�E�#PXn���4\���'���IwzFXieL2|�j.� YC���gX��f`B�20�5L�@⚸����@�̷`���F�!N�d�qV��̝+��p����5�z8���C�ׂ��T�i�JB������p�c�(�\�C�'��ʋ(����Fuj-�ɃG�C7�Q��!�A�=
��(�/�o}��;Z��1r�_@$�o�[1��W�*T��Xlq��OGT\=F䒒j@�
P*7�S��A��$k[���W�o����afO/F�F��gq�rBrA!3D ��=M�\���Bc3u��6]��j.@Ѭdh����i|b�'a�d����Q}�<^S�Z�Z�L8xsW�F���>�c`t>M�Ք�}Z�UD�s�.�1=��j��������HIj���	��P������X\���';���Ƭݕ-��]�h�t�Yp}������� q�<�B%11���q�nF��t{UG��O�BQ�7��7�U��	Ӌ?6g�����B#ђ�rt�R�]u�^&��5��(Cp�`.�k����/#Ҷ��4�f�ϴ����Ÿ�� ]�m�{�6��1��%VL�S����i|�� �OW�Dڠ���\Pz8�������B�q#T½��'�ܔ�w٩�x��d��A���㣦'BJ(�>g�O��3)i�ˠ>����$�_����}t����<���~]	�⹒x�I-�o��Q��9��9�esB;.��C��f���Smz���.��\��u�mN�s�z=�����
�q<Iŉ_
&f-)z0�]��G̞�ټ�4���իz��m�w�$k�-AŽ.��&�ήXn9�o�ǳ�����&�)�.	_+��i�� k��M7w����Њ[T������a��l�C�����X,ǖ9�� �Pa��a*g� ��������û����͸}P6w�0j˛[W�;���� 9�)O��̻F�e�jA��6�s&fU$<��<�J�p
���oDa�EҰD鱧�Q��3��ɏ��)0y���L�Fx/�l�7�bV�<h~�ĲY¡���Ł�+Qy�eo�s(Q�+g)�φof��R��s ���F7��8�Y�g�E�γ��AX�DTX��3���A�.���=vyd�{���q?�?*8��0��/<C��e�6�k5�F۹����?�n�Er��63����Et���3%zb_T���+�p�gS��Q�%�Dz��ܬ�>�-)mK����>(�,�V��
��r�#')��ou��֙:����Q��T���ߐ������]ю����y(�}�z��Rp vH�NW�Ϊ��!mKV���7��)&\p�"+h[�}?o��GR7㚤�S&���8B*�I�|ʧ8:ڌ�*l3�a^&[���m(��A���O(�[��u�Uʋō)G-�����	*s;�ʜ�j�0B�X�L�_D��Ѩ�3�/�}sU�^��{���a &����紇� o�԰�Ω+��7}�XT�] [.��3��5�lh�l؉��X\���<MxX��	���3��.���U�ZY�Ţzݲ��+�#�{�m�J�v����bT'|Ki����J�E��{:��iE��{�|�H��"�8V��iC/�NE�{�I����gxZ4<�-�72Wj��	��fѳ!�8?®^<��{d�LW�p;��c2���C �vA���^��p�c�۹�B��6�?Pc8I��kZ���1��tf�m��T�!>=1�2�hoW5�J!�����տ����7�9�����]�e�f�z��Yp@�:�t�����|p�;V��6� �m5P8���GMy2Yї&�;؏�z!���������9_�	A՞4�s�#LHLzJ���-��l�g?9��M���`��T-�o99t�Ğ�#�UZe�C�R�.����ZT	���~z�"%x�A���|�}�H-b�J�`�JOB����0�͚v��8A6�3���:����Xn!��� m�"�,t<�s���ͻ8��"LdE�A��$Y0繇��/��,�� H�V�0�7z!AحZ�ʛ�/=��C�A�@�2����F�8<TVE�J��;Duq�~	��q#U�sF�?���G��Yz�7sMRV"Q݋������x��I3(�r�FW��R;ÎLO���?��4p�;�<n)uQ�j��dO>Q'k�禖�'��aqg�C�ۿ��¥�L��*na󥪣�+졈#��l�9)k�ٮ��w�6�C4�ȰV��6b7�k�ve"�-�te��6=����n�k���F�x�������lfv(���� �၃�&A{g��f�v��x@�ɽ��v����9��_H�S�5	��a#�C�U��q��I�3�P�H��1Ӡ��}Y)y�*��|�$�>�HZ����=e��I�Rˑ��H|9"ҒS��vF<��{ԞR��롯1����⽎b�
MiA��h!���+�y�U���	�s�p�q|��h��n�GP��ӉV�:�&���ω�KQ4T��'U��B����'�	�L=�[��3���<w�E��bC�+Y,�)�4�1PGDt��65��zҖ��`�V�����T?��č��<��AU9�T'xpfZX�K�.Ѭ+-�WbJf����c��<��}����\ס'o{-?�Q����h+�y�h�-��E�
��B/�$�UK�Im[��B�VT#�|&�G��-�U�?�Z�Ed,�H�x���r�v��%V&�Ja�o�Ol(V'����ՅF���4�Bf=���P��}�������Dp��Jjc��#_���]0����4�-֮��L6���R)���pu\�T/.���1�wg�@� �f�oѦv��ԇ%��1R:&�]�?e󜃂�0�G��v�u��wN��&2~(��k��B�q��k���x�(E�/�=Gi<;/�Җ��t��]�����]\�Y뚶����-f��CC#Y�c43��	��g��3Ն��׸O���2d����:vW�ɶ�4!�@$j�k���(6�@y��Kx���͜(���I�Ngn��)rb��6R��O�uf-�9�f�%�%������Qo�?�ܒ�8Bp�]'t`��3����j��g��%�����J�K���U��;�7W6;���7���kA+��^���Q!� (��s��Z���'�~\q�Y��%|p�}���5��>�	����9ޝ��5�xŇ��ئ�.l�H�t�!�
j¤�k�u\+�D"-?}�[�b�sx�a�-9g,����*�R�2c;TP���A0�),k�ָ�[���c��G�ų;�cvy;���va�?��G��2W ��c��K�w��eW���S�V��3��j��
p�wR��v�
�$�u+��5��/�m嗁-��I��}��u�>�@���v������lF2�B��L�M�u����V�*k�k��T�[��!R? �p�0�cbS���nVy���j���Ɉ�E)F�����s`^t������I��V�8��7з�fyش�E�y�  ��Y��a���ij����fL��k�#�k�]>I2��S<�R��D����G���?�Q�՗��(^x�'��M��k)��C�"ǂX��Lt
<KW�`�'Gc�2�<�䎾]�[������G��et��8L��ղ�L�d�� 
��0�m׭��܎�����rF�UM���R���j
v�nI��+�彋D�_�wX�FP���$!��쥩z%=`}/�G&�u�!�ǊHF],)�7�<�$��-�����wX��=W���\YU��RA�� &'���3x
��æ>8�T��3JJw�J,�|A�)�PE�1����fLJ��l��p�&���D�{�9 �rY1Wb�u�V���l�!)w<�b��)�ł��"�f�C���J�#*l��e�P��^+wk�>��V��R�q�X�1��%AK�g���0��|vN�6*{����J��$$�%��`��Mz9eo�="X��+�{�dz�0պ���g��!n�ZR�%�/�}��1欌�9i��`be�c0;u��t����|L�������L�lU������#�·�&rԹgڕ͝�˶d��ef�����/���z�vT`)�Y��p�h��À!;Ml����1t�ciq�B��Tx-��퍧j�"�n��yI\@[?�B6�����%��D������TR�����"a�x/�|Y�Ϻ �%�^��W�N���G�8�
��*��?���&o�[�	��PL�X��4���W��*:9��M����q�h��l�Yt�j�u]	<��eMp�zqs6w��*���P�D�Km�ڮ+�gJ��
��Љ0��e�&��E(c���N�7��-�7�<������c)�+B!�x��Ӭ /�����@p9�9���UWi���[�"��,�n�t:�� Dԃ��!�+sl �4���դ��fD�2W����Xה�nGQ�e�+��ks�AUI0@$;�ϡU��N� X)�1����綌��. 4q,��&��0w�9�Km�#Y'~�-4�<�/���lĔ��"�"f��R.e�t؃G��7Լ�}ęچ_K)�f�U�ڈ��g��ӶFjl��J@�<`�u�j�u��
��;�������7󏎚�I�-RN�L�i�q�WE�W����Ť;@�J��'8s�����Ϙt�՜#��>�v�@�����5M<��d�4 鬅t?O!�κ��	��r+{O*1L�����B�L�p(�k3����ݐ y@*����p9�`N��q���.���/��ʵZ7(n���}��& @�)�lQ��n�i�#m
a�ϊ�}���)s2��+Rt�j�1FHI��KW��y���n���۱���l1Ds^:������oǐx�P�<�l��Q�lkI�[ުl'oGǠd�{dn�q���<(����~P�X.^�<#�Z�Y���O��\v��"�p,:�y4���99�m�@�/���
&pdE�Aw!N��䤲=����~`�@� r>$�}�ۢ^�¡��|-�������
6���A����Z`Ϩ��Τϴ����Z��h���!���2a/�����H�tw�u�6�)��~@�~�D�[��� 捀��u3�������f�O@��
b�BD�����-EB���w[��iBz�r��vG�Xs�)z wx�IX̬c���(I'
i��E_īb��*}��{����;]d�[�0(_l�&Ć�����e�{
��>�b�	\�%����@u��%�(�f?r�_#�L2����N.i\2+_��3��<��[�z;ކ���M���;h8x
�e@�����hy�fh��ڽ��Z���DdQ�acFA��?��Qљ��O�Ɯӕ&ebF�C�7Zո�s>I�����i 8(��J"<ɘŎ�8�-�Q��*���	����pNB�B����Q| �yW## 3UF��էk:�R�N�;��ʮ��+?Bˊ@�C��l�k��fsk1���ƈ��2�v��P��B��ro;e���NVq��P��q+��G����k(0��	�n�����ӫoI_Լ-/oؕ���V��'����8%�Ԁ���J�"~���?)��M�⍚���Y����x����b�m�ė�2j]%��D!�5'�pImolzx�=����<��Ai$����ĥ�A�vӍ��ׁ�ŉu��-6�ՙ�9�U؟���To���Wz��(I��)�鈩���VP6�sb��7O,�#��2֔���:~�l9\�\�NWd)`6Ƌ�"��~���T��"V��.3�G�R�H��������j��⽤I�B��԰�'��G��3�X�E^>+��d��:�0++\̌o'�O��&�����@}6�R	��W��ءE�C}�"�`��:��5����E�y��I>`�M�ҵgI'@���e�*��\���mG�TR˟�vb�ד��[Z'�]3�c_-z�d�:���Yg�3Uw��;mWo�����C�?�:�#TVG�7�4{�;n�i]mR�8t;B���YC[�}u4���|;A��f���E�6�����ε����t�3:p3F[4�� -�\,n�L���g~;���f#Q��P/�7u�>Y�Y(M��6Q�y|��b!������WB<nT]t���V�O�]Eu�x���/��g�]~y��/�Iz$^�c�V��M��� */��q��$�󶵰~�߳N1�m}^H(e�:���s�ě����U�֘�mbo��k���o`Ʉ�Jʌjv�SF�o��4�6���_3�lz$��������!�J+�m���Jޟ}�j�w	�D��o;���N���4��r�ӹYū������[m����M��hi��ݣ>�a_�Ur��¥��c: ኩkr'��ZKxӒ��.�Z8�N.���i@�s����UR�n��n��)vn*�����&|��(�[����b�u���m_Z#�mC��scREMs�y5�J�Q���GcB����
�K3�{�e�l��__]hc���:��5�U8*�61���p��*^Y�5fl<R��7���q0j�� �sIU�u�rU����Y�2&3�� �&,��-u2���TjY4�U���Kށ	.F��V���v8�+�����w����[%i܆鯽�kX�*�c�M�-��í�tM�YÏ�	�BV�k������ݦ���!�fuə�]�3���J(������u��vE �N[�L��P{ܵ���
	�J𵨩K�\ʢ����=�Y�[/���ҁ���0V=b��,���6A$�	�A!�������|'���q?�H4��z���|���Le��Y�'���S"hw��L��w#�[YM�W��gA@�]��u4/�w��¸눰O��٦��6��}.�G"ƒ܂���L���ݸ��
��+��P;�KJ�g_PV�0��B+�K���"P�����8�ؾ�	�{�U.��p���Q��|.��^,7���3lU����� C��-�Z��H�Xt��I��Z�U�ނ��s���׺�i�����s4^>i��k�>;����[�i���v�K���rm��\��z-H(���zb���(_���/]�W1"&��\�(\��~��i��mrw�龺����).BOʏ#�/�
ǉ��&��Q���ڠ�~�DQ�Đ}q%<-�h-�?EX�����t]uB �[�!rO�p��ְ�J��H�~�e���P��c5�t�C����8�����7R8���8�Q�cU�"�:������(�q�2b�֋ӘD�X�����P��!Uj�����.�A��5a��8f�']5���-S�����Sl���f��#<ɻ�n	ڛ`���, NbO��5U�޼'9��g@dP��З��0�k7QNfxV��>z�bF��_���}����Pc�$�ט9 ���
$��w�P�.��%�f\��F���=��Q�8��e��:&""gY}�J����"���[�	TG���[�������2�Vs���LUk�Lυ�q6"Ml��9[���G�� ��h����M��� ��y��ߘ��_٫
"�^O,��@=�D+���Y�Vw�GUߑ���m&0R�!r�C��"��l���c*&�Τ&�;PP��\�~����tw�3z3$(/���%x�#�qѺj�i :�����&ȬD��Cw8ݨƫ>�Y0��A��߮n����^�{�Ӕ�)��t�^	@��P4�J��)��f)������/�\�Z2�Z����oٴ>��B6<�͞w?6�#	t|�hR� XD��k*�H�Nv�R�C�(���J�r1�	�d�R����A]A 8�Ժhۊ�}Q��~->v�U�����3.�����w�o^ךC���&n���$��S=��g	�3睉��HbU �v����7�����%[�h<u	m��Crh
z�UC�~J�Y�GX�䮽�(�+����b�5��s#��Ґ�|+������8�ھ�Ь����<����Z���_o.]�����t1��.(3+�&�c�ȥ�;��N�����s88�~<TI��U�w9�NLj�1*����M�W#:A|*S�l�Q|����@���LI�]=��X�� ��ioЬY�w�!W�,��V׾*����O��&d���`a���r�A$.?�S,����qT�ȕ�ź�8�fOp�S��bޢ��<�A2�FғM�;��P;�݊����1jv���<�ؓ��<�4-����+��Z�łtCh;�[�?>��A&0�,1���͍�$�\neh��h�S�2���Q�ySv�5�o��fId�O��#�a��׸o�.�@�� +:� x X���viL��r��+jo̚������i!I!Eoj�`J���C���ܱ�9�p���[�0���9���M�&�B9/��k[���Kz������FF��-�(吰x�G_�I�I�ˉ[�HI���E瞖��F1v@��_�?������Kf�&$�F&29u<�5�����{Vh#�p�᳭�&�Wǻڴ�G|՞{������a9�%��K�l*\q�:(�gt�����=πv��n�N)�6}���6s}\)iB��!f�,�n�`g��kEzo(�@4�r��wS�G�d]9���|_U�'�
����uz8t��[Z�*'=�J*�o�v!�_#�K��)�5@�G!Č~p����<h�E�j��3�hO���mv�=8��>u�bB9X�b
�F�}~^��͉ 3@{�&�䯆։�lˢ��Kj��4���@+�6R�4�l����s�i	`�ѝ��\��7tg��)d :.N�����2��W�V|�,g���6�����v=��6����h1&+���f3�7uT�$j�jh��yD�Y\�l�f��5�=B�V�ܰ!��,K
���yz��t�눔�e�_K� Ԁ��8��|霎-F>��1)�e�̋�p�S��%���Kw����g�e&��^4)�%��������B��]ӂ'�B@+)���͘6?�,����N��}�`K JbӼ�gG��qT��p�i}w��Ѣ�x�:��v(Ҭʁ�I��	p@[K��,�"��`����d����;*�i���bd�2����F��������d��PV�P�Ѵ��p!��õPƬ�g�u�o�xU42�T��������)�������Ȅ���dt��6Ț��������2ɝT��c�6�70���`U�P�8����:�����<Tt��� j1�x��gC�<��������"&�DŚ���
5�����9Z�7�!	���S�S��#���@�b�0�Xa� �Nub�).��s�a�1��=9��o���)S;�A�Y�u�r��������`�rǬx������{Z޽{�(Y�9]�h�y.ܴm!��?����_á('xh�A�t�}��1�Mz���&���)-��#���¶�ć�|ڽӤ�4p�8��l���n�T�����������me��o���X�FrD��v;8�Y�A��=��rmW�KM���8���C
�H���+3��m���hfY��tR�����=@�Wq�i�M5f������К��0��SZ�����$�Ѯ9�{2��_$�f�J�U�y�S<�禗ߙ$�uL��6�yG�Cձ��O�4���%0��P�o����H��ܓ:��nW��� ��9�� uk��l��S&_z`xO:�ܶ`<޼�<g�aGI���Ǚ�t��_�GMV���oO	p1��H����e�f����"��`F���C>��f�l����e؈6�@�����ܦ?ZѮ�Is3��:3AE�U�R�����A��@�yU%f��)"�̬�j��r�:t�ۂ�D4����B��B:�鉄�l7�f��S�4� ^7����A�4�c>H��u���e�V\�����;��IN�B]g���0�y��8��Q8�D��XXn��=nͭ����X��r�zO���I�H��}�%�j ��J\��HZv�)e�3X��Zhż&��?�Y�fA��5�;����Y�4��Ws�Lӛ�
���}$�C��]ш��*Lj�+S<����G�q��
�l�U�>�URy�M�j�>f%��w;W�7_ĔV�0����
�E��Z�ӎ��� ����4"�Ѿ��ÔV��)%P���^^��D�o�O�i��#�ئn����:���$@�0��S�С{V��Q��u�xCxH#����eF9�y'��@P{�lr!Po}�H2U���Hʏ_O�	��p#��S�F������Է��q��aEd�����9��m���7P�Yd��&|�[�gk/�u��q�]��8$�:n���ڌ�0�%�+�L��f�蠃�Ҧ��=~��'?����[@9�%��B �$�/��ȏ��J��$߮��@:��~jJ&�u� �o�5�4}Q�:�i�p�75ރ��T����d��S�[>Ǔa5>�����^\���}��u�	�v�.dX��q Z���bұ�_G�l&����\�\"��Z&\:�u�D�,U�����d�s˾>�b%���ӚŲ��Mq�����w|�v��Q�x:N�,��M�vȽI!���D|L?vZ<l@I%���E��"<)rV�q�v��4�T{H6��n�׈��K|���~�P�Ʀc�* $�X6/�������9҃V�-�.�rc�����6�t)}��;�y��J�\`�ǏȑO�%���a��
�7��M9;����oI�l}�]>�lt�Ʈ.����,v!]]��sB9��븟F�M���YZa�	��"j6�J[Z�ڢ<�����s���\=�!��Z�~@ �y�-� N�, J@*��"�T?�mMb�勤�	��x_��#w�y2���}����w��NF�zgֳ>mX')�����t�<g��FE�tNJ�h�w�ONz��~�D_�����tI\�&�0�ЈӘĿf��D5�b�Htvx�2�0�-Z��d�]��]JiR���}�8�I�/Q�]k@�� ��d]J�6Fi�*��Sq�m��PV6Z_���D@5�y�'�?���S�b%�.��eޙIG��:�d��y�b/Ց�hJԽ7����ǈJ� �?V %����22a!f�y߇�W��O*�5�LM��0[d Jm	��G��\;�z����b�X�{���L:���R"�YNsJH�[�Mk��OW~�6m��AF�kL5��ȧM|4�� /�WDL�\_�fꤽ-��/
�^�#QE�m��e�ۤ5D��*3�~�[d�x�_�'���'AۮTFs������z��h�<+ԧ�1	�~r�s�p�h�f}7>ԭ���:+Vn�9�"�� �(��R�Rű욯��{.�Ǩ��&�XA�`��à5"e�����خ�Yz���ՠ�!!ӻ�gӘE��هg}m.�=c���I��֎{%> 5�ۆ[���a�}��Y��^2,&UE% X@
	19O��x���g٬\{�ΰ���#�h%�)[�S�<d��=�NdBe0D�ʘ�z��N2�8�6��>�L=���򓚞�"�$*ÿ
~��ev�N��T?&��3)��],t���T��(��B�N��w����}�&kTU���!>��>;S:���1��s���������NE� sM��:���;#����:f%]z�]�H������Jw�o����������ʇAm���!��Fq��N�n��$�y����L�`@��AL�Ar3�$�253�f�p�����ہ�����UD�GK^0'\ �����ړZ�x )��hW�� :�Ӎ����G�W�r�-A[p�6#���<���߃�|��2��\Y�Qݑ_�O`eu �{{�U�f��ն
�#�D����/��KHj����r0Z�G�rhU6pHK���^e6��N�~�=�ks��y2���W�U֎?M��N��]~�7����m^}zD��02�Ӱ��r��8��W��[93�=���7f�s���Q�(�7jvG����:*���L@�[O��;�B�/�[@�f�s���J��=f�m��y��W{��y��c_!��@}_��Y��@ѽF�<�軉5���lN Y���b3쓝���S�7ɝg��]�B�nX��15����?r?����H�]��+H�y|$�����&$~��=T�m��%��tj��0u��T������Lv��9i3b�!�C�kR��RHՉv4C�^S��WeĐeg�#ã�����J�Z�PbѲ)��էN>e��o�z��Y��q2
�0˄2�~�l�H�������T-E��i�f��
@�ׂ���M�Mn�F|)�TP�%4�4��
M�
0��s{
��������\Q�Q�Aa���%v��}���@�Z����z@�������С��~�o�+����;����~-��U�p8�F[�u�;��RY?��w�-��7ɳuTr�] 6��;B
���n�5׽�qG�e*�4H�������L7Ŏ��[E'�Y��x��W5���r�6��[�󃭷���m�a1��1�n��.l��/�n���,`J�j8m�X<�W���z#�ȑ.�3���6��IR��~X_$f�%u�[E��>s}-e�?mm�'p*����	�C��n�ss�yD�3k�"'v��#6�������g���pu�C̹>CF�5]!�)C�c��������a���|�&���g�
m�ZI��܏��(��y6���iV���KO���]t����<���emj���' ���V��Ilt��p��=-9�j#�p��/TF��1Ǉ�ݾ��AI�>6�c��Ũ6>Bd|"��2z�����h(��]Zu�Li�w�*�����z�5��B�
j2����&�_���7�s����U\����:/2|���
%�>�����y^������-�{��(�kQ���y'��yvo��9@"� ���y�O�k�
�yx�g�4�m���y���`��Ѝ$�� �,��P�}F$���fE֐��1���~vnj�Kט���ac�e�P�{!�E-��i��(��p4"�I������%��Q3hiS]Jj4L���m�WC]q�ϭt��8^�c��K��pw��-��L ��u��=z��ǚ{#&����W����V4�-u��S;��a�{��lء)��&��{��va��j0�vKFH�V���f��ً��Wz������y�������`�U�u3�����I�K�+��J��/���T&�0 �t׆mV�(#�3��hr-:��U�{��x/��g���$��m�
E.Sd��|���}�K�	�~/λ�ry%$ST����V`��El� ]2-��K�x���̈́�4��^H�7V����6��h��pi9p�B��%�J��\N�y|nCB� ����~pbܙ���}__����������#aݠ��Er*�JR���,;�euK�����Of�I5P�)q�=��&�9��/��&D�a�s?��D�xi��^��?5��h����1E��e���0���"]A��YOtP�߇ř���b�k �K,�M����#sFkN�i����=�'��m�bD[n�w_���mܬ�,LHXͱ%����3���rņk�c�ִ��7����e:�j�SI�:�Y
�%s�H��u��8F��������zx���L�1�KE��,e�j��3���Szs�p�p$����߷��[n�&��ܻל��a�7��LFF�N���U���R)�N��JH���V�#SYQ��6ܨOo�R����i���� ��/o�V	��v�B���`��t�W�!"�sw%�p��6T�M#xv
Ni�jz*�^�����C[�ȰYo'�"�;7QC��9��[	f'��#��+�ϑ�vC���.����Z�g�#�� i��D�����2�*�U�|���8�`�|�����l�}�m���N�gމ(�/E����5�0����T�l�6����&���GF�4��b}�� �a�&����B��N՚%��Fd��d.Z����l?���{�����x��/ʻ;_L�WF׫���Y�S�K��|��'�l*k�=�x�ȰUD��:�f�e���j.ڹn�X�%?@��:*��t������7�����II��[��ى�����s�>}���S ��<�Ж�A�lJ�u���D�|�B�H:�~��|���[���yz?�t��>\{�Rq�F��^2LU��Q�Z�H�o���pS�V�����Ķ�h�Z�	�潎���ZdY:7�O�mP�6O&Y�Ø��@܌BD�ǟ���Gj��j�]��ee{C&�:�f������ϭ��W]@��|rR P�u&�������7���o��ō��D��S�%�C��L���|E�w:(�d#Cҡl����V�r(]r%i��fȉe.�4nP[�uH�;2���*�ĳ�U�9!6^���e���.G/�	��g-�=a����m�D5�p�u��|��L��m�8�f�b������=R���F/�h��T*��>��%�,4�d>�J�iE��]�M���ru�
8��(��K�W:+�nrq��C�xoo�W(N@O>$�G9��dA���UY~
����;x���*l �͕��S���ĉmCl���@u�Fb����*�c�06����(/go�jQ�7���:k�*��Tz�_)���c �;%��������J�7��s�q,N�^�v+�rg�}��Aږ���{�?K��"�*a�GN����f����B��	���[5 :}>Χ��Zb���|�U� ����L��%
�������'�"���rP��h�X+��j-��-���rN�B�1ҺK����3�f8�3u������<ʛpIܼ�Hދ�@֤�K��l`؛׶0K�q�����[2�q����Yw�<_�yΩ��q>Z�{'D���%�ʳ�>I����fFz������w!30g��甬�����,�w`�3�1Xul=4O���YS@+_��<�b�N�; T�8�����U�!A�5wlى^���SІ "?/~U$���t;�g�z�J�3����F�=��}a� �3~��՝]L�ղ��|h�0����t�S�82�u/"	�P�Le�����Z9u�����,��d5����	��O���&�Ή"�/����u
����5I���^����6�{+jQb���R��PQ*�d�g�*ܺ ��n� �����N�a�1�Ĺ��z��4�az9�G���tR����!F�8th�~��P�{�{��M�#�~�yX7k��t�BL���2�-��4'1�&���p�竺�jQP�V~��|
��*2#?�F�)���Ui��G�u8~9�v'��4���zH��:�b�ώ���e��o����)�X ��f^�9��<��HK@t��>�zքw�����x�~�[+������d���6Ϫ�@M�
�)�"~�*=G�	���,)����u �Ys�?t�=N����&�C��S�v�Pr�-var�E.�K�"��D+5D����!���j8���C�"`��zz�}:_��A�CBܔ�������	I@5@ j�*�����i%0÷a���P̼���%(�Q���Y�`�D�<��D%�n����yq�h͍3r�J���R��e��T��ԓ�T��U��Oj'i7�w�~��"��B�BvQ�Z��St_��x��ڵ񍤗dP��R3Ñ�J�2�Ut�X 6�M& tk�<3qO �l�9�$�M�I4)���3��H#�=+����3e~"y��p�Y�����K�^�"@�=�����+�?��C�wP~��qԤJMpzr�%��u8"b��ױ%��y�o���v*�t~�����Cgy��y22hfo���6���ƛA6��@����>��1�A�,���蛝��3���a\��l��&�͔i9�>o`\����J�Р�!E3��ڤ{5�z��OS�?�i,��`Wj�Ǜ���P:��mD����ː�ל�S���_W�J!P�~�bMb�5{%�m��:f9�2�����H�|S������ ��[FOJG+���_BNR}XBZ��e�Ǐ��{c����@�۔�\��o�h�`� t^̯su[)S%urx�� �x��D�fז���Q f��(���6�nGȑ���x���E^jN	�D+�]v��
}M�UB�=cX$��E$z�y�7�/˯|�k�|lr�Jי6(9C��'��)��My|�!�j�>S������*�i�����Suf���Ա ?K`Sc5g�[�`=��)�o���)�9����1�P��k�Qc�	�hl%��H��� ���;����P��*N�򫠱��ㅪG�|m��כA�����{lFN�__�����L�p���,P�196l����<����ї�5Y��$3E��ZCr�d���za�� ɟ3��2�PxV$�=63y�梢?�2sl�J��U���㳾�REMo̳dc��8�/Q#�������r^g_� ����aS��>�U���~I݀X��8^(��KQ�kv�a�ʬ,"��4FV׬��HL�S0�i�V��$���*���f�8���NʾA��|���
/f׬Y��D���1{_���)L�@��fnv?4����7L0����;�	�$�<�i���!����/��2W˩0u]VJ�i��SLXKʙ���$#Jd�3:���c䐵'��,M��tg)"::9���r�ӔTC�is�"�5}���1�q�#ioLܙ�ybY�����m���m�.p�1�>1]�|r��\P�>	�0r�ߑ̖�[�S^�4��e�g=� �ƦU䢨$?!��W�_�y�FћA1�c����O���oJF��^�|nŭR~�䇳u=Z}reB��0}�B�q;���PLr��^���~�E��h^��a m�{��!�����,3�/���J�~���"�d�OsA�^�c����h"Q�N�"�93��4x��P�c�u"�a��:�^<��h0�p���G�u�/w\.�Ǆ�s�LC�3~X&����V�¹���m�?5�i��hi�G��J֗]���5�{ѧ��H$dW�~�S����K�E����(Ij ��i�e���_a7���7�uTWk� � �,6{z���:gy3�k�|r���� ]�ql���7�v\{��
[Ԕ��U�����6�����t����RbpV̫�Xgh
��M �i����)�6L!��O���qR�J*������I	�0����-jf�ax �!fi�F��k4�צ��A�d��е�� �������%X1&+ �����k���gԭ5Ro�g1��Ŕ1��Ȏ#FVE.:-���n����6�|t�4O��;E0�I��0S�i����=�T��"��o^!E�����*���D}8hZ�c�$��;7(�G�W}ޙ�����AK3)kgD�p��b������s/�b��[�K��&\Gt'�_��/���y���Ƣ]Ĳ�E �#�]
�>�iC������>�O[ސ4�v:a��L���ҹ/q��t��u�4�|�l?���h�_� F�h%r�� ӂ���@c5� ��g�8u���@��s�z߶��sq� I��sSn�y7�����Z����E?L@7���/���[�{�,�����#-��㬐#V�Ѕ��&�	�$�FƵԀ����I|�涤 㓠��ы����:�Ο����j<90�$h���U��z$��,�՘�
�o��s�ױzZw����p^� D�$,$4�L���w��N.P�M����Y�@�M�ǔa�%��	֙�${v��)n!�o't���rY�iF&6{'�PZouZĽ��wh�Qt Kb�s�mR��v�s	�zX�=$Q��29��Ux6�t�=�A��t�V6�5�q~y{���,+�XD��K�V��b S8�0�!�*޴���o]F�N/AiI��Mu7No0��K�"�d�{�Ϥ�d(�v�D_�Ҏz�x�����*H�d�]��f ���A�hdX{Z��k�'���G��J����2p���M�������\ǘ�1� �W�4y��'g�� 6����umH�cS�{��X�M����>En���:;�8(:�J+e��}xUD��=ª�'�m�MRځ1�'��������=��?A!(��/`�g$�5�Vf��!JB��qH��\1�]�˩>s�uݖ��B�
��c���b�z�}�BC�m��Cّ�e��*���E0dk�;s���h�6��>#6��!���_�o�@e#���K��a��)�ƭ����@?~l]bhE���ؐ����wVK��B��V�1����^(<����;C��U��į�h�;�]f7&�]�#���z��s�$G���ou80���� Z�Y�EO�����*�`._�)3�^�}�qQ ��FH$Xo�;��|a���P�@��N����V�;Í�0圙B�dh�� ���q�H�_$t��+}f>�d�6v8R�.�1nl���4��%U^�����. �j.�� ?G����5�W�l��K��m��V$o������U���V;	,�����KЫ�D����j���q�w��*����d��Jߣ@e�����QZQ���
`3���������(NJO���Nr8�|�����*��H�S�з�>D��1٦w��TY� �Wo|�톯#��f14㢽�I"7xkj]�S�9h�j��0J7-)���h��{匡PJ�XO��<�j����3}�^J!��0��+o�+�e4����k4��C�$���'��9=���jv=��0�g�AP!"��d/�c����WH�DV�=Sx2�l��Q�ז
��/e��4M,/��,�P�e#ח
&HSm�Xҋϱ�8�D1,ߡ�I�q�;������~{7,%o��	⁀��Ɓ���������2
;�9%�D��]UfK�Z�}��G��v����0+d�h'�}L��\�%e��[:ܫ���;�u:�Tb��]��bx���ҝ��S)�tX�'<�)�4�"�-���O�]�T6'ld�\�i"��MHa�j	*��o�]����v6���#|��M�G���L��:��V�\M���zT6��3�$�]'g���w��$�4��94�V͈4��Al%�9�|TT���,�`��� �]���2 �!a��eR����F�����NH�7? �#�|o:�i�  ~�E����d}N���VX�S̈́N��8���X6�_��Нr̆s�2d�2÷�'���{v�͎����D���Q�I�T���ku��L-T��*FЍw��t�E$�gXl>y����@P�^��%M�p��%����f>���`%�v=��$՛��]�6g���a�M�h��B�� ��рMV�����|(���ܮ@��ò^��6I��˞���,�g`(�ұ�������.��F3l��*���(%h$���H{W���UQ���mY��K��u`֋���y���e��N�u߄��q���'�O3;��G\��'p�̤*9��8��z�_F�����a
T�$���U�a��� 3e{bX�))��e$���H��IdL�n�p���!s.�q4K���V-�m����1�B���)����#c�fSyiI��;h*��o�#AJ���'�O�J0t����,Zr'4f���w�M�O��rtv��nT�*O��$� 6�m�74���2���G&���21~�"Չ�����õx�@8�M`
�,�<�0<��X���f�2��	��r��%�FΞ��D���b{�]f��ę3klTV�g	��`/�{0A�<��(题���?����o����#n�ȫR� 14΂G��bj\b�\�����W(6?F�%�9�HI�����E��>����:^�B�X,W(`�X�Æ���������g�`��6�c�_e�k�POĪ��"� .�n˾)?�����BL���Z�����wA�nX�[����N�r �ֽ���z�KxDq;���`\�j��z���b^�"�͸d�[�,d
$�׉��_Yk��#�#y��6
��f���
��
W��N������^\�.Vy
u���=�2戝D"���L����M�
�X�z�YС������q�H/y�l��^(��[�ˬ�&G����?3�c{a���	o�j*��������1�xU��\���3���h;U��_�`߭���MUR�ޤ2��C��i�����P��]$7���Pcɂ�)�:��RF�He
)V��	�i�H�/�LIt���WAe�M�`�).�u�/4��vAffI8]Vs6�����HG��A7='�I=�NHe��$clpa��-dؤ$U/e����	M̫b�2��[����gZ�`�X����[����廕�S�*����x�g�i�[W<�N|�����e}x~��/�rx�yH�a�ܲwB��+��[ `������?�B��rAv�#��}.h��5�z�KW5ú>�~㸎���V^��1��0�"���L	F7�X�G�����3�2�������6Xe�!Z�YM��{�Bhʄq�MJ���i.���
���v����I���F�+�����9�	C\�jnNu���u�
��N���fV��]��0fg\)�-;��}/�2��;kFSpO��NW�'����>�5���Ȩ�F�IE M����͚o�o>���&l�!���(<g�w��M�$$}D�a~$Xȴ�_^���<�$�����m74V;�Tb�
�������E���n����8r��7���@a6H�����}Y"�z�D$q�Zu��B憵���Дz���ˀ��;�4���o�#u����]s���)��^Ѕ%�PՐ��(5��D�T�4g�~�����j��sDtP=$��CX��Y/v�KN-�/� K%��Y�)FO�I7/V�=@c�9�
C$O� ����Ž ��!)�	��w�w.�L@x�iz�����"�i�/B���Cz>͗/�3OZDV�C�Qx@'} !�*��a�]m_pؼ��
����<��ĩL���+�2����� �8��Q=Y�Z�k�rR~��̫ai M��oh����4I���s��I7� }rjO,)�WQ1G�YL^�LЏW���W����_C��YI&Y`!�2$���E��,�
¾Y�],�}�M,���<��Q�^�w�Gw������ũW��`_�N^JԊ<t|<QYq����E)8�8_���_��S�\>�;oH�;
��FWw3y����ϙ��f/&.}��vO:&��E|~�V@�O��`vS��鬰s*��m0�B.���
E�ܺ���p/���7�$��Ϋ*#�&�D�2�-t_��������<�n�w�b�Ȇ�DȺ���U��i��+
�åG ' ;�d����#c����;��V2��M�R[P��� �������D���� �P���B�|ti�Oп��������K����]R��s};K�x���.���+�#�U�Y[M�������rx2�zeXo�e��*�Yy�ӗ"Q�ykB$���2�$k�h�v�>>H 3��{:�.��%�^z_�7��v�;}{u�|vG��ȫx�'Čݥ| H��Ȃ� �f�(ԁ�����?Z����M2"���W�,�FRP�l��������}>C�|;=��	u���/]Q��W�K�
�ݚc�}h,��Mt���
���vX�����m&��aE�q]Ş&_Ǟ�����a�Q��K_�F3���&E�S�J��ك&\�k�L� ��i4����XU��f��4�)��Q!���,U�|o-Y7�0�F���dP�7�سPl3V�,����ׁ�zC�Mo��]�p'�ԙ<�B<��dC�Z�ڗRS�(o���Teϐˍ#�X�2���f29n�s��'�����?u�Ͼ�X��\J�v$9Y0n�-��&���N��̉���=��)�i�w��2�l�1��:�gk�ybVAu�W�ˮ��R)�ڻ��rmI� bO?�w���ءZ�X��mWYd������PA��s��W�ܳPɺm�w�^������(��E��?�z��6[˂�+��*�8=��Z�נ:͚� �Z���&
N���U��R���?��K6�2z��w>X�p��^).��x=�BA�̣��;�A�r�=U_���y��a�ӋDyZ�aD�@����v[K;��'�)�4#�.�c��b�$#%�}�QU�������sҦǜ(�e�8��U%�,�s��y�u<�����y0�P���"���Xז���}dB�B��:�CO&n�r%0�y5qh��NA�찶���+j���
�$̓�_���f3/�Ң�{��g䠴�)t���(o[s��a���D�6�#��`�5�t������Y	d��)��i��EF��T��A�?T���
�Ў|�A�L춰@H1P��'�h���#p{i�c
�(8أ����`�##p�T�{3����8��О��EN�=_	�:֦�Hǔ���i��N6��W�1�}N�[a�X�z���1y�{'9�܅��o*�6�Y���V?ml�Q
'@9��;����L�N@��?�9�,�"���39IK����t�h�.���OU�T�[Z�;�������w{ ��xn���Y[����`H	��^�-��x6���N(���]H�,�MZG��xSd�E8�9/����C�m0��
�2[�c2jiQ��ݛ79EO��lg��TJ�̫ȃ��_��Tw~���������m�&6�S�*A�l��P���F	����E���q���ɉX(+�F���p�ir<̭�y_ĨK�&?VT)�1L�ƽ<��hJ�\���!�$Ѣ�z��f`JU%�k$���&疬z���2i���2%��ܜ�>Z�`sk���n�b��B�+�t��n�1@hJm ������)��U��Ѡ���pO��1�_�Y�]�^i{7��B# T�7��5���0��`��+_9uT~ʨ��{Ћ���R�]��o�Nl,��$@��+���~/ ��b�w����P�lo���:����i�ES�t���l��B[�<�~]tP`��Ԕ�T��t��\˕Z+�T��M`>	0�
T�[%�	�TF�g����󎭵��C�+���FBqzs�Q��o�o�uT�*�-�L<{lص�00��A$��ܯ@��~��He��}�w�g$���ǈ�E�8L��Ǜ
&�����><��{�F3�|�jP���ۉ�fA�:@�V����i�h7hWL�ai��1�$���T���Ӆ������cӷV(����O�\��6����A�tA�����/>�����y��������G�w���}/u��fd"��Z�.���f\=V_i4�-b�"����[0$�-ca�fX�"���3�"Rem��Ͻ(���&��3�hOa.ȞO�����`	�M5Y2��h4�1�jj㩆T�Uy���v��E���
9ߟ���;�Z"�8D�b�8 �2�ţ@l���hC�zRq �FZ=���#vU���6�{�-�h�p�������gѧ�E��P8����m|&����ׂ�R�"�XZ��`� jwFU�"&1x�G�h�^Y��vxn]� ~��[�N�Öc�*�OX������Go��kk1�¶ʪ�ZiMB��a'�������#���'8�Y��`�m3r�$Sḋqq��j�$J��}�����[���Iu^��=V<��4Bn�2��"Ӗ�l�4�9	�ʇ+��ѭH���F�-�[��SxS��Ź�#'OW=��	I���/�Kk򔇳���z�D���qpn!i$w���\&��X�nu|&E)����]��T���#w�BP����.�m�����mQ�Ts�S�vj9rM�=P�Ը�C�T$;k��,Ǿ���d��{q���
���y:H�&��D�T�{EaO�Dkł����l�{S휛V��A�5�����-�"}ʲ�l�DRZ�щ/�_���ei�*Ej�u
[2,�-<��g�E�y.���/�jWi'�k��ik4a�w|@�I5'��z�x���N����v/� !�S���:ٮ�H0Ւ2����8N�����J H,u�Bt��x>k�F�d7�[i6(�jݕ��lΕI���n��L�������4<A~�T����f� yj��-
!�C]��i��*a-�Q���f{c���g.�>(Qn'0Nc(ƺA�&w��r�d��˅�:v/��~��p	�Ԉ�������: �Sл����ܱ~��t&���M	�%��}^���Zl��=Ũ�4����R|�=��,ć��N6��)�Pd�oh�Ѷ�P��;ɫ�s��ĳv��`|!fES+\��oə����jȚpꧣ�y�����T���v����y����@��Ӄp ��QΣ����rɨ�f��ݑkg��U2*E���*���HN�&��D��c�C�e��~+�z4��8U�C�b��E�{H�|��V@B��I�:��G����A2]rЮ��Ul��:��;X����  g�:��ج���!	�R��զ+�(,���C�t�F�h�j]ƴ-�^��w~�Iԗ
1n{9��c��^&�Ĺe�M�L����j��I�C�IQ��yHI��i,�Q�ƜșV����l�ͩR��2�T2��U�/�.H�P:��9ٳeU���e�	�4��:�
���	ό�N'��|gk���~XCН�&S���&�Z�W�]�d���I�Nb��[9��P�����zA�O�@���,�;^]3f���~���N>E#��+M�m�8I���q�v�!
w<� �BV�ۃ}�-��d�8�+�4��{�������3ZԩtY˧/�o�P��@[Eme^�r	b&R�[y����?����]�X�!�d�{G��湾�ZZ�|�<uϷ�8|M)�z�{���3���^���H�줄��~�����P0b�VTP�����e
�6��"�ǹ�:z��P��E!� �/�%"$�����3Lś�y>�H���sm�q��\I�S1�� =�T�d���m�!��൭��8����=V��f(��o��kIT�Д�4�%��}��VɡsK�[_\�cvs����-�{���P�Z�J��cߐ$�^Z���b�8�>�W��F|�<{�C�Ɩ��V�1{�G*�S�5�N\�7pD !��R?�U�����
����;)���[�5�.���i'��yA8�`�߲1R�UєX�Θ�F�h�ן��B�,����j��ܨ�~�g�5�h����J���G¼	��pև�y��\�t��)I����{)�����H0�~�c0��[(wl��0�,޼>�¬KV������"��G�}�q.�����DN�LD�,*�"5K���y:�ő�����	�G3��(�0x�'UcAt
� �����|g�� $�`�s��k�\c�ŀK�y(�1�W�wi����Zp𕯑v6A"���G��N�>�.cP�����$*����Uv0*Kۡ���Hn�H4I����XSW\�������&R�{�U!=ӭ��#�ە�"��f���n� i
eX����i�/�hn���@f�*�wet��i�<��=��gx��霤�7F%Z�������1,6�ݮ���Q�T��G�ރP�d���@��{1�������V��~xx�4�$��u=�Ý�(���qu&p�E�*2�?OX�6��9{�N+/�Ј�J�'KR'�'Y}�^S�S�q���F�-��=kPmR�.Fc*��*y�#v=7S�t�i5�d����2�������~i���������*T����(.�u��ݨ޻�?'��'2��p¯Od�(�AtE4���&�#�ɛuq?fG�#� ��E���{�.(��.(�ƭV�~��w)bw�.v�e�����d/�z/k�f��Y.�Cyｖ
ѥ)� k����#�l��T�x�KS�:;��v�%�H?���#J�;�6��N��	��L�6Q��t�cK:�a�'QP��OC�"�o*��e	-�ނ�1)t��n�X��Ϙ70�����������-�&�^�� ��Z����uv!}厢�Z�)0�\�y/2�3tc�"����VH�+tf2�/�7�l�p��3)�{�<˧-�-�<��dg�0NC�a�o!��=谁��k}���;��F �9�W.'l�jO��.�}�*Ho�g�3�}���L���'_}�.m�0�^���c-&�7O�,�ـ�_֪��X��J'Io�xsR�p��_�L������s�f�������$��z�rR�ք�����t�T����x�'�0�/ς����KOX��A䬜��dB�-w�'�	�*�`�+J˭Ikǧ�K�J�<�Qi��bn�2ԟ�!#�@B6�~t��<�:{"�B�q�k.��fv,
�W P��Q�懏��Hk�����SMv!㽮*��f��t�̑\�u<n'b������ݘ�'����$��VؙF�+KTa�z8�=�����L�T,�.��-����������ւ������7��(N�)_4-�#���(��Cc�2;�"��;
���߫G����a|�pEB�%qGZ����˾�㪉�Y^�8�M��d�ؑ�K+߷� `٬������>E������4�x�Q�^��������&$W3���+O��?n=�srJ��}'�F+���!cw��q>�������jyԓ��EO���5 OME@&�ߛ������|K�mf΂���6���qB�r��N�ͭr��\�o$�(	��C����ո�T�u�0eC�
�� ��G!s����aaN��s���I�̈́
OfJߍ�d�5Kϡ��}xAY>ܠ=�mz�,g����3��ZԐ�KȕcC
�$����N����{�:�;����	N;A�a���vo<�S��Z�+r?iLC=�Y�n��Q��uP�-T���qV-����������/M;�kK�p���-��R=y2�E�v��E ��*?.�3��m�.�WNE#"�f�秺���1�۬�4g$͚v�� �m.7��ی�I�&T�ɜ�;����qG�G�BŲe���C$�nַ���E�6hR�*���h�jN�Iv,�����JF�6�����ݯ�� nơ]?t��¢���gF�M|�Hh
��a�S$9��/�����r��/A�Fqĵ?�����Gh�W٣'!��熯sA�Q�%uJK)[�>#�����<q��YR��Up��ލ�c�2�"2z4pH���0,���u��"�n���nw`/{�l�UDin�n��c�*�A�d��
@������;��5�K��+�u�.D�;i��%N�Mx���]�kT�e��xLRt6~u�m�#�	���1@�ް��U���� u篇���ve��.�gb��_Z�6��v��~j 3��0��%��o�E#�����P����Afr�-VQ1�i
[�RLP�|5��
���S�x���S��C	�lI��R9P��Q���Î��V�i3���S:,wb������ނ. < '>��4�5���ξ#S���I�u�`W`o�cj!���/�9
�єq�+)�蘨@��*�[��|:���򾊋�������r�6C�h6f�N�y�NV����D�1k�CBu��JEޙ�}ڀ�l𼃏Y]��^��^c� ^]��y���ŨBe�2�s�l�8�L�Z�E�P!�!�UO�ۑd�,`�1�0<q��2[:-j=^�$?h
�^oTg(�yn�r� &�N���JSԸl�����Gq�q�V���	�=Ko����7^0�yV�ig�wL)�:����uS�R8��&gg�sG�C��󜖥#^�$O�LZX�WlƤ(o��J�X�ҩ(*sZ�mfk�n���0�X)Hc��$Y���9�f�#�EC8L�Y:�l �N)<���*�S�J��}t(�NQ�Wr��~ٗ��{���p|����n�u'e���D ��E�>Q�"��Z8l%!��Q(�!�b��L{����H������	�Eb��D���� N�`�Ph�����t����q��x��z,A,4��F�R��;��)"ݯ�hl���L�yÕQB)�.�'�.�c2��G���a��U��1�f��V��{lu�1�a7��K��x�D��܁5���Տ97t��2/�K�NJ>^���s�]�ޗx��F
�&�ѣ�C�$1�bn�2p�1���OrA?1���G:Q��!@fե9�+���Ԋj
��]B�y;X�Q�%YTo/33�� �* ���y��T��U��2���lBLי�KaϑT�;�`&c�o�D�Y�<�q�I�E}����]����xd\�X��>9mng�q�{pk�Q=Db�(V:��DmY^�C�j�U���#�D|LY.��q��R��ܖyW�g�A,�s��xg�=t��Yl?F��"�p�opq�S����Wd��U���]�,~���-�x����&N�%6v�R.QUDԭ���uu����b6����eg����+7�$٧*|W�`��y�|��32�t{^7 1����nxspz����fS���9�����}���9?�h�=��e����������;\����D��an�[5!�X�����예G>�!2���,�UF�km~���Z:���P�@��u�|}��ܶ�]��y�tU�t���0���Q{]B�sܳ����=�����+y�kM�2��o����u�3�<��%|������oUf`�k�jtbxE���Z`�z���_ӎ�;|9�5U9K{�d;��L�HC
b>W1��	����[�OM�a	��%N;ո�Ɨ��_cB�m7yEZ������`٘���#��Jʿ����g�������1��[ �r��&��.l��c�.@kz/ҹ��T3`f�λ#ȹ�9O�*��B>�g�����v$���7�z��B���hx�֠�2n���Rw�����g�v�p$�&!�y"@2�/01S��P�loR��Z#G �_{��K6WykvC��ȑ-��h1����(WM1j�QU��4	7d!����,��HTM%p7�f�xNgj�
c��|�����
Ɨ�qp��at�/��o�w뿾��@Wei�cp�hE3T����7u����KR�y����F�>JA����_�E��A�w���a��%�������g�9��i�|s��L��YQӇ�8��ܤ�Rj�C��%�+a�^uɲ=^���)�����f]to�qX����H}z��=9��PxH$�����xl|�4}���2݁�Y��ۿ�c��G��vrb�)��屉J��uɿ��,"i�UG/;�nѺO��ܶ�/��ø�ǖ�4Kp��l��!����?N�}
/ѕ��E��z�vh=@KCPԿ��jhW��&lkRD�
Sf��S4pEI�����]c��R�(%彔 �.���~����5���6�\D�@Ys��,vO?�!��x����j4��}���z�G�R͗�k"���"��1�̽��I�(O��p��5P��������m�r�m�*��t�8,O�l��U��&�����L�<���=h��+!q�Ca�4}�z���Uh��Վ�KA$���uh�Rw��Vd�����g��m B��Ci�V��N���㖥���t�|ٍ���r��E$���Y�\P�\!N}�ݔz�U�:�#̈����jN�Ѐ�˚l��ɧ}�nn�zm��`��ח�g�-q ~x"������_w���L^V��a�y����fC�r���8��G#�9��@Щ��M����u� �����R�eᒚ����T �/i���è�G��
�V+-�Ny&\_yز^8N��;r�+���
��$h�'?P�:���R̜��a��v��c�F������nG�?��Ç�0=YX�*�&�6tNi�(��u��9{c���l��Ğ���}8bI��]I@e0��}�~4j�n�w�(�[�z�X��2O´ff��5�Z���^�gT��UU#�V��&j� ˺11������*�]G���:�I�D|b���ٸ�/hH�za<��n�����������Hz���I)[���!�#�O���А����A~��ʸ"R^$�Vq#�jU2k�v\�$pd��lb�)V9�_B�̫�E�r_G� E���*������6����!S i���!���������n���Q9M���B���	q��[%ƍe}���3�Xk�e�-A'Ƿ|^�eÇp��y�܎��% ��P�R|���������ILM^Z�h��(�����P.��-������D<C03A������1��|�(s`�nHm�M(��V�@Kzk��+F����piL8���f����g��O���F���xL`-��^�l�d� �vYDj�ݼ�"��>ٳ���I�Xʗ����z�#�h���?���S:v(���^���u�c!ӭ��P!.f���7
�a�[+�����yP��?��?�J��������M�])�1���@]�;���Va�< ���OU�.3���x����������P������~�P��1��R�Q���v����EB'��K����h{[>�t��'[Y��Db]�0X�j���*�P�2�.*���"X"����.�_/�-�ZfMVr=\$$<��W��y�>0�_w��6�i�^����u�k/��}�������5P��>x�#*�i�q։K��uqY��'p"yN�!�^�Ӱw�G�q�V-�r7���g�묂z�Q���|lsy�FHt4��H�N��b�����u>�ZE���F.UKVl�ѳ���kl�иf�@�'���m���0(vW�>����V���m�H���������I3��I���2S���-	~e�N1uI'T����PJ)��g�N0���V4N��X' �o��>�|�\���@�=�C�9�hv[�K&F-�A�rH����?�EU�W-��o<nʑ˄�M�$B�&��ݍg*�%�Xw�E�̇��­Y1<ݟZ��G��U��[嶡q
��$��{�~IҪ�D�-�Wd+ɞ.��i�(�5��J��!k�P>�[���.{Y�'B7�O~�i���C\���CR 0u�h��ݪ��t�v~c*m��|Z,42'�)�(�C͎Ҫ����O~���?�a1�����D�r.*�����Td�}���n�y�7n��$2��sӍI�+��`�v'pʢo�S��G/�y|�����k�z�7�
��p���d̼��s�����g~s�߰����G:�(g��|��CR��r�[����)�1��ؒ� h17������L��v/O�0�ۿ��u��.P�n�[�S<��JI�A�����Bi�b���#��c�y������iT����� ��
/��R	�K�J�@�Ԁ����a�~	�j
�3x�Q�i�C�QS�Ss*�{�_+�Y����	��bZ���a����x�T=5'Ӵ��
{WW�J �E�l��~EJ�A{8u�f@㏬�nĴ��YO	�P�y
(��eM�ホ����n�}O9�/���/�͂>8p�z���"�;��6����T�Eg7<�4m�La���4�MQ�|l���f�-%�Yds�k��7���w�e)��lW���|@�����5Jři�Q�i���NI�_K�ۀte�����W�r9+ߡ�I�)��G|e�o�*�>��"Ca$O���R��13�%]D�+7�!j1�=6>�s>�?_[1E����YkS[/I�Q�1e��Ow���V�g�sD���}&�>Y�r�B�/��u�N���sT�z>iw�@��~,�K��.��@Z8��"��[T�
�p���/*ꥷ3���f�����9h�Ê����Vr�n��ѕ��*s���|�\wq-�`Ds���E�V�c
G��%S�W���.�`E*zBm���^�WU�I��2̃Br�(�f�9��kn�=�y�ѷ�Z% <g�*�6&��`��<�^����S��c��0>�ԁ4��< 7�(���vPjN;�/m:�5�̦yx����%f>���Y��DFɺxK�!j{��-Fտt۟	�q6ou��*�*��ujH