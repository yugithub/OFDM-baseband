��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ^c���7�oR����|=L�x/��)�.�H<^~|n���=�I�O�f"�|Ӭ#���L���"�/!<O��Q�SŁ�@��V��`�#�UXJ�>���2�B�d�R�$w�����ˀ���	���ga�h6x�.��{<��]�ߓ�Y��K?)�������+��;�D\�_A���s�nSU)c7[�����k榥 ���7G�jأAL�*�Zl�.�(�(:$���+wa�"�Y�r�1Ǜ�~�m'IX0"�I�� ������3�_�N�6��J%FSl xr�^d�,8����Y<NN����[R/U�._/x�$p��������'����9��f��I@#�	Q���E�{���	�m`�=��W�3%��d�p ���_=�R�?�*�sM%�iJ��4i�<U�č�%�v"��R��\��9�*<��i\:dF���5PJo���˹���������=;�>?V����x�6b��l�%5b,kS3&��K�εò�PG��c�k��ld��Ni�d����5�c��}x?�Tә���#p�GQ��+ՏxR��G��Y�@��=����=��z�a��xlAib�#x(��eA����i�W5�o����]Y,�LUM��#�,��O��/�:�f���P��?�#��~��H���Q/�M�S��JHAL�nQ�,�)�s{C��
�w��t�u}��A��w���=��p�H��"�܌�� ���1�l�#:�����}V	�4A"<CE�~�T8�-�tj�$���-Ť��P訌�VDť��@��R�5�@�g!����1�9��*Wu����2<�,u I�-[��ˋW JP�M����<��g����g�a�ɰCq@۽N�-�A��E�4���ǘcB���l�U���Ə�z4�_И����̓�w����H�?�r��@zj;���{�+�ܻgd�g,��G1-�w"s2'��(�?���� H�"\�}�P�҂V"@}�Җ3�BKg����.��[�ק��Ф	I���%�H�{��=>%�&Sc�=)~��	=��Wj�q��
S��g�L�Q�|����!����\�weI�UR��P5-d��F�m�ZA~٭��T3*!�^���|�G�4�&�>�/�b�鹉��*�<�v�U�¸fZ�Lc�}@��$��7��]փ*:��cs�3��k6�i{~]"�+��Ϝ�����gH�紐�5��tȐ��4��X�m�/��K�Uڕ�r��XPy��l˰f���N��:�����j�	ͱ�!�,��#�(��gC���#�C��8k��,n)_�����׉�x��I�ЅQ�L���i���8o�w]�ԂF�^�l��<�z<c�R]�0��m��k鍳H�,�P#��L���i:�Bc2օm
�جJ�4��(���a���3��Ro1�WΗ �ɣ֙=3�v[�0Px��J{������|�������~��sw����0�g�FA��\�2	��T��*	��XQyE٬��T?´�!�
��J)Z?�(�"��^,��4� �Z�4b�x���
a�+�#�g`�d(����qݥ\�~AՅB������-Ûˆ�����<*�iX�_�Dё��(&�9��3χ^���>~	V2�Cɾ�ˡ�n��Q�Ċ�������{	��Ba�P��	�9�&��B?(Z�A�|.���T���������&I���M$4.�jH���| �>����U������o)��} �HU��H�R��CW:��'�֚�-u���!:њzW�7��h��FiT$��/bW�p�'�i�u���6z^ykE�0��#끤���\;���l�j;��� �����T�o34
���n� �r�@k��q�V�$%�}o�lN�|��3j��e7I�x�L^�#m�)K�F����Y��,͚�����I����BAz���	�q$�y9��ȵ�|��2�eJ�2G�QX���d��S��V����E�9j�(��Hߚ���m�� [OTJ�5=wR����0{��+�b�9�w�Ҽ��Ț�M{T�Q)6�d�[PIX��|�_m�c���1Q��/
�������#�.]\;��.��5�-f�Q�dՈLe�ق���i�:����B�E�d6����r�(*���A@\-�3�0�sKԼ�6��qgw���] Y��r��х� �z5|���q���;CI�̨��iG���aZ\�ɋ�q9U�7a���&�
�f�>����`|�2�����~�b�^��XL�h8������T������!��DD.3�S�u]�R>��S�����<ݫI z��K�:�Q{�H��~�`3��H5���}�����sI1���|�x���KX�'� �Gw!O�5�L��X�s��s3M<Ҁ��:I���q��i��8�f3#�ɦ=[�Q�F�����O+�����b��=p����8���l� p?Nou�A풏�M�T'�b異��	C��E�/(W~���A�䑄V>\��1���ou�T�D�?E��լA�!X/��/��t�#�m�y�\�̣J�n`2a�K=�!1bW�3lMK�8�iF�*0M�}��۹��WC�~�Kq��?��bqZ�j��b'��z&�!.����>�����f%���eЅ���������˩v���q��>�9r�5:�mO��Q���(`�G�K^?�7/a_���|%ȳ��d�ǫ��(��GE�S<:C��nM#j-����U���)�U=0��^�0}X�~"�6?�7�������v�at�0n�(簪%��[��
����\��M.�;@ #�n�lC�w]e:Ε���nW6u�F����0o|p�x�cxX}��i����P���M� ��������:ױD=$��"p{lw ��A��8WI���Z��3J�}�c�i����b݀FH��C3r�iAĹ��G�Q#��~#�+e7�K���
e`�HkFX�57�
���a-ѱ��7t�1t%h3	1�5B�n�4��� [���4U��~_�$ұ�*��M$�5Ƌ��"���D�
,��wd����D	� �>!H�),���͝�j�ն^v9%�pa���`"�z?�8OjG�r�/������qݠ6�ujX��6W=Q�d�+hC	c�	�Zi"����w9�Jg�
' �X�=H�����SWe��VЕ�S�L�r�]�c��O5h7���M��<`w1+`�݃�$�d�C{�B�^wr�_����T+����l�۬�R�_�`Y$p�}����4,��?Y��M'�݆>vr��!z��W�ߢ=>�j����@�5�����ٍ]��Zov���<��;��nk��ؕL(@7!bI+����1[�~����F�.s��6)W��d��kYNES+z�N"�h3S�/�w1�3i-��%��U��1I�U���LQhЯ��g�f}�F�	A�L���E�ݽ�6 �/��.�F�p����B/Z�L�ߎ������1uj�^9�*Nnv��t51QE�wA���#yX��nM|I�
βU��nŃ�����&(ڱ�uZ�[���� ���Q5��EUߛP=x`�9w0j�d��k��q���^I�ul	��bÅgeY���nsѢp�}Rl�"h�J{Iس����2�@KQ�s-���R:ў��S��2�X�$��>���(�Mk�}���"D�XUi����t./`�c�����6��F:N �aZ��^�:g�;����3��sDp4<4Z�`pM�}OT�W4�Z��p�Z	^g�Z�R���	�6��P�P��͵�;�������XWlռ0��%1�`��Nm*#��׫)���cώV[uuu��W�)�ݭ�S8^賮)��1��aW������(�6iY�7H��)�`N/���,:��j�mj�rBͻNC���m�WƔj�9?0M�� 
��B9 �51S\V���ڏW�����K�>���Ԑj�/r5޷ʷ���{��Ci\����N�]���2ت��Vw�u��U�&�H�H�gF��:ٗy&Ⱥ)2�YJY[ yuT��	=��3�.�D�*�g�?2�����ҜÂ�����=�u�������DTxm���9�z�%=����:�)�h��g*�9���w�1��z�����I����5� �y�IJ�����ß��~Ë1�<^�"�^6�rZ��^��~V�6��*�T��(`붂�Z�ܼ��`����>�jA8[PE#���qf1�����F���[�_��B��b� ����Ly�KN"�Ef�(_�؏B]qgk8��N�Z���kM�P�ek|��)��sA�}Qߖt�`��'��r�8]�gkh����b�W0X~�9��j��a8Q�cHnO}���߇9�z,��'�'�c(��G�ZJ��P���O�A�ݴ�@{��5z:e�?��_/� V�k>���c�Z�0/��U���z �V�<h���%�u��M�^���j�\���.�{��؉��q���ޔ�2sƨ���rRʄ����5@�B�~�H�.+�}G�ZoP��l���o��E����/Y���8ÑT*�E�������%�mxi�˪��LCM�����}���M{0��iI7t�&ũ��ܩ���!���4D�M��=��Sk)8iۼJ^���K'�)R�͏请���?Е೬�����JostmT��~��cʭ�'�����l}�VB�W-:�~�� ��d�%�h�4�p������6��f���ǔ��M_%�Mhm���8w��#K������\A��b}��S^|ۜ�e6�6rǄ��Zy���Xh��v\�	�sR�~{�\lzX�6H6�yK�/F)Ф6{\�v�ⷁ�N�k��w'UL0��� �,�|����!��T�^��`V�*/_�x��L"��
�� ��,:����<d����Jw��"��7�,������DL!Kш�{Z���9/�vʭ����P�H���5Ǒ�k��C�`���2������{9i~���@ry$.�@�C�]Ɣ��1�s��Yv�}��c����=��A9�3��y!P�������R����ul�#y��ϣ��O��I�AX�o��,WL������Xק�g ʊ5�O�����KX��ⴳI��"�ڒ�k��F�v�&�6X}����i�Z[��O�p��������y��������9'�ݱI7F��"���<��G��/��}_�/��W"�^��"��?�l���RuC�������9�8�mFz�"qc�华#[���5�7T�4J��T��������s%f�rn�e`̱��iTG��${O��ɾU$o0#_��C��i�rl�e�W!+X�/]����&?���Wm�a��a���8G�GU̒��IGtv���ǃ�,X/��A�aOU�K�9vcb�~��)8O@��TN��W��,�⼛q�N�}�{o���Z>l�)�9��ם�ި)U!���a엹�.�ё�3���xk>�;�l/�uG$�6���	h���Yս�i�me�͐�~�����ĸ庆�+.386��q>���BҌ�@U�'Y�X��͖C���[�{�Ʈ�΅�~e~�[�mH�,.�s��r�"���?��r���1�[�p�-/7�=�v}͓��By ;R`<<a��$T� 䍵eK�^JǮ�F�ѝ7y��_�s��p�����Pr�0w���	�`� ��9�1�Xlx�k��� 5� �a����5�!�^b:q,�}HU��{��VL4���LCP��7�۬�Q���=�$�Vf:��āi�9���_b�F�ܜ~!& �UU��Ĝ�LU	�:X�sB�#�p�����~az����toI�_yT�����a�o+ǳ�r��b7���s(��,S!Hy1��TЭ���*�hPO������@HҷG�k]���)��2��J�mx��/A�P�
K���~�#��b��3nHp i�ӆ�H�����!�-�C�Ki0�g�6%��$1sw��ew�.֓�c�9�M��mr�Q#���?4~9����[���1�PN-�����S������e]XØ�]�Jq{l�B�稟C�6����@�T�s�Z덏����A�ܕ=R���ً5%Ԡ�	ӐI��ʊV���`l�+�6������B��;�YW�8D>e
��Fk�WR>'�,|5vŷc |��x�O�Uh)Y  _�����ć����a����z6�4���ݾ��1Z�"���0'���*���ڎ6<�Xh�k�s=@r%<V����eu?Ϥi��O]ݫa-,[�ɜ*V�"�����#@V��L%g�i-թq��G��/d��U0e"�����E7Tz\��7���I���*��B߄�ƻ�!p{�T�ҧ*�za�݈� rK�� /*
콈�-tUhE�§�=@�<�jqda�)�i�>�Θ���v�#�D�u2|�\����.��v�ڹ�!���'�}g�s:���k}���/��M3�O��j3�헏eo�8��e����͏?` ;#�H��[��*K"��F�q&�)!t$��e��f�_�����$�;�Y0�\� �h���S�Ձ-^|�����E'KQ9��ֳ�0�`�螲��{��R��S�;��{+�w��o-t���-0xq�s��\���f�9)f�:hŲ;Yݢ�j;	���3�TO>��\A t��ТI1"�&y���;���"��53-�|4Z��(��2�³��C�6ܢ�)���A4 �)����aJ��&�7=��a2+�:���|���\�9�U���ʼVh�-�)�y����Y4M��AS�3�1�xs�iA�7�m�a;C�i�� ��$��� y?���׍@.���+8�ovy��3�n�}��>�2��ď0��;����)�=b�K�H��"�~��#��LH��kQ���6?`n��5<�m��e7��)�o�t8��5��s�g���#M�1��޷x�w�QzL/�q����y/����<c���dk_�(����64����Y����5����$��%B�m�0���hv��8n�t)���!y�\�!������x��C��C�~8���4(2JE�cA]��Rr�G'�Ѓ�1��$���&��	D�wa�\���;C�����ل�A�;x<�������!`�o���a���c�`��9E;��5��]�=�,��}����P+��.(�$[�P�u���^	�GI#A��O�{�;���]������A����>�<��JN!hg�Î�[I�:�[w��'|��Uk����	��;$���vaw�"�9��`5�����X��Q3l���{|�(p{�H�ry��+2��/�Fв��h����a(U|���p�1��b���aF�G���
�*�3u���կ�%@���j��!e� �����CB�KU���[sg�	�G��T�
�����*���
u�K��RIqv%�����H8�N���k��y,J�OF��r�����W�@�E9��!5�M��I�;�o;|on��`�g�m����N�3Vy�忠�G��I۸��e�<����j�l��� 8�ޫ��ڪI:�s#W�^0"�G7f�'AČ=3^�F���q1�Ot݌`J�1�SD�ݰ��<�7�N���~F�1�0�݀Z�����u=�����?Ⱆ��>�Y�e/��y�&�ÿ޲n,�F�r��J�͕˳m2N�p�����+�W�`O���� ���̏�I��τ�TW1ė�>pU*�(u̬i�)�#�O��VhERzc�f:J*x�cM����z&��l�de��{櫣���o�ݓ1$�F2Ƅ{8t�?��fv���4�>�Rha���S�]����"[�tg·���(��`�5�H���Tk����>����b	&����%.�N�_�=O8m'�Q�/XgD�^Ι�
�shtX��M��]���f�F��À-(m�&�R��!���"�SlJ4%��_�J�&�_h1k�\�D�B������mj
�"d����'�Z!�����`���0��} k�ڤQ�dɑ��y\��Ƶ�"���h���4%�>e�Vis�`�)�2��4Hc�Y+���@��H$س��٦�J����N�����>�%�S�	 �2��i�������=���N<i�x����g��V��բd����]��rW��[l>5���ۗgi�k
�+���F�He>��Z7�P�a����'xs8'~�w��ms�zNc���8�� �og�W2�	�u��I�@5<64����F���ͳ��Nx$�铀܍�ϛk��9�����"�~ˍ�/	{\�r �+�oIZ�]\	���L��r5�Tz3�������`ހҾ��@D�\�o�1N���a��ҷ-vUy;X@��C��{��zR��J�h����E��d׆=aᒲ��yJ���	4�H�!I�3�G|�X �m׃�:~��""g�0�.�2߉��.�M��!�B�k���ԁ���r$�R_�����1:�f��N��e��Ɨ�[S�:\J�\q\���t �z"�9��8��.��F�t��K]��2�&?�����ޡp%Ue���rJ����Ql� 3/]܂k��}�[$�A��5���)�Q�)�F7���	j�>^�R�3C���{ρĘl�_SO��y�#�J�*�y�޳���N�R����,LD]�Sɸ�"D�%4+<2e(��a8O^�=%�	k����o�kx�T�RP��0鹒f�
�����'�"��(�'4�qHЇ��S��2�����6�� n�Z�帊�d�Wכ���Y�N�ML8�2�ϯד�-��>�·Qc��S='Z�YJ�֪�B%�u��o����;Ӆ
��˂ZА��ev���O8:�`�~!M(����=�Z������mX�4�EE?Hd7��P��w�m���R%��~QtT{��¤�see��o�J�t����wX�G��-����c[��Km�@�����_z�-߆�2�������?|��(�nD@m��Lf��F�GP���r>�I�%�~T�����4t~�������<�^�a=��ɏݼ����j�5ب����ip�tY�mF ~�,��J�<����I��`�*Ř
�x6��F6�����GrH@dz�ҫ^�v���s��4��&]:PL�1>�T��N���@v<�A�sի���qUR<�ht���E �8pD���1�[����l�|���x?ߚ����XG�/�K��.��N�
�}:�W.p�i��̟$$���3�b
��:<�����J,�
*���W�Mw��*͵L�>?aMކ	��x�:��� ��1(�%�0�g�1�Y@W®ݣI%|[k(EX�������\ӽ%̿'���_�e���;��� &��>�����C!i*�~[	����~\;��`��ӭ��mP9�r���;�`͘7�ky�~Ⱥ:#oOV�-FLm�q�;�x�̢u��lր��Qʹ��13��T�g� 6�͟(�K�k�G=l��Jԫh�T���e͓��T�9�J~�P����m�[�~B�l�6(�Ɋ����Ы�ڬ�f�"�`Jו��C��FC2�F����2VdX�w�<.�L��O?y9W����2������Ƭ�䥁�+eL݉-�L��k����Ȉ-�a���CIJ�w���|_u��CM��>NAl#U�Ûx�J�F����Ê�q{$��<���H�x��~�'��:��F$Ivg������@2�@�,�^���]�5�F�'8�F��#�w]��(�/mكC�֘�|��+�����W����!�P��ol!0�G�h�A�����@{]��ü�7��������_�wbT=wj�\�)?��S��c�ҧ|B�I%w��%����;�����M[ڂ9��9Т�Y��.�����Ӡ��R}�px����`�����	S�V�K�ۡ8&z�Y)`��F���ֽy��cJ�.,�G��rpS��\�nVK�w���4~��)�x�\�7D��.�g����k�ˁ�鐦3��."�����M��\XP5N�D-f�\�p���#.oү���lt?�'�����2&3c���c;F�'Gd�0Ï�^����6R�5�Hm �������|$%h=�m^He� �<#�+K𱍅���h�jŗ\���.�VJme��9��參�DG3@s܁|��y�+��+۵�X5��v� ��8`L��sN"�:C���Q�,������q�M�_� ������C~�G��W]i�������\Z{bۦ��$+�U麁죙E\0���1��_mD�T}֞�vbT�2Ws���5���YZ~ ���б���8L�)�����	٩o����7����^[h���*�tj�?�S��V��_X�ٵ�Ǯ?N���+u���� P����f�w���ӊ0(-RI��5�!
��ٵ����!�������BP�����a[HD�%�p@1W�m�C�/�;�s�ݾOy�g緔�Ǽc�o� �\�&o�J�����s��KG��Z�u)�ܟ��зq��M��r߼��޶�P'�����.WZ̜�s*�<�r�WJ#����Uf���Ѱ���DW���H�(9}�c)v��B��8�����D�;��L?}j���o|潩u-n
�68��g�O�s�F�a���L��Њ#�Π��O;R����=�TjiE��͵?�]!�q�}��A�W|6�M��Db�Y�oN��#�Hu���d	w0yN���jF��J&d�˱~�Tn���4}w�J+;�ecP	��)}��>��L5���(])��!+��O�)|I��0��$��*���󫆵���S5�M[	�C�� xT�h�V�ݰ�Ʊ�F��7J*��7;Xt\s���ף���a��O[ɷǴ9�����(�$R"p�"�+_��Z�.�$dڧw�������	�0~}�рB�ana�-9��s+���h��T��6Ġ\��a@�ͽ"��l�W���%�.��D���uׯ+-����3c,�bf)�fq59'
_w��̤	S�A�)�S]����Ss_Jٓ���f
%f�}�AT��ϔ@�/�|��a8��7���Ĉv\E������1l��~�;�!+S� �9���>x�:�i%�����ޖe��G��z@�MP��|˪��A��:X��Ϗt��"�E�b#K$N�1�+,#(M����9]m$��_X+�#�Qy� s�qT~����p�,Ǌg�'M�o����y.�^����4������S�j�����6���LYY%���@ ����S�[q=���V�oE�>q�3�F�7�A�51�V�1�<� $�H�QM�Oiv
0_�g>_�)yɋ���m��B/H1�8/�k� ��u5�`����W�tؖ������D[S��㩄�>n�aE�����jph��HhNVoй�
eZP���?���t��e��a_!��u����u��1[�5[n�m���F����;OK��R�@m�����:j��z��8���F_��G4��(��?��S�}���"qV)���߅F�:�{�U�̄䦮��H+�4U[�&�,]��p([ݬ��Hi0��ً�Jc��QC��c�Q櫜V�yw\���^La�Ӽ�s�Y�攲F�,��N�W�OI�\�5�`�P������c2�|�섔�k��E�e��O���@��C'<F˝)
�]�[)_�s����&M��G��n��{z�y�s������˲�wT)2Xpv�g5 �x�tWTij���ӑq��m�r4����lXqbK|��+�O�AI�?��4�Ӆi��f�򤴿vU#��h��^3^�!A�*�޾��q�Q��ҋ���)n�&�+p��i�3���㞪��6.�O���O]�(��"���Қ@���Ch�	1 �U����C+`]�[u	�Ww�ū�k7�w��'E�dR�:c��0�V�K���NI���a�}��mEr�R�}� (9N�����#�-�:f��T$�i!h���gD���u��򠜦z5!������;��7��+��q�r�[��k���7:U���/�Ų��Ow�K�Ǎ��T�c\�5��&7Bj��p��E�8}��pI�e'�V�>��n���ѳZ�R�/m�����g�x ��2�q�V^����n��
X�D�R�����,S���{6��� E���]:]�Sv��`E��O���߲0�q/��!�p���*��	gW��p	��g�m�d���Q{ItԗT�fCݖ�~e!����|��L��SN��6����T8��٢��gz�G����l��sb��ޢ�����"����[.�ĆQ����kc%���ժ��g�E��bt�0�O��eG��VK�u~>��8P����k*���	s9�
�urg�?�w�U<�3��?��k�ɽ{�J�ʏ/&z��z��z�B�� L���Ջ4��/H"��T�����J��U�7`�&׊�	�蜓e����.�3��0��\�tAs���qݡ)̴�S���l�)��# ���T/��(yg7��E�,Cg#�� ��NJ9 ��������T�k}�4�6�=��ް�O����P� ��{��6U��5/�XϷ�q~�.�}���@��Mj8��mj��Zz	`����uD�6��a!f͸����A7���{���L�c���j`O~�טgzA��7�l�䯬��@�:����ۦ�	Ac�|�L]H>�vI���H("��c�{VA2^������1�L�E3SN_�J��:x�G��P�����%#���c�V�e��
\�7��ۦ�%�W[@��>tT����7S��b�
)T���i��˥��U�����w�T�s�KE���u��{��=�ŋ��s�DF����R�~�����y+5���[H<Ħd��Yr�����_r�W�i[y`��2��j��H<�q5��%�kh��r�#�3��l����V��dD�&��#���Zqy��X�?GϙY�2���ꣀjcGE�])����0���{
1(=P���>i�ز��3+AP��!.Y/�`��I���P��S�!>�è%s'g0�'P�=�Z*�x��/���걃�����r�o)]�O��7���N�J�nYx�� |�˥���u�\��-D��m��'���.j%	I�������AR��up����b���E�{+|𒡛��<+���~Ԯ���sr1�~E��9��C>cl�l諚*f^�x{nP�n1RmU���d�56�E�B���2���d�7Q�+Yޛ�{}��l��p�7v�7�T&�3LE��*�G��2	h�n����,Zi�Y`4%+�$o�i�%��P��	]��`��YJ�OK���/�����U���Ė�e��V*��P�ߣ�������M��+������Xt0aW�M1�pCi7���b�u<���j{�z��mOU�5l�d��Q� /�sb▦��4rR�|�]ڇg��R�p���e�#�7��)Siٝ�ɉ%��0<�����f���qė8��W��2wGJ�c�o �o���t��Rv�	2z��1w�M�����I���˝#\M����>����U���ݯ�%L���b�(Yz����
�B��9��B���p?6��]��U��7�c`ﻃ�0����j��(r"n�϶�,�^�D��4��7��x����?�;�'m̦OC����XAt�=Xc���2�1Ì�9jJ�D�C������Z�e�p��w���0�+D6�G;\ן�|/ �+8��U�u~�	b$Q(�'´�J,ͶO%�C���0�$|)o�*޹���Ś�9ا :��ND�
����)�9p���d����mע���(�����U���f}m����o~��m}�|�/%W�i=��9}�6�����2��T�;���ݼ}"����Z���O&���<��븗�͖�q;�䛤�S$����RG��(�8����c�T�wl��Z�!�B&ߙVE>T�eUƆ�%̖$�@S�d3�K��	���&P���{fI�|��Z*�GhL��H�AVB!}D�?��D4��Uw5���-τR�����
P]��X���z��/�$r�*ʶBσk%�dd GN@�:v�|���\ԙ�j`�;�!qy��!ޝ{
 ٢1�/�g~;���s-����WGo����#����ͫ��?�t��*PkK3I ��ϥ��2��,�UE�b|4r7df�`FDj�2�p�a�o]`ha��v(��s+<�P�7\^v_����ջ?��
{�)���ocQ�JO�^�w�og���"�dĦ,�䎋�B0�S���1�R������qQ*�P-_x�ӓo0d��K3.tFj%��Y���_8/T7U�-=�!p��ڞ�۝���)1d�������Qg�!��װ���f�/� �#7�Jg4�.7��ل>�vrXЀ�KA?:"�K�ńr0���4��XMgE�c�wf����(
�w�Fl|N�"x�~����}�i��D�h�O!�^�;aw�a���u�(�E���zt��	q\����JrӪLF�{��D@�k�{6L�L�Ox��P,¾�x��)�[O�- �0k�����5{�m�Im؛ኻ�5Ӯ�(��e$��"e�����y�/��.<W�����J�Y_]��Q���f��D�f�5�lVW$����$�$�@R��AD�b=�p��.�^.�Ǡ��?�����u�3#�����[�9P]B��P�}N��7?��6��Ps�O�I�MW�ښ?��T�����+��q%�6�<��U|��>[�bU@7KC��E�8ŕV�x�0���0*��@����!���*��gw��3L@�!�W@Oe)�Sm�_��=zQ+��u����{�Qw�Q�dZlV�q"�*o�}A�2i���yP�9�f9���&0r�E$�دC3sì�(�tÃ�P��W<p'ڃ�בM����t��&��4NT�����E�U�
�ߞ�OK�5��x�Mގ�e?��S�B��q��P?�N=�D�rA������?A�qz�X[���xM��`��S�\�B�	A�e��Q.wX�[��B���F����^<W�x��7\��/��>9r<�Ҽ�k�s�&�T�H��#��ٻ}�j��T𢟆���2t�|��d��Y�c����!����}<#�PRl%w���ړR릸�����v��B��:������f��as^K+J ����)�&
`��`�b�} �R�ox@��fsY�׌�a�����J�Be�xkO4��¼�'���@G�).� L|�'��h<3�w ��$�\k�2��7� rp�n8���BUq*����Y0���c��=� �j�C:���P�UzD-O�i�7�����N��`���z�Ș崄A�+���{W4Mm�2���ߐPٮ8��d����b�C��2��yW<�YD�^?�zM���Y��q���5=-}�z������Ы>�RԾ&�HD;]���8d�����{�F����N�k����F�%���:��V1��D���G'I�xZ<U/��� qQ�����Ϋ�n#�5h �����3+?����PĢ72��;ص��A�P��ᬷL}(�hA뿇���1lH@�e��o��Ƕ:aot���.��T�~NJ̇�}Ȉ��+!Nںq�rѣc�t�	�Y�$��gqЎ����D���z�S�	�HD�e>����:�ǣ��'=%�q(��������K�CXM��!5�>�o9�3��Ü9����C����?��s\P��?��J"�l"�Aز�ܽE��^���a�əZ���.�vj`��i�=�����eCG��4�YI-d��zYܯp�e�w}GH���t�N�a����1c
q
��]`�y�%p��+8t�Nd��_���8Ӥ^{.���W���4����0=��e�H�vH��j{{'v���Ι�I� �Ҳ�����P�Le^W���Q��o�E���޷H��!	`��FR�����$7��d�@1���-���2iƽ��&�fL{2Y�r4(-t^l"�ݡ��c�

�+B��4��e������Ws7���r��}�Hҕ���%�6��d�7nl�<�{��$A�W#MO�Q����_E�s��f���<  4y�-��I�d�퇢���-���d��<��~���	\梋P���B{s�a��?l���|�����Y���� � ��bl��8@z\���u@�&hJ-I����l���Y�B�%3��3x�c�7�ɽ�/���u9ZGVmN�I�"�:Z�1���Y>L�dG��ٳ/�A�|�d��q�Pt���,�E�ڮa�1�9F!9��6�{�.�&l ^�V^���H�д��[J_T��(m���Q�1����G���8*��fi&fM��0��i�p�dÜ[�	�����C�
�`|`Պ���7Y�rB��0I��j���JෳY e���أIe2�]�l"��ԁR~s��ު�5[��[OS�  +]�>�"�R���3�i7������C�ڽ�m���j8V���k�?B�T�6�i�f��V��|�*d֍\�U�J�U�_��3�����G@ƿ�Q|�n1����:8�KfQ�]&Cɩ�G���M��&�G�]&�]�j�?ρZ�zV����o�v�q��ME�cnK?��M���X6ԏ=(��T�=b�o�� ��'ld0T�
��'Ь�܉y-*k��TK���}}�̚I�a�\e�Զf�b�!-��r�窜oÙo�Q)?�W��V�H������� qf�*�_u�X�J�y�{}��h�պ���sYR�Tq&.Z$0�	���=*>m!�:Ƭ.�O��D�Ƽ�&�P!F(�Ԇ�XD�\�ҋT�Bo���a�өWy�څ�jh;(���?���@�:����\$��ڵw���xA*���G�Az��y��L,�G��.]�m�=�6�.���+��qH(c�� �[�jA9��t�S���^9�eQ��+V�Zm >�1�a�BN�4�әh%KI��x0���	5)Eu�f+H�/�9v�u�gWKa_�I��3�F�fE�{������2f�e�)/�i���4(Kr��3��%j��5� Ŧ����O��ŲVo�z�B�RL�g,7V��
�$�Tk���q.��)X�xm"��h�k@ѹO�J�zL���P�..���.�W"����5�Eż�^�́�~����X�K���B{�����
b��������t�6tBM졠H��2	��A	b�� ����G�^aB�&P{�1S��,�څR;�M��v�Ư�����S�9�قF���T
�k"� �aT�I?Nk�tl��l�u5;�"���m��
���Rͭ*�u���������l�<jn'�'�G�\B�8�U~*�Rl��$DNV���~C��lj���i�n�(����̜��LCd�c@�.���W����a[�=�� �)����Ql8�Z�5
�A�T�ml];��i�9�F߅��I��wA�]*R�X�1:
���W�?�]Oѳ	C��Eڝ����v����z1;Xx�����6�l� ���u7"2���n@�L�j�O��D[��@c�q���-/�p#!!~�.��nA�U�����K+�{m�� G�0�������g�k���Gz��8�;���4Vm�7��`�xwX�az-v�{g�%p�Zĩ(ԭC���O�7�y#�Z΁Ir�IMK�M0J�w�"r*�qˍ2��C����4�3����0I�X��'�6���	6���c�|jqؾ�(D,��Hp�n�#�C�NsIR^s�Γdcr���;���Z���;Ew�=�л&�7�U�`w�)���%���yX�|�u!�^/p$�r�].1�9i W��𥇧������<��d���Pe(�'3��LR�%�����h�|�_���!�U/�E7,�:�.����S"�@&�գڿG��"���e �xIz����r���@Z�g�A��l��*���Z�т��$WIgP�����,�>k�.T��zF�ҳU��\T��y&���_��𚯂,_�ZϪ�m�B1��60ϳ��xqǳ[��~�9��]�ﳈ;k�ʛ��	G]��K5ϵ���<C���!�){$!�h�x���!�{�� %�Y��4�%���[�I(��,Wh��6�8�iف	�l�R�qI����c;>����܁ބ� Ҭ:�ե�_���0&W����pŀQ��noVn���aP	��>:[2.���(��PDo�#�f/��S:�Ä��Gv�q�MO)ʭ-���5���.6E��#vXU'nsiTZ\�g)%3�-Ne%�
b�������Y&���h9?7��xc���u�v���dc��r0~�Y.���c�K�%G���D�gj9�@7-�,}3a���ׅ��M�{A��i��a��CxU-��e���i�Mӓ{߀Tx��KhF���	���cI�T2.2�Ip��v�$+�zS`#!�>�ք���h�x�����5��cz>�"G�͚�����42����ኚm�����pb4������T8m(y`�p���4�����s�d��N�xo'��y-.���xO�סjH�D�����-��wh�[�*Z�6�z���8���.�/��4��SHH�#���ǲ��|/�b��6a�c��T��id.T�;�	�9���ļ���l���f�BڟN6��_ۊ�t���T9������4g(�2���P��l�:|��I�gE�ۋ����L�o�W�G&����Sw���=��/�T���O��V���Ԯ0�:��b��k��Q����?��qw[,͢�O��དྷ?3��e��"�{l��
��~}
6)��f 8�6�c�ILC����^�E[�3�jfne�J45��x�����P�A��(*,ܾ�r�X�W�Ĩ��J��L1� =g����`Sk��_���/�tQ���M�#7�{�6Gz8w�M���d���'�Ҩ��cR-�T�x�\;�L��L�Irc��K���g8��f�;��=��s���¦pk�������K3�v�i@M�%�&ki���D��-)�$B/F?�͉;�Y�ڇ�jƍ�x㪶�w��-<���l�1̕�d�gVX(��dL�hw�`�7ERez ?i���3�7oqipl@�����lt�|>[���:��������}4�|#��usiL�3�2��7���ڀ�P<8.6opU�wB�3�Y��O,�G�\�°�iOER���Ώ ��jܘr��zo̲���PIK��',��`�d�B��G�fӏ�l���1�QVucҢ�t��¢��(�Do�x�虽�)^Z���Ʌ��}�4օ\(���j�xh�6N�˵�6��z��)Z�'@Ug��q�Xe#)t�����%�U�U{iƖ���S��e6�����
e5�[ưB�#��J: ��h��w�u�B��4���$X��DW %t1�Ǵ�}7L��7,���I�Y��" �S�e��a�������D��oV�u��+4q>� n:�A|tU��� �*�ѿ5*�ؑ�Ap �.P�l��hl�W�З�>��@t�U[���� �&�.�(�_��6��/%�t��/\|+�A.���#�O�j��G�����[OIu����v�6Ur�{�G.���}��Du,m����#95N��̪ء��N��������p)|ݔA�︕�vB�z7��N���guK��Qo>{���E�yj�nH�S	ba���5����i�AZ�gN � Q��B�-�k�&�=�:��i��\;�2�}�&WmL[b��B�Zr�5�aE�����%c�[p�L�gLk@<A
���N�W��̛�pxgv�J|u�7�]ɲ�g\I4	�@�e�?Ξ	e�"<�`������*�ƀ�ͷ����[\B�$ ���ڎ�p;�{�G(AAZ�~�K�&��2(�a�;�Z�Zj<�7r��0��,�nֲ��� ~��(
Cq���A[�4<�aW8�"���#�AfƓ���~��/B�36r٧��;�0ڞ�`��4v�*���\Z�:!~s��O�Gf��8DQ(�/;�sC��LXA���#=���9������Fӵ��m��}M��b9^��s�C8r�-5��W��U6��M�p�u�0�Y��J�Z��8f�5`�
Z&T�0�(���?�~4�Y���L�.崁 ��hR�,�Zw�9�tY���q�nvs�����P4�HN���x5p4�\O�j�k,h���ܮ��<�;����d9-���D�|���J�Hs�aR)՞��������/F�B	��i̃bK����fV�{d�6�����]�O_|���������9J�If/Yݒ>V+�%kZ&Ss��� ��"�0���>iŝ��</�>W�v�#�j���܍��@\Ȣ+�Fۈ��~�UlU'DɁ0����ԏ��w�@��M�W��M)[��%��n�N��<��J��p�6D����^���@瘏'M���]i��}S�R�-�C����{���#�lQ�ybA����0Jx`G�~��ox�'�I	M���(8�*��D��C�V<<E����W6$���Nw�w�����Wª޶��&%]��_o�� 9`�d�� �PM3�F��:����%�4u?��.B��ӑ�]	m[n�����u?��DI�ܢX���b�˓�4N�]
��9�/��3qܳ\��^{O�$u��˂/�b�.���@\
���]�>�T1<�]4�i�F]�3�/�͛^-@��?;��L�|x.��!��!���A��{�·�Sd���D@9�N^���u�g�<i����ܹ��]��&ҍ���s�m<�Yq�w� |�f�N����)������ �w��D�@ߦ��!bZ���.�j\G���
O���A�K�M�[h�����X�d�K}c����$��:����Џ(��1-�Ydkhv���x%��g����F��6��0�9��2���v��;  ǒ*�a
�La<n7^F�����eB�e��,�κy�� 5�3��|L���Dt����P�����/���ݍː�݇�0J�%qB�1�a�8R�����GU����[��y��٭
���|N�.�Y����"?i'�Ul�v�������b���M� �}�BT��\f��@�%�e�y��� ����?Xp�%�����<����W-�$�ի�{��WQ�>?W�rQnof�"���wqp�a�J6��i�D�`0v���	#<�Hw�R`Y9���J~f���X�(��+�z~�c|���+��۽eڐ/qae?��S+��xײxި�U������(�r���Q�ɬt�دﾇ�"�;�EFL	AK�����B��%��|�A"�4� kS>1-���4��[�)�r���6t0��q6���q�Kȭ�B��L��>��w6&G�R0=��MP�OK[倣�3:^Ԃ7Hnx'�Ɋ �~"=N��58g��s9��rBโ��y���J�G$7G�:i�AS�pGy�n�h�<'���wH ��&>��7�2nCO���<��+g�i��v���50L[L���i���sX�O�-�5rt��m��VYgu�KS!�F��&�ܟ0�%5DA����־�in6'�c>%A�.ph���W������j�v4]��E m<%��B��bH����V�O��S�j����L5_��̿���ԁVUh\��"K�=�EJ��M�K_��d3�jL�M�f��o�N��� �pu��vL{f�(�m�8`r����P��#�[d���k��2 F����)�U"�0w^�wf@Q��H�r�3���HY��,NR���?a�eZ��Ȼ��l�V�x6�V��),��]��P�I�c\�~Q_Ra���+��z#�'n�Qy�3���p��#Q\���k�j&��Qv�9�j�>��ֳp?^�γ�6�=�3{�Ϙ)d��kgu���):�gc�d���B��C��@g�9L���^Xℿ2ץo��ɍF%��w�Gw�:��I�}�[�U�Ea�����t��C\Y��-|8E`-�-��4S�U.x�� ]��Y�w'��!�\�e�k����+\v�1}���ƭ9@���]��C|dt@�|��q���N�����]��.���/��������9u�o��\lz�Q��7cC�>7��ؤ�5��5s���e?��%�,Z��i,��Y#i[��BMtjl|j�j���f?��he9[��6�v��m�Kߪ�=Mx
U,1�3�H�<8��Y���A��h �pӆ��/���p� w�
V4e�u�<tޒj�R[MՊU���){�l`/uR�c�b�ayx����>��:nu{��� ����`�]}��������©�3O㜰Ď����_}�r�n[�u��-Q��9%���QJ ��Qp������d)�oV>l��]�����o֏���b�|��i�q���?����+��=n_�y+-�%1]c�C�D��I�ͤ��di�� W�B�Y�gr9h�ݗw@k��d��W�W@�.��dx��ƨ
�q�l�} �轍�-��^kEX���?��g�!gf�~��2@���ΌwV���Kߔ6Qw~^K��Ip�cP����I�?6�����@�Y�����bZ#�׹n�h��e��#h��L��� �d�{Ķ���B�:t	���AT�E-�y/�=�6�B�QtN{��?ٕsF������W�I#ւ���
���o����l� �	�3���4�� M��?	�ͻ�`��&Y&�z\�	��(���R}���zR�����	�l�w>��7�*+�h�6�g'�y%�9���]YE���{��t�.Ev�e?:L�+=.��
�W��>��y[(��o-��������\J�:���/��*�hVS�q���jG5�#u��XS��އ�|�1#��F�H/������Kp���4��VJo�Y�}�*3GYp��bF2��2�;h&�|���9��9Z�5:Y.qcc|t�L�������Q�ڥ�d��ɵ���주4-��f�Psq����<+BP�g�>'���l�R�7��d��}�dE�\��_1 #�� Ў�O���]�jJ�4��#�W�����iy�+{��*����?m/����Q&�@y��,>�0Z��*��V=�ْ���5�|Z3�[�}���Y`aKqG��]�u��f�b*!�QɗI�Ԏ"�e&cJ� %�{(i(w�c����=d�S��)�w\�6�p%S��W�o5��jf��:^��/�o5T�{�4]�!������n�s� L6��v^������|(�4�C~�/��6 9C�����Nm��C��6���"QD��D��QM�gC�&�̟]�4y��V���̊��h4�-�/���[�;�p�������?Zz��,�����C�1���uᴇ���3�w�KL$���e����&q��h��+��nѝA�8�{�V�;CR'//����7!˟�&�".��t�pa�`KmcE��dOAՙ],H�D�#FL��m�L��)���DU�T���߸���K̷�5E�2$�V�V2j���)r���`Ղ��3��XY��q��W�StU|a[�9Ub��^�ϰ3r�8�n��\�x�˺EX���VRv5I�>�6Y�-�|{*��p�e{�.�<GBO�Ȏ����t=}�&��f'���vt&����#��r��;���v �I�/�_�!ԭZ	o��pL��d\a:�XH�G���G�㉗,&
�����wt�ɽS��ӛ����f��׹.�N�MG�
��cOFJ� X8ҽ�0"�h�%���OQSMYyʷl�׎�k�|_v�+�<��]�E�¹[k(�ƣ��ˎO��~���a�[�u'4utfU�����>�-�3X��e�k�ۗ�vY�rw.6��_�ݚCQ��MPϧ�e���Ƶ��*�i]f���}��μ$w��c�$S�M	F?SHKC$���f�l���|@��4І�8n^� P���	-��������n��	�l���4c�N��z��6恈�w��Q�wh��et(�	�T8�HNBK���&�ᒳ���v�j����8gs�I�@4��'Y��j��[ɶ��I̰����� 0�3�~������=mY)�!@�f�ů�w���To�^<WhMc^�au'�菊��9�А�Ci���o�W�+�Z�d��)gd��6�aG!m��Zo=��m�:�{��%k�7'�����FJgG���6X�Nv�R��h�׸7*�n��ʈ�<͢���#���܆�5�@�Z�gu�7��9# ��U�mu?V�[SaD$xZ�k˨�Arr��h���o:�Vp��os���<	��f�MDq��ټ��q/B�1��&s+LE�/@��W��f<ک׻X�*W���t9o{D�{5��5���b9Q��5�d����|�z��O����b��U�����I���(p�Iɍ����b��fP'��,d�".*��_̾���c�}*u�+�M2���9�i([pCYC�>_y���r�:��o�D�E+;21p1P�g�Cr��HE�O�5s�-�E%~��+��6-=}{J��Xo�P�W߿��Flo��r�'�UHN��{`V<���ya��\)�YyRmib�j�|m~{s\��.�s�&�YjET���_��r��dm��+��뤔�s�C�Mi�8~��c���T�n�$�d)�P�vp�	5Î�_>�`Ǫ�~�k_T�e0μ�3�b���S��?��>�G����^��z@��9�\��0�r	/^l �=Xu���9�q�h��p���m�������OtLKN13�-�o���hp���iVYg��t��:�C-�		��ԝ����_Q�h(S-W:X��1�b�,��O�_s�pt>�C;�b�7������=�y�SCW�
L5|�ޯ�o�4[����{[�;K�	'ޢ��C� 1.Vy+S�m{�śY�p{�����>bے֨�~
[��F�ֿT�g�W�s��B�����.�����mLV��lw-@����IOF"�"ϖ/^4�&[���z2��_~S��0
��;���$V�6�sB�g�732d��_�y"�q�9��ٜ����T��nZz{l����om�л��zlv
98Pb�C��"�o���[(�],��IzOx&䋠$���C���9`���}rt"XS�.7<���x>���꬇vK䞂=1�{6}��hS]Kb�E�&L��},"[��;�ƭ喝��0Hc���#A���I��.��z��c�@*j�#)��q<�)���ynR���r�j�����D"�̀U\��q}�W�Qڳ�P��}VOY��	��n"b�p����ְ �T�ԧ��&a2?k�k0� �r�����N�=PEsŉqx����������Y��x���=qΧ
����g_���0C��A�jN,��F��-[��mbB����)����P��
��|Z�i	��V� ��O+��T{� ���#���O"��u�zV�W�.�5y7I��$��s?�ٌW�n!�ͨlv���#�s���o3�Ĭ�h��g�j���v�^���۰���Lm�/�(��8{�3E8bq��
����b/$.��i���͙]�����+�� Kp�*A'2Y岮Ў�[-c�D?���Dy��1ޤv,7S]7W������ׄ�.�L�Kj`iz�y��g9ƴ$�ik���	�0౥�� ��~�SP@�dރP�� �-�QA:�k�t��	�����ꙛa��{�"sA�T��x���t�NIK���w�UX߳AF�~�[#��A�5sE�(�|UP�&�f>�����s���9?�"�k@!j��į7p#��{���8���Z]�����س_��ćTw��_��@U�T#=�3\�m�W�N���v����vG1ۉ���erܫ~r�����̨*�z�����$����<��`���-��+���\{���@l�g��ps, �q��.���;��m���w	��C��y�'�`��GJ�o
0���bF��ҷ.`�G4�yL��|	��~3E�Ha��4����W����%�m[(lŌX+_B��
S�h	����pI��S���GS����]S�ڠO���9�T�LK��Q�z�g�-�Mߩ��@&H]���|S� m�Sۦ�kWCP%�0����2�j�]1��l=�8���繚�����~K�3#5�
�2�P�	����F��wD��m�����F���b��+!��$jq��`s��)����:�E{�W��1j�0�9Ϫ�o4pr,:�&�j'�w��g��/���Uy�nm����\�]�6���t���B�&�������P桉ct��+��i�ʌNĺ į���rh�2���m�cJ�}���W|���#X�{<���G
���N<��c����F�z�`<�L��$n*��d[O�Ҫ�n�ܱ]�d�`���Y�]
X���5�[�hɝҡE�w��T�c�����E�C�)��6B���xR	�������vRH�'���*�ː�{{���4���p����*f+���#�!c&u��6�q���h��Տ!CMᏸ��9��\~ð��>��,���+��thw�G�=���G�g�=��� hʉ\_V	�ִ��ץ���Ħ�Ӯ�%:=ci"��t�)R����{����#�7m3��,}�r{�'��I�v��`Gs���FL�M&��íu��I3?�H��?��h��ó|�
���0tT�� ��%��_���������	ز�Pd���21����������j�&>b�s�I��������H�u����8���/XƬ��\2/ILBּ�)Ku�7�Bi9����M$l��z�6ְz�\�5.�e��,�ՐK�W>s�4U�`���8��%8�
IX.���RBN�B+4�E-P;��W��9�<':JN���tD?�@�����b���q��o��4�����JzBy>��3�XP���m;o��w�
��'R5yf��х�_
M�r��޸Q���{0���^ǩ|�r{�!d"�XLǿ_ ?WC�߄Mj���@�Z���Ł����ڃIS�H�&g]!|��9��?�&�Q��<ut�Ҧ�C��He-�U��ص漌���s£�i���ǖ,�<�mB��i9�G����#�0;�k9;J4�e��O�HŢ�n(�y���@��Zg��W��Xr)竾��p�[s������UD%����04HMhe��!۟����<+��dŁ��M<mJ��ϴ^]ȗ�q �`a�`y���b8�n��5!��dd��w���hS|`�dT`7�tG�1�����]+x֫w~����yuV5���.F����?�Kae٧�B�Wz�#:�F�)`:R��!d�������I�}L�>9X#0��	[���A8��Uenz��ٛ����Ə9������[�Bbڋ���;n1�=�KM8XW�"�u�͒n����H�;��1�����ؙ'bC��(�l`1O�q��Y����7�M5h��6����4/vړ��<���ͣ�t��Z� �IO9T����"<�����j�hhL��Q��t��W]P� }�I��wR� �tuE�d
�.0D��T��y�U��������appd\�D{����ܒ�삊s��-����Kx���F.��"E���#�,�Zr�傳�/�ۑ�d�ǆ��<�.�ز_?�R�+�N�
�v 4G�Ă9�7�M~�}�IG�I<&n��6v$c�I.$��>��"W��>���O]��M�۷��9F�t�ͻ_:4w��S��R��������TBu�\��QY�'�8�V�$�|-T{U��Ǡ8
NJ%��|k*�r��ǳ��U$���������Q䲎�5�$�o,�L(1�f�iA[СTs,���B���˂����3yr�Q��\���.�[#O�V��Pv��Y�`Έ6e��9Xԣ�||s۲{���٢8T�b�f�BpN3$��v�{����S�* �/�Ħ������b��`-�.UM�q'�+��<����:���<܌<�����6�[�7X'�+�}o(�{�XE~�wk#�_��&���fϩ�颟	n�AR����Zqd55�m�; � u1lD\�}��Z�{��n�4��iǙb�ސy�Ԋ���N�wㄸ��kBX!r!����J�
O}���d��\�p�,|JZ�=Ԗ�� �~���c���_-��3b��5X���T~\v�_r�q$��%,�.�k��i��Cˉ���r@�}�^����i�eQIQ�/H�����d�ܨ#��f}��ۻF����ѫ�s���Y-�B��o����u��Lq2A�+]��J[�+��ԚuW+�)�,tm�石2!Nb��yŰ���8_dێ��840zE��f����PI��~`�V?Nԅ�/�!=�Ƭ�~����.Y#�+����}��P�I�Ub����5S+�W���z�h�EU+��3����:R��BB��*?�ؔzd�>�U��{�&��Y!��m�p��1�ɳ�,�=�F��3:�?�;���X���7�]���P�Y�FP�C���h�A^��K?�l����g�Xm(�DE�%S��e��TDI�G5�~p����A�	��e(�°�e^y�Z����FZ�<��8�Ee|AT�#�||6�� а�x8��wx�PZ�W�"P@TB@JhB���~��z���E���%D�	�C��X�)�S�[X�Q�;�aP��)s38�HN�����z����&jbNX�,��ɷ����*Q]c.�`I,�W����+�Ϧ�l��}Ϗ/K+D\ą����{׶&�ͽզY[�5|�.��j~�&��V �	w�¯Q��Q��9�Z�
���W���݆4��3�����G��2�؏�^$��ݵ�E�a����h�N�d�~ҵŮT.��FI�!��2�1�6��bCP�KQ[��'X7Q���s������e1�7�۵zB@�a{�!�j�q�M��o��2ާI+���i�dT<W�؅�l�@�@M���:A<����E����d�<�eN���`����,������c�d8P���N}
��'���k�%Ƃ��}n;Ey[q�w-ELa�8`�o���<e�fIT�����out�b�,zMѩ	IϹ����v�э��tl _��3`�Ĥ��D˖���+f�/�߬��`T���V1a�p+#�Co����,�K���yȶ�������ˆ��h��qo�*WS�l�*����7*2g�
�Hm������轈U��	5��@�Ͱz�ś-ۜ���W���:�5�K�h��zhQ~Ry(�6p�!.�z��XVw��5Wŀxv�,o��le.����Ĕ���{��'r��3(��h��`K	�&��Q3&����}�Զ�+�0۵A*��$%q7��uS����N��r�xjӗ��	0u�þ���v�EDAA�PK�$`��\��m>C�$�f��5S�ی�}����H�����k�k�p	����3�+�etj0S<�w������h�IPnn�v�Z��Ru�g�3
�dt�Z�\n��e��~ycW<���9c��_hN�X]�Z?��e�� I+��ї	A�������(��g�!�V|������C�����؊4ܬ�UZ����=8L�P"n�B�7�~�g&���]Zd���k��R����fōr�֗����$邞�T0B�=�9s^����r�(B�X�GohS��<�+��s)�mA��*���b�����\�rl��~^�#���Z��A���Ě�Z�t>tD��Q��Y���T�l�uI��7���.�	F�bF�2^v)�Y
�#�e��3�/[�q9��؋��7)=�R��[�"�	�df'!.>Xw,5"d��+�6.;��������~g�F�n�$��ʁb��v��n�_�ݡ�#Y��d��Ue���SSj��繯�t�(�ø;��(᦮|�!���\����9��#�q�����*-r�ܡ�|�
=��R���u\r�,o��Ԭoz_��C7�ϒ��;��h�^��� ���c$hrwT��ÿthB�ϓ����Y�Rh�MW3�wgn.r��N�
ס��Y��9Gk�fޕ5����Q����T�`a�@P�go����ƌVҙ�l~�zV2�_��R�q�#ި�h��-�G�,#���!�L1g򶳎��trg�z�T�֢c\�i�H�?I�暾�a؉%��S��=>�**��g�5Q��q5���RY��߿ ��Bz0"�<f3$9"_�M6�G%�i��9| ����\(�@�z��b{�o��?�N�i�oֹ�_��ئMb>����$�Tu�jk�Jε�թz*���@����>(3(8��XJNI��Aݠ~�o�,�1!b��״���VV�d��6��b-�L�r��9���t�C�WO𪃪�R�.�,Y�<<��Zퟝ-f�#��>T�G?6H��!�Z��w�⤒�����)]ӡR�C!��X0"�(�JޗYy�7�qq_�}
H��QK=7��E ��r�&�\�#	��#�g�	���֋�K'h���̔�5D��p�Y��]���VU��V
t�u����=�NM��uѡ�憜��m����(<?$�4}1���V �<���HK2�\/!_�_�:TZ* ��nʔ�U����^vݡ)�Y�oƑ�ڌ�J܈yç Z\�e���vj�Q�ӉE��=��y�9C9�Њ��Y��.���f��J���K�`�Ó��La�~�ze����sz�rW�����|l�o�^���L�����	���[Zc���b�4dP ���-yKlUq��;������}�ֳ�q��a�(Y�@6wus*������r{l����c����<�O ��.`"�H�������L>��@y���L�_�*f!zD�<yA���.�o�Q�rg�t(P��PF��?�4m(���҂�z��pY�'�G}��s;����s
y �.���VK>«e������U�|d��Q��0� �iϗ�`�*H1�7璏��\m���t��r�
24ʳR��(ef�n��E��v�
������.S9����y�T���o� "ڃX�t'��wX����^�Q���E���)E���S:(��߶	�󓗻�NUNH��z�aa��OZ����R�	t6pj��/���5��*�x�|�Z����d�L�����FkDn~��'n
!F������k�"�`tr�FA�3Z���̿�b�����(���g��S��~���0_��{�s�AH�����?��u-�=(��9> ������ۆ�O�2��b	ӜO������Ok��@������m���l���њJ]K�_X�A�m�SR&2`Mq4���O4K%h���`/>���T���n�3�Y������#uHGQ�}J��j�gP�4��&�Z�ݕ�����ݳ�Z~W���H,��6��p�)����`�!&���#�w��x~v�p(t�k�6V!���q��h*��0O�#�[	}r5L�2��tC�������a��:�ﯣ�	.I�1���@�m|�{�1A4V'^�ذa�-Ao��AFߦ�y������㍏���Μq��T��lU`KFaSl�ʅ��:7zcF���J���é�I\��@�j|��.B����T1�O����%%T���à3�8NQE�x�[��8�b��P�y�p�Z\yP�6��DQ�I��g�RXtD:Y�h�{�AP��˄�᪭N$��^֤�0Šԧ�E��&��'	�U ���=�eo�TC��s�ĉ��y'�aG�Q./�͎��=_�M:<)�E7���3���;vB	�A�6é#l����{a��aE?�e�2����j&:�6j�7�����P��!�M��C���ik�������;�q��V[�6����o�JT,o�D�#��g�:���ᆼ��K�f�5�Cܴ�����HjW$��#fn^μF%��+�O,�>�at�q�D7������=a[��+X�q���f��:��75��Z6���Z�j2\�b���,:�L<�o�y�n��m�5c��ák2�O���D�~�Ѿ4��aV�c��lD�53Y#�+->z�ޚ�m�ք�(*�
d�l6����IKj�[�$��Rv`L��-\���m�m�Hj�3��Vg6]�Ii���� It��."�D������*����I�q� [��s��c�g�r�!֡SN� ��է1��w�@���em�������=��~�H�֣�=����|�r�;2(�JGB��HO�Xd}3b�yR�RW��e�j���$�Mn�]��q��RZOP0�brfC�RBC�}�((|l��,�a��E8`'ß��,l%F�N#���h�<���Q���HG��+�|�Y\T�6�c�:1�(a$Ul��G@�2�ֵs���W�= �CL��/�F M�Y5~�%��k6�B�5�5�v���S�{����D^�C�8��:���b%P���{x�7�sR�eύ�J?����.sjVatv��	j>�CL;M �~�����n�8�	U4wܙݕǶ,�G�1�L2�	X�u��n2�������{��)����` ��#�'������	�8nz��B�̀CC�>�GH���Q@(�e�D�:�(3��h� A)r��~�����8r�H���T(}q����~�ǎӖ%�Ƚ��V�r�c��@��2�$R)��<����qN�r�Q���R�Mk$��	�ڪ
�a7��K~k{�Kk�'�z����;2R`Wg�cl�,,?���t�F���>s�O7�N���O�D}u���#Z�d�p��j�\��vcg:�'-��F�'�@NѴ=��.�n(�ْ櫰�
�s�J%��9����&�^rN2�o�'�A8U��%e-I#��� �E�?ܿ��ߒ�O��=St����tb(��K��LX���S���A�`���:`7 ��J�����lz�: J�N����B��*s"��Idl{C��ʛ���%<���&௅����`�#,\�����I>i��z��<��T�����1^$�H[��K���n%����?�J�K�%P��҉ڲ;�Xϖ�N��u<ZY��$�W1&d�Q�ԕ;����������3�_���������ܜK����o���P�r��c�NU��w���Pq�7��ƣ-$�U��)%,�a�krV���P����}��u���'���R�٥~3o<�P�5�6�.�5IE�Jk��}�|U�uq�����2�+ʄ���,�	�i�Ѡw9�9l�v�v#9"3ia��`א���	���X���!���QX4�lNj��d>U��-F�(�n�܉�s�dO��y��=Q������4�l��G��I_�o�\P��|8b��lM���]V��c��w:�1�N��wE�T0�}#H��;��N?~�"�U��\�J3�>$�G��f� -QP捱�#E������g��ul�9
���HL���ۮ���((T�z�u��&�ps� ��^�+�d�T1E�/:g7���l�� ��z�_�lNeX�z�t���%εr���%ϻ#�#��,y��4XB����I���.ƚ'(����pג�"�\�Kkv˜��4W���ѱD����:�ۭ%��֋��_�����n�l"��H�� f��l��i�@���w�������m0��r�	uE����5)�����k?�Mҷ�-����ڨ��K���+�P%<s׳�*Vu�f����`_��B���A)�M�\�����'M�R6��0=z%D� nIe�a;�N�0��D:꠫�6���
²-��_�?qӻ?�IL�����-(Kj��S�}��MD��Mf�Y$���m��� ��쩡��PƋ4�J��Щ�xev֜��~ܚ��W��O8�����Y�M�GB�t�ģ�ө�;˅�ɏɁ^��j㴪,��L�ay�
tP�+v��o����l�X���}���꿭P���*3�λ3�7m�2(�⚉("�!�Hdo���EVx�H��a��w�q�o�)�)}45#Y��k�����1��+DMe\20U�5y÷������'h��L�m.�V�H�J��JxJq*(�M�S�p��}�;�|]%�ee�M4х ʷ<�V�O�֏ T���v_�����E�%�t���NȏҰ�u#_�;�ʞ��Z=�Bp�S��yi3�<j��l~|�2�c�5�Zo=�/-3��Hî��z���F�pkSη�ن�	�0�`���!eM�d���������@�L�&������7FI�ꨏ�ʲ+Eʟ���Dg��_����/k ����<��Ր�C��I�ζ>�r�ؠ:^�+�߉t&)�`'��ɡ�G7�r$�v_z �2^�j���[�G5�S��ގX��)0z;4��-��Ls�f��23ƒ�ہg�ʶ��u	����z�ऀ���L#��QJ/ʳ� DE�s�H�I����ޝ7&W�Qhe'�L'q�./���˩��_��q��������2����̅�(�z2Jm=~������}Ri�#��"Fi#��ȍs�F�;�z���"��D �\X[�Aٷ0uV�M&m
p���:0�f��^؈P؎���_2�.*����s@�w��߾ͦ�`Oԝ�?V^�3�@��W�f6��I�?���j�?Xe3qN��`��tbi%DG@�
��>��W~o���7�q��-�)�n�19юuf����y�}�_�f+eR��Ђ�D���^D��SG�ь ^u*J���h�;� ��j( �αY^��8���&u�x��G���$&����9^sP��v+���l�a��\t cs;
�-T��VEO��g���!�7�lً�˟S@G�톚�*��:�@�e{Ci��o8��-lWɦ'�d�1����e6�g����G^�l��էrV	��Xs���E�(�ľ�s�T�(��4$AF�����%N�G<�7�����2ǩ\4N�:�Zd��1�bB��BF����9@�O�zR2�\�z����i�wԉ������{���A�?�?��N#ᓫr�1�!pc�:����ʱsu!�������ӾeJ���sR������wh*O9�M�g��'��ؿh1~���DY;�m��x>{А�V����xu�?3`�E�j��\S�F�D#<iBj6�>�9,T�[aV���Eyz������S-$�=Gʫ@M+M�YV�o�*�D,6[�B~��͒`옎s+�����YS��m]}���y� ��!��f��I\j�������h���^n��g����<�_�DG:�����/��^﷬�����Lݜ=L�
 m�{�G�����$6����
|.���?Ϗ�<H�����ڱj�IL3Q�H�������{�0d�}�C?�E�D��%����t����#��u�����$3X8�4�t��D���u��_�{O��K���۵�ŵ�T*J+�qV�1-*C��֤s��ݻY����w�Tzɼ8��G�o��c]m=�Bc���@�l0P�]#�R�fW`�I�0l=3���n*�hu�=���=O%��h�%�V|�(�#�!;̫3�~�Sj\�n�:�~3������+�d�e�%��?x��/=�=e��p��n�|�'��ZC]R<�y�S�.�H=ǐUy��S�&���t('�Q�Ɠ�?����%d����
��P�I�-u/�H�R/�`V�;AG����ȁ�������yhl6�)�ϐ|���v�e��g.瘉��iZɥ�Vz�Ŋ!`F�'���c�ow��BS\�,W����ֲY)f�K���;���f�	�	�`�`�2&��G�FQ�L��p��}�?TBm���eO�*�v�i�����Xv$���v���]�z ������z�EW?�m;M#�@�n��"z���jX4��]Z����UKͳ�����?#�`�:�����-���ZQ�sgصffi#�Cl5�ШLr�]���]et�"��.w$�� ���9�B��w�49+1m\H
����N��t���H��IQf���z)�Q_���\\�KES�|�Qj��Jp(f�K�T�,��0����C�^z�=����}=�+8����pn]��a#��/�౞66��^���=��@� @;�3|y͵��ံp�-������۹�����O����F��)@�H�&1��a�Vzذ��l]p`�z�ry�
 ��V#C;H'=��=��]�_�<i����o�J�Ս���Y������ɖ|�5�R��u��g���?�HnT�C)���%������'�Q��`����l{�/|�B�;�4���)��J��Sq��W�A���Z\D�b�!k���|y����5��������F9��1pj��5_�V,�4�������
�C&������ֹ|�q7)�4��P���kqY��`�C������I�-�jk��)�#Y)�{�W�-L�*���=G�'�6(����?q\��=q�O�4a���NKǜ�I�.DGY�`o��0��N1y<�̮��A*��jH��"����n�u��	�J;���
�Gw����e��∘����)��|	��HD�]�5�A��q��v���@��ճ~�PM�)��G[V��=�i���?��R;�ӗGً�VO��>�!x��Z ��g3�G~�hD�Y�6&���S3&΂�6��G�+"Bw��ʍ[jg��3{�k�/�C(}�CL��� I�a��O�G�xa^jr���M����<l��8�c���
F��ʅ�!!��$pga^� +e(Z� ��vuB�#����������-�i��Q��<����)�S�d=�Y4�*���Zh<o"��y󲚘���>6K�!�'Iۛ%�<�g��r����X���e╄*{�2����M�s+kG���1�C�	�72�Z��Q�/�[���=�v����J��׿�v���p6���=�Z��-�I��LϿe[>��a���ʽa-�Hf��-"{����m�d��*sV��M�g` 2Y�jrdW!gP ��ִ�W��$�ly3�� e.�x�U�L6�8��jSK6O�1�_�p�x4��֗T���F�d�����&m���y�6K_^w���a?�>�o�p��4�NZe��4X��H�a�Z>�`&�+�Q�G�cߐYO����MU�����U�B�el����q�!3K��-p� ^rN�7�����n���������vR�ȡPөm@VI�j[�A��{�أ�B�M����=�#����Yv�5���8US�PT�H��g��7-�v�Zz�s�YdBtx�����º���.Γ��+B��Ӫ�i���+�c+OxL!����O�V�bd�N�`f�p�cs�(�,GTm�C�E����1���"�`��t��He]����2��Տ���ģ-���������?���,���q���i!�7�H@u �z���iʯ��E�#�Vx�}��yz��h����N�4�ۼ���g��F�\jS�׼V�J^���X
G�q�-������iX��?6�H[ h�_�R���2%�f{�HlЊ]�l� KNZ��9'�Y��HO��8M��òH�ɯ�ˁ�*,�B��|���+�]ܴ���"`ǐ*��|՗3�ܹ=�m?f������@��^����	��&o\c��@�P�U�:i�Dv��t�ք��m�#��z����\����z��5���#�e�:��t������{@��a�Q�v�^�]��8�$�4�R����P���ԕY::�Sp?.^�!#D <��6����G���O�t�ݮk�n���C�׍�&�oi�_�~�z���u��:I���Q��C�HW_�e��1)?�.ځ�/z]��d;#.
��IqCk�մ��/����ڥ��L��1��a�J��j�q���洣7j���vUp;l����#����Pz���?���ͦ�
 Zz�����.��\"�����E4ӥ���i�y��Q���y5xA�w�ŉE��2�Qy>�W� ���KO��R9'%�B)�U@��kԊ�����K�YuW*���O.+���}�m��J�3���?.�_���8�W�?S���j�gxL�7���O��(a��9�/�9V��%���瘴n�O��*��1���S��[���+Y>���\�i�贝'J���� c3{�^�p�ĸ���"����q��������]���ܩ����  ��Y��_Z4�v˿��'��v�ᘌ�����6�H�rMB���/���&��7>���/���ske(��٢��$���H�rw��X�/|�s�i�����@�O|�=2�I�Y�-��`�|�b����K�p3�0�,p��
���b������	�#RD�jC��E��mR������<\��>�7�������N��ط�&q?n�����5�2����~:��U���JB,��%e[f�j�x�� �Ǚ�u�=%,�.l�= �_vpM�a���i��q����Ֆ�	)Ç��H
!�ט1F����Z&�&�L�cI���XI��v��U��a�Ue���d�x�� ���#��`��mZ+ڃSM��*܅��EËV��S4�����Fė,z�}� h�S���[yku �}��pO�p4�Hz�j�7��I��MLoE�g�SSN��s[���-��d��$�2��eB����ig���-(�Qe�k�YWu��2���+����oF�!�&�Lp�BE�瀔��0L`����\�=!�K�_��Ķ�Q0��H�퇤gN��ي��C�c�"V��Y"���� g�S�9Ӛ�*I��p��ID������6Y^����*iAuy`a��!�-P���,/�-4���Ƚ;���{z���*�!Z&;���Z�_3�Ͱa<�8��#��{��,�+uMDR9A�_�3R�n�w��xe�x��)���=�Ε����b�1�x�Z��ҡ��8m��]R���g^�X��)t�Z2*��x�M�33X��H��l�C`�֭
����x���7�x��������\]�C��{�S.��Oمm�-�%NU;�����!դr� �K���	}{/��oIGkǆ�K��i�r�����2�~<�U���-�;�B����[޼�$���`��f	���.�%"��Z=�/�8N�����7Hgӑ��}�X/ğ��$e��Q��ـa&�0�Q��|�8�o9�~ ^(g:�QCe8H�qι��ϟ0ȩ��O�&�Ϭ��p�kf����m�ޢ�Z�XI���,ӓ�iʭ��-��RP4���}�q��X-�G-�!Ǵ�g~���H�o�m�՜u�*��T��$��|	�c
�QY�u#�����(r�Eّ��|2�.���p��	X ��^�a�GI8�u	H� o]Qv��XG�3�w>�ّհ�Fݦ�
O�DğrN�q1r�| �g͵���Zi�e,�&G\��T\r��ȻDJ���*'�t�eq\�j� ���J���!�`h7�#��q��� �Z�>CLV�	�#X^��E��|������*�����#y1��C��ɤ�IYt��HL�3MX���7�ˉQT�Ԉ���j���.�b���y�����ui�.��W���jR�vO"��~�&��ɪ*��G�M��9!o8�[R�!�Z�i9]����f%ܷC������8j�K��X�"�ӪEQj���~w�V`[�6�>	��L\ަ�0�}4_^(��)�U�D�M�8v*�(��簤#�4��x/�Fd�<�H�� jS�Ӈ�<e��h"�&���{_a�2�Mt``F�,�D�hW�@K���c���Ql$�V�����&<N�4��?��T��qd��0��)m�e9��bɚkQ,`>ϣ~w
���fϲ��`hT���,��bU~H����-�?2��6����6 Dj�Q�d;i"����	";��)�s;�H�t�!��e��*��-��uT�k�f�C�*v��[����A�}_M��fB�ߢnə�Z�����V]y��d����[�r�o������r��G!�5�8����`te�~����:����eS��ZмB�ߥ���p[��H�`���?�y�=�KT�e_Ћ�|޳@���"Hv^����%3;�)�(�A�7����ڥ��]���k�_;�_�E:�kԤ����PU��x��%H��5���q�x�Mm>@w�"O �x����b^0����ARU��l��J��%K��^3-G,V��g�s;&�]���{Q��y#���4�.�>�B�:�H��2�m�j�����.��j�]�5n����~���U�K���=â�x:���O_��w5�k������;2�Ιh����X�B��4ӥ�"��scN��t*@�j��,{��j*>b@���}t���O
����Iϙ����P@��ed���˃L���]���Ky	b��X����r�����Fu��h;s�H��I�dH�5��˲�r9q-!����������b�U��|ԓ_

�(4E-�z������,���e��L��*"x �\��c���2A�%nomԞb��s�,Y�aJ�'�� �]�Z�ʈ���/N�o�wy�-=�ËyeR5�̋1���x7�ȕ�4`��cNo&h�;eе�p������w��6u�� e���>���I�Z�;��
�X���a1��;R�HV#>ֶ��SD�~, ��u�^D��+�]���~�JzzG		�^}/^�=kt*c�o�|1�i=�1���B}P�d�P {�Pౙ��4�x�::�;ҏ�k����u1��F�,[M����8�		�~R>"D#z<���R�.��_�T�� q��q&�En	Yꗛ�MO�$��y���ӷ��L=���<k�7В[!YT ��Wa��ְSǲڗ�B�!GY��ڜK~�Amm>L2db��\Z���������t���=B���4ɒ%��P�ٜ�]$f�>� �Ϩ��?͞�·��,�b�v��|�tt[[ѧ�J������P����!z������W�,�n�o]u%P�N��%�)��YnI����z���MI�c Zynj�^�x3{�d"�R�pؤ�:U���Y1%�: ��O%IU.�z=Jm-B[6�$?ǫ��/nz�.���To�5��T� 5���by���͋��͡ѿ�bDX�a��ƌp�H;y��8t~�^�dK��eֻ>������n4�V+���2�{<�0&�������,����*Rk�(pXlN	��I�ֻe�
X����@���pN�v p���Ny�l|������Yc�ߑ���M�&�[&��A����m�FG��*RJ�U�B.b��'������F]ʕ#'/
�zQL�PE��:UF���MF��be���=�A���Y �r��B<3�}�Igd�~�.Y���}C��sa.�5����b�+W���7����g�H��P��z��������{M�GMs2�,��@Pz�-�U�!w�L�1(b�_T�x ��U5�t7���6���q=R�ĩ6XL�0-�-2o�7O穏v(	����u��U�oxE{I�^�Z�:��F'M}��(h���*�s���aBĉm�F@~@2���8d�)�|Mg���3J������!�u7��]g��'ߒ��
�\��u���S/��%��|��9H���3bl�[̙�8{��DFo�� %�m�p��?~���m�K{����CcG��,��8���a��ƺ���g5�R�
�I����f�/�~.��?2?L<�"^o5���f/�jV�	���&��&��n5��9[9c�89�9g�L� �5cD�dҦu�x,ֿ
����)ͦ2�y����	k�)�����4�{��Z��=A����(ڟ$؝��A�+���/ɯS&���+�b{�CƑ�+J�S����)���V���mR𧺅�1�m��=J�A��k~�:,'�T�#k�u=� ��g�=�>T�pPn0Dt�r ��X!$��GN#�$��{�7&���O��T_�UP�D�mτ�}3���i��"Tw٦�x09;��TN`�)K[�#+��ᵭ�$�Y��[R�$|�
{�L�7�mNҧ	/�-��d��1��sU���U$���}�0���N��5�r�c	�S��J������kf71mt%�'�� 
\�3�#�����6�Xu� 4^�3Sj�8y�%ӡ�������N�d���e���6�A�.�]�/;�9;# ���gm&�O]�U��vK�ڻXt��҂���0��˗32���/O�����¥� Mճ.���M<G�@��>����6���3Chk���]P�E�n����& �GQ�P�τ�A�\z�O�J�a�BEra�� ���33nP�.%YXe)�5�U����~gm?����z~��ѥ�5����f����i ~|{(�3SvI��H|H���G�XɭƧ�(�u2��g�>d�2\�{*�K������l�;#.4[��f�uI��f��L!95^�v=G9������XU�~*D5B����-��e���E)���?�ᔖ�#~Ś�TP���J�_���r:�cz�>� M��~S�D���|&.�}~v��@:;y��E�����5A]*�*���sѱx�O#&==*�'Ͷ�>�#�V��Y�=(�Į�O�`�����o�\٭We#z���R3��Snx��cGVZ�G#��lC�Ǚ��������r��o�=(P�g�A�<A���Q��O�|�xO��.z7�z4��:��{M�K��`��nCj	g�y��#�r����d5#,0�jH5>�z����>��s��x3p��� �@�ъ����ϟ���e�g0Y�Ɓ��Ǘ�<^U�K\�G�����<H0�:��I�n�~o(I��~
/߉�jf�3J�Z}�5;���j��Tٝ�;�c5u���'*��ʹm=("���hD`#�:O1�=�S��=cc=
�����Qp�;��O}�m��Q�D|ˀ���'�n8<����jت�X?��V�z���C`�W��l��H{�c���R;�c��腷�,��,��#���: ��Z.����/��>�� ���^Pk�g_�sE������!�_9�V!8Ȫ<�Y"z��i�����G�\���B���#C!|��zj%�ջb�>�����@އ_Y�%׈sL��%���4UP�r����ݤIt�$^�����mfN� � ��Q�T��[V$7��E��[���B��>���5.����d:�y���
�Μ�H����i��Ƃォ���5����*m>�_@��n��À��t��OB�̗�w�;��c���:��b�T���/*����ш1�����P-Br���<�m���f�B��!"���e�:l��7eh����\��ṃ��V!���H�N�	�A�!��,8+o�J!�Y�Ͷɤ�vX�XE�Q��1����̱ذ<.�:�/5:٦��%^���!�de�^���˰SG��L�\W���]s�~����"B�b(
ˋz�Qǵ��	]b�x�P�n
��� �5/��m�b9ú!���~�x�	��Kz�w�A� ����M��G�gG�H�m6tBŕ$�A���,���hnB��J�#����ms�)̫ʦ
3l��_���1h2��,������i�)t��J���/y��"S��Q"'E\���r�+��t���n��"������lx5 �DJ�J>��#q�~� �}nQ������x*sv'F�t��N�g�foR$�ZY/y}�^|r���6U��������</?X��"�ʭ?нx<��2!�߈����a��a�ZNb%E�R���&3J���t�sT��5i�O�����okgM�r�b
�ퟀ�x�� ؆S�{k���H��4w\���cw@<���ii
����q^6c��/_V��i�Y2$t��rC����uu��$^C�M��v��ߖƼ���{ߌ��� �쮦Xk� �?3�u"�-}=#�ſ'����&���q^}����b���SOn���@K0�E��}
�{-Ua�H��Y���F���G=�\��V��T�\@W�g$(2�'"��Lb��oeL���E��bw��,#����c�v�>��šG���C�7���`3<���_��O*s�:RO��،G�5J!:�$ZjA�%p�X��rԥ��B\jb�Ug?|�?������u�E����.-��zN�c���BW�[-�k�~�W7-��r��Y�;�*Fk���l�������?%��Ľ��	5��ѱA�Z�0s;ܶ-_\�	���u�<#���K�6��S\=	%���]}�A`���,J���`D�.Z��y�qN��i��Ǩh�V���`����m�Ś= Y<�.�1�q�/��~T���v77J��zK����<�_�>�m��}Ծ��)r��Ap��O��)>z�$b�=�Z&�5Y�.4nS-?���݃!�&�m`�q�tjt�N/�\���fΎ�I�v�X��myt؜M�����q�{��@��U5ET�]%l�ުk�̠��-�tH6�j�N�_$٫_�k��tp`����� �k|��91�L�O8�/��Wa�+l�=^��!H[��--
��������|��7���$6�bX�����=��F��Iw0*{wV���&��n�X�W��A?z�����k����FUn�D�ڑv�`�i��M���,�0ˠ|����;�x���{߆�XvZ���`7qX���4j+QqQ/��ᓺ�]f���.M�� IdyMZ��������wn$�9��8j7����M�_0��R��0�{�;����Q5�Z���75h �5R�O�1���P_S���!i�oXO쪀O����4����N�"%iB�BK�O�]��8�L�3�D�"�����->�~G���(��g8]�_}�f���Ʋ�/��	�a��/���	4ja�Uy��V��W��!T6Dwh4x^�p��y^���H�Eƚ�_һ���MGG<�p��I���10x߾{y�kKV>�j\�%���<��4R��_!<�1n���۞�>�aTQ�i���?���\H�I���~�d���w}�)e�*K[�����:�Ȅ3��ݜ94��M��Ԙ�o�pr0�I�AY�Gs3��5YQK2s-�c��h[��Wo8��MT�7.?$xA��6l�2�c�b]�� "���!t�y��5�^�dh׵ EU�f@Y[M�����o�!��je[����rX�g[5z[�u7cwG�s��\>3�Q�g���bbM��[nzPW���pBa�LJAS_�������
�>�S^�� X������Z���A(}dø/- D(�L�RU��$}��K/ݼ��'���^�>�̓��@�/��PX1��)#�7Y�諅/��e�Yd�]®XT���
$0���4����x�t�ߌ@�͊F>@2�J9D{���S��H�3zD'wTBK	!�)[O��eb���`���s���8�2w��l&�$4�!�t��5��0��\�胳�4�xwy���
"�2��Ql1N�E��>Q�z{=k\�i���ة*<wq���=o;ˉ���Ի�^)-�xx�ʨ%8����5����U�]�b	���i�����M��=*Ǭ�A/���9�SD��;�� �`�V��pc��;�k"����o������T��6��[��e�J�}�?�������/
��͎b��<�Fz8�~��v��rJ�(e��\�R��r���8/.��k\�G��#^�=NL"�M�4������퐑�]�"��}ܘ���	���$4i K��V�Bcfm�:�|p'�G��ONj����ts������]}�Sكp�%Ń��!�{�L18����&^zk���\��\A]�]��i	9A��SC�$Ra���񞝽����u�H��MۘL��LR�>��l�Q�A�8��xk�E`�j}_��Io��~�P�SK�Zf��>DgfS�b��o<|�H�"yZɧ��Iͫnx�xHIF ����ԟĆOV����CbH��Jx�S/��a[��j���ej��1�&Y���d'aͯ�)c��k�ăβ��zk#�:Q���� �>9��!����v����_���s��	�Fm q��H����esU�ծ��}ŝ��9��� �\1c�T��������`��:�G��fd#xۏ0��;qAR�נ0:J��/���8�j�����}�j�̫�b�#:�5�b�_j)*�X+M��|j���\�Gp{Ǜ䣶���<��� �����.=EMѫ��/��0ܱ�
�ޮr�6h}Bh	��T���][�|%)�됲��~�_B�	~�H@�4�	k��U�Ѝ �9(z;8�p;���{��p����ĉ2{�~�Q�߄���{��f�X�L�PW����: \�G(j�L&j��5��2N�DЕK�$i�M�l/��?��PĄ�9Ѭ�0"��x
k*)I3v�ͪ�5�&M@�6��|�j�X�`)��ll������-�wR��3�)��{P�o�F��t�E����{ٲ5�/�ϗ��3ZH�*�k]�fbԕ/ف���.��Ho��oN�zPʖ��_9��M�J��� ˑð�g��H��ñ�%�盃m�c�ٛhWЩ~�� �n3�	6U���n) ��p�R�d�̅�T當Y����r����N�2(��AT� ��&��r����#�� h�����B��zc)p�1�r/��qs�����\˒�Ս
6o/�W4�%Z1��BY��Vl���F~�ul�@[�F,	G�f#��H1 �@k:1C���i�/����m�u<�hϣ^��*Oc��5Kk���Z���b�w��P$����^�fg�^�����(EPl�-dh�Cw	�$vpٽe����vMѭ/+���|��̊B; C/
l#>��g��`�,q4O��R,>���/��"�ﭩ���q�l~��ӌ�Z<�x�8���f~"��QQ2Q��\Ç�#d4W~H�8=�w��ېC�}D�; u��T>�
���Hn�m~u���hw�@��sT�pK�E��?t���H ?^u\�2������Jք�����H�I�9�h�(F�}Z�C��T�O���#�#?	\�� }��zG��)��!��,�#�gN��X[������a#���h�"s��.a�ӰɉR'�L^���>!�H��Ӹ��Zz�a��#�1(��>�ty��R�F}�A�H� � �FO�˲��NJ��+�s���=��:�eE�j��m�Q��[��h0�E2�t��/t,���~���/�W��5~~r��b�?^7���q��*p?n�ť�@+ס'����@�<��P��Ӷvn�ꇍH}wq8'�&>�gA`���vE7��"KȌ��(�:>F�#h6(��9��L��Ho�-�%�kn���_j���	�%�9SZm�[���WSt�	9��gƔz�h�o�x��ǽbw����7��6,V���T��L�k$�88�v���~ܽaIru�X[����Nzpg�0��L��,_ʮi(x�:�]o%x8V%����y�Vt�BZ5�n�5���WvZ�g&��n3�]>Mə�{�m��,�0;"�&���/J��k���-�&@��!��<�q=�jQ�S:(��	��2�$�A�O!:���L���"<�>�f�� �Z���\[%+zm����eV��K;�6��{#�;
HJ��ѣ�0
���MGW<�5�c���s�8��P���xV~1,����.�hR�� H�<3���hH�p9�� |���I�G�e(Ԑ�z�U���5�:�h�Bا��L��++���UV�)^�!,�-�%(��綍sQGO�C�n���uywWuq���c�0������mn�zGk� y53�[��h�< <4��a3-�n-��_����5��"����������Y `�l0�p��w
�H[(a)���ǻv�G� ��IS�&� � �"}Bz	�&��a����еZsh2g��AG�4:���f2���o�%�yJ�O[w ��_3�!^ ��8VN<����%��(���`�#�ry��߉��a�D�d���� K%���R�?be��>�٭�:��?�Ƣ�C�=3B�[�/��K�-��_�ީd�_ؔ<���������\�BFA��>+5knӝ@ς��>��-�N�	�mI����ڛ6b+{��6��Z�҃��.��RF*8�+z����� ��o)�%�-�zJ��@B,x)0�|�ӿNm�iK�?��3��
�);�P9�O,j"�Lu:��yAI���;�����_�ܼ��6	n�#~�¤n��@��rBt�8I��n.���iib J��BB9cו�������/Ǉ��]E�sC�� ��y�� ��W�;ԁ��$d�s���|�A���B�_A�9�� +ޗ��<����")�Bl��i��	�gL�Ƶ�it���m��Ur�Ѿ��X�KG#��*��+T%�l�W�ԡ�W\#����ǳpIc��|6U��o��-�\O��%���|������l�]�j@z�"��:���/�h�`���zR��B��t�:>VMߦ�Wūo Q�g��F�u��Un���e��M� hd��>��0��m��|~�Ҟ�?�% ��7F��Kr��Ig�Y�|=p�����h2^�8��8���?zΞ�LE|�%W~�>E�țC�Z+M�}I�ղ�^ �F��hbo��1x��6M�������"'�^�0����E�OG�4sB�?W��gA��$]�X8d�A���M/���	�#���dY� �A#2iy�O�m:�᫈P6X�i;jF��Q�Fޢ�k&\�&����I�͇���	�a~��C�)`��o��_����1�2����4=��8+  ���5��j^��!���az�z$a}��H"���'�ţ͌a���+��w���<*]W�<��oU��.5��}��[>J�t�rcN&}Dw�j[cp��?)����4��9��h7�,]w�TZ<�Z�OM�z�B�B�<����!��$��� ޼H�#����u�!"<�s�)Uhd|[H���!C?6#!hZn����%Ǘ�>K�I����`�yP�d�4���<� ,�ƳdD���B����ℐ����%#��˦N��M�4q�)��1+���\Y�O?"�<|Bi�*Ӥ�T���_d�\�S�<�����͸��p������p ��2���\O=��>|��ݓb`91�L?6eK4�7��S�4�%0��z�yf��d�l���GG�ާ�O%TN%]-=�J����vKS�����X�����|�t�rR�^v�do6��5��z�N4:�^�h�(Ժh���ɣ�Ө5��5��Ɓt��Ӎ�,�E�/Ȼ�����=� {�������Xt�i�M6�2��Ú~�W�b�I��>{NI�O]��
�_�B�M�aa�V;�X�y�u"E�pjٞJv:X� ����0�Z�k�3G�ǖ�h�!��z)P��^����wB�oD7Նc�8H[r�5�՘��U�(6 ��1��];23�����5�j��%��2���-��[+������2<[�N
)��^ a�Gw��>�t�'�9����h0P�z}[MnV����h1����G�2�!��/��j���5_w$�i��-1N+�J�f�m���C�C<�w9��W!��)t����g
n�	��0
���i��0A����rů�x��.��&l������V>��5���V����,�h���$��^-�#�����5��x�wMm�O3�%� �@�����8�����Mط�Y��?̕��9�
����'���6ٕ��Ъ(�h��r��?1z`�󏖲�}}Fk<90�ְ1E�|1~�a�oq2�6��0]e�*[DWj��3$�FS����8!�/����8�q��M�i΃����s dE�����&>�Yؙ��)S�2n�S��*�F��􍠸�xLu���Z�Dk@�[�����αb+�­v����A�_���r��	��x뗜�T���_D�S*̉� ��<�����r�п����E��Ѕٍ�yS2$֕Y`Xk�6/�-wd�� ��X�u��/N����,��<y��2���&�Ͼ�a᭏����8�����ڦc�����&�b�.�―�0D{�*��v��H�ލ.����e#�����L��z<�4|%��8HTpL��Y{�E ^����`��˽���dV2�Ou-��h��с�ͮ�%bA�tvg
���o���[���!"�}�&�m�������Ϙ0�7��2�`&�!�*�~i��<l`o�7ꎡލ�qŅ�P�2Tcoo����j��L41���m݃�i��jjI)CCx���/�zf�@��X7���#��Yx�?r���?��
�=O�VE�N�@l�4ۨ�0�����9�=51R����%�]�,��o.��]6y<�����`pi�/��b�a��^^�)�4�y��ڟtP�o�dw�������ZǏ4��s��� �)�a�p��Tj�I�ވ&��v��É�d��x��ɼi�L@�U�[T*�zp�
�jS�R)�9	t��V���z��p;(�NK��0d�ޓ7g�=�Z.a2<�Jr�]I�X R8��0� D��8�m��v�Z�v}�$?�G��a�\H�[2�rߢG $��p�z+{BQ0�έ����j�#&$(�?�鹬k�f���QN "�`�st�	1r59� �����[�=�&�V��d�"������G�Lw�<!i���8I��캗�up��{n�$����F�� x��ˆ���t_@�ϻ�P��ݗ"~=!2mވ�06er�6�II��^�h#��T�G����滄Ԃ�їnq �֝�4MN˨�F���ؾ��A����k�v�Tu}�!m�K�U�֟2O6!�Jd#�yh�C*��pz�C��\�^l�,<i^}q�h����aIF%:E�
	�-�I�ͯ���98���1��rU�Z]��C̕b����/I)�PHa�����Ś�4�}i�pFe�DAݼ���'U��8:�F&r�ܥ�4#5B�����J�@2Cȏ���i.A��3�=�ѻ�^�x��yd���J����(	[�bm_�i���"����S�C�	[\~j=GK6)a�F�4"�"v�G�d`}���rQ������?�!� yK�z�K̪����8mC�q�*�+l�,�����X�c�@�5��1
�|9�vԽhU�h��(��gZ!>�"�����fͶ@��u]S����r�S�k@-uꝩ�&�60%$UT�����qkG5��)DYN�p���RmN"�L|:���e�Y��� �n��yP��r�l��c��|�6�X�'�? ��'�iK,��řP�Rx�.=�@�Ou����TG�K��Wg����,!�*��|qqlV6�!�n��ҋ��x��r^h��i�'�R��O�S�T �ya�[�C`����lKr��[��gn����N��E[��R�;G��%�E����� ���c��{�T���iX�{�$?���|�o5Vg,{z�����]s��͑
�냾��b{ʧ���y�UA�<��?G��/����D�7�+�|)���E���e��U<g�9G��7�|U�,XZS/��JQ�-�w �<�HN��4|YB��H�(
���(#�<�y�i��f��3V��
��+ۙ�x��̓ay��'}���lCD��uQ���tvʄh�,�_Hb�����3At��W�b��d0㪰&���3���7�������Ԩ�4�ê$
�^ͬ<���ف��-z����5{���N鬏*���<�VB��,�u��b����G�����^��B��H���>��mP ����w��(���/���(�1�4��Ԯ�Ŵ���*x�5�g���\�b@y�Q��ad���M*�}��L�Q"E������6T�FG˾�2ϸ�ѕ��/E�q�_���4�ԺIY!w1ub��G�<��)��������.�5�|�U�O�$�pJ��<rL����U�l�U�� ���KLk������� ��.p����J���U��O�fM=8X-�o�Ԁ�+����Ps2pX�[
q�9a��g�Pָܡ���.����osS6�!�?j�H�qL�z���&�Zch��������/I��9 &��0�j������6h��������%��w�g+6N<
�@�`ݺ�Hm���dM�y'_|�$ܤ�?�\zx�R�fK�L�Ne\�'m��"���+c��'������j�2Z�gJ�=){vJ�K��5�٪�s_®���?3P��p���<�ԧ��б�}@F:�ÙK�(ЬD�K��v���x�4�%�ET(<�$�sZ�lo���0:?��d����(��6#�;��M�
5��btp���k�����^A�G�#��TK�WB�m�-c����h� �/�>����!x�;Ǘs��	V!y~�嘜P��ޠ��5u-hg%���՛��ih��fiyi&��&!l����J�w�f�_��َ��_7X;qt��m~�lj��ǿ L�}T���O��А������S� rb���Y�ű2��=����7�w��C>Y�m:�F�.Twְ�^�1j��S'��X_=l
�� v��m�;�w�����V���518���d\����p{/TH��DI��l�Q���`d�ߏw���55��e��-�9Jp�3^^��\_����Td�v���e����J����Y��ᇅ���]-�GG�~;^X�<C��()�.��	i�B,İ����/�8+�]��u��.�6�@璥�LɪQ��
pb�h���@�?zھ
�#,��شǽ����7!�L[�&Eu*��=5�r������ϟY�)L�r} ��R�I�����[�KQ�Z�5�&ҡ﫲���A�֋��g��5����
Y�[&�zWq�Ӳ�H�kWX(����j[�5���G�e8��hIc˸T޴
���"�bsE|�'4�K�F�>��QW���I��:(ϒ(���}S`{���ӱ�cD��^��,�V-�Ŭw��Q�x���ߠ�[�a��W"�۶���̻ZZ��&	"DO���p��ګ�����������ĕ�]�VAC)���@�q����nL{�N��Q
?�ꦿ�i�m���7)��m9�1�����
M��P��0����
;�f,:�4#��LU.�)s��b�����Q)Q��s�s��<+n}�����*3E�ו�+�S8��z^��KX����ui9��J�C���E:�?����"�{�~���ĸ�ұ�I4
0=��2���L��#}>+"��EJ5.��Y�y2%���(��GΖ][ �/̹aM���nɲ��P*I�\��f����eֺ߻��L�2r3~�Rh.[y�������lN�?����y�����+�M]��$?iI�'�T�Y��lUj�ɋ@��4�pە�el;-DO��ۭ�b��_Rh��$l$�t"��m�خ�i����%�;���`޽�4��R2�_�֯�B
��~���$t����L��J����-��7Q��mn|ש�.1.����
ǣ)/�q1��dX�����b�?�����|�V)G��(o!���i�ίy��R	�c#��%y�΅Q摤�1��q�s�lKrE���-��Q�����`
":��딛�<���*�oɨ^������	2C�+� �Q-9��,�ز�S#�d��2 �R�E'Ǆ�@�C����L��_�L:�C+;s¿[�vT^P0j��&L�(,m;�ft�>�Չ) '����i�9��%a0n�nM���ظؿsf}*�����ʗ� �33�|D���Z��r�Z��[-q����Y�����ݧ�`
$a�H#'�J��x����<��i�A��<it��'	pǻ���XK���S��E� va\�f��ȩ��Y���\U:���ߌ�W^�)�����["p�*��,3�l��D���g�w{�����O[Y�i���ޡ��.���^P�6@�(Sܑ{W^>}��:s��@ZN���GHs�?�F�QXv ��PG�:�د?��&ە��w�g�;��gR�i�1��B�u^����o~d᫽���s�To@��+.0� ��C@[��_�!���ٯ@bd*���f�_���m<&�Q��e/��bj^�:��n�]�;��h �8���_U)x��c�P����( i>��;�ou�k�6����Z��p5���Ƌ�r�ʎ씅|�4�n4�X*�:�O�' �v�a׫���ݡ���@�� ��Ge�����4'c�ꎁ.�\#��{꠴���+�2zհ������{���x�	.r���@Svj�x�Y�Y9������5 �ᇱ]�F�9�O��� �;ne^Z�l_���_��ߣ)k永�����r�q�X2p���T&훻��7viA��N��T�L(���S��U�٤avd��R���E˸
�Y�ub�(ҵ�+m�w�X�#��:�����g�'
ߘx���:��M�cXD�Y�%
6�Ac�Jpp
��cz���6��	���|�_�\���KVb�v��D��������/�o�^���|-T=��ͻ!�(*@�.��L�������6��c���9�����b�j=Zc�(���2j��*�?�����v�Kk�<����mO�
�K�!yi���+�y��{���l��.A�����T�q�P&�a���V �6>�a�e�����&쒓��Jm!Pa����YܰIڭl��N?ގ� e#Ġ�3��p4�D[l憏l���n9&��ZO\()�҇�Wiߒʀeix1Z7�x�@6K��^=��B.�O(q�\a;���|ʔ~���a}Gj@�w�%O?��
�Q�G�?� ���ox ����� !�Q���V�c��\�|�3�¼�a�	Q���TX��б��,g
��D��=T}\��G���b�H99�'���R>�Q��ɱB���`� �o��h�eL����Wr������4I��h�j��X����N2��N5��Y@�� �`db������fT�;ľ'���Y�5"�����JXJ/U���ԣ�)���c������er�$R� �C4�)��R=����a��T+�5&ߨ�v{>�ZJ�4S�14l;
�Q:J���d��xq�e]_@�$�A��Y_C}�x_�@��(�K&t���ҍ%�O���ǋr
J���2�2Ke`l.�ڭ'y�}��g��a��`��k?5F�<��hkv�J-�RW�Q�� ��4Sү��������U��cj3
�>|����u��Cg��t�!�h�5+5F�g�/q�"�+�E��(�;U�sf���7�U6�����]*Â%�� F��E�E-���G멿[�Y�ƍA�4���㶊�^9�o7I�#�Ȁ���F���
�C*��V�� ��c�5kP���T�*�O��I_�0��i�)p�2���Z��bSrZ`���Rڗ�"7y��|�D��J����`������~'Lv�V['����^!�jB�*�Cg�x�Z���Sx��O�wp�k`1a����!th�.n,��Tv�R�vy��Q� bL�������lH>���bHow�5��9O߶�38��4�����f����M�Fu	�ΐ��hɜ7�Y��-R���i��y��k"�����7�*����}ϗ
u<]�@J\���*A�EeȬ�9\���D/��\��ҰCz�H���Y���lB�*������H��W�F&zb��
)Jy7�e���g��o���f��
�|�𷾫tvʾ:#���փ0?DéF��|��%�9�ˇ_��
B�ĖR�sb�����4���I�Ԋ�j��$n�(�6����i�I?!�R�a�6g[O����Y��L&,( 4��u��v��qG��� �9�����w��,d���OD;�0N��"	��d![T���4��]����F�H��X���Y6�e�"aG�C���ӣ�$
��<H�7���6�AV�⇤<ʖ���U;������3 ����o�����H�?.�x�w?�\K�)�j&��{�#@/�-O����-?��HtT�	j齎:�	?�U0V���u3�e��ӎ�>R�[�����P��w����~��+	z	�ӓ	�$�ճ:؆����S��\�I M٪�1���`f�	hoM�Bs�qȒAm�	��w]�V�O��)|�F�4�s���Y�t�	���_Aӊ��A��a��J��dO�?���q�
 Q�L�@��u;riMI7�z�5%��o��~�{Љn�5p�X�@�0(�"9C׿s�@\�Ո}�R�7��*����[��t�Ɠ���*$˩�[�d��T�$�N�,���)�&%P$6�6G�B������Eu�P�Rs`�8O: �~6�]Y]�?/W��*�%-F+k.���7d�E!��nW�q�]�(�ᶗ6�kGǋ2^c�f�(?�^�
CϠBE!W�2���j��ȇZ��:�9?�	�r�H6s�d�� O����Oǰ��<��8��5ȸ�"_�y���� eeم�T�ϲ���I�0�����+'��vR��I�Az:Dr3$����Ӿ��I���4��i&Y��oN�Ͳ�𛽥ǀؗ�w�͆�l
��a��\"�y
Ôv/E�(5����)�h�L��.��7g�I�d�����)<h��)�ß�5���L��J!�^�]t�xBH�~�sm�4��H-��M,��j��/~�[��P�^�T�9����P�б��b�$ ����<>���-͎��|�b��>�r%V�<wa��(�LBybo8�P&���Yw"�)4�"9�4c1l�yA>�1��Y��_�:$U�K^�RQK$�_THL���ܯL�-5��ƹ5�!�Oo���[�"25����ۭ���fo���
����W�I/!�=hu�PX�$�(����{t|||���<����@IW�|�R� *�ȇ3�Is�;4M�>٬Od�ϛX�>�b�����(*v�`w��<��M&���;�1�`��+̳��
��:A!ؗ �'>0���.i����ـdܟ�kQV
�<���y��{�]���	b�`Ѹ)Cyh��O�5\Z����w�Wȑ����,�K׼1��E���K��@Q�D&��FK�('�%>!��L5tɠ����5*oWg��W�1&"� 5�Z�x�E�e�Q��	4{[�'b��Y��-�w*����pW��<7A�����1��/;��C�!�4��!��(�����exc'벢�a��B�U��#���}�Deד�� �4�9��^���%[��L0bZ^-C�/�R��a��J�Ep�i���ێMN���JUCи(m0-��"-X�-��&� O-����_�Eu�O�ɛoA�A@}h�Cus�U�%�S�_�����a�Vk]ImZ����$6������y
�'�r�_*Fƚ�B�2x�x��h���ѕ'|�f���P�<�V�}�G�Mn��NZ��a�����d\��N&�ɐu�~{�9��g{J��f����+"0/��1B�a5j�E���:n�A����-|3j��Z�+Ğvi� ��hη$��g�'�27���(dD�0��h�t������K�#io9����_K���02�1�Y�K���Kw9-�4A2�`��z�%Eߚ�T(�R�Ͷ��U�.���|y�Q��p�=%�W{�=F�PH�}�ȷ�}彇.B�g��Ms��k����,��ڑBi�\o�7
��]�1�ˁgj�+�+��9
,ѣ���D���L���AD@ Q��1�1��E+�����^���y�V�ǅ}��H��&����m����Lh0a���_�E���5�WU����\H�����4?pD#.:�,a!+Ⱥ� �Z}�`ٻ�.gA���YM8��RO�"�ap��Pѩ`��?Ѱ���O��ЉG�G_�F>�#��S\2�2K����1��1�X���1�\y�l��O���
����,�O��=zƪ�,����U,���\�R؀�[����?�I�k<�CS8C>㼱Y���d߳���T{b ��p�' ����o�`0�9@���O<M�x��v�Ø�5���1>q���I�R�e��oN��XU�4K�+��r[���5４U(���̩��n�b��p��*�>p"��r�����D�qjXL�����;��;΅��sZ0�Vr�	��S4�
�T�1�Ѹ�%}���
J�l�ä�x^-�Ͳ��̓UcQy��ș�u	Bz)�-U�}�R�o��u�tw��%5��4�]­*橛j9��7�f�W}��V֭�Do�q;��:�n9L$#�����mV(�*�dQ-uD�#@76�FG0+�	;rc��ǐ��U�j[��T�M7�,G��q}��΄>��2�.9k�q�-ހ��s�%�e��+@aj�՜���)���H5��ߗ��T%��a���c��w{`	?��+T�`��9�i�R�ov~=�\ae8�:�AA����.*\��v�T���L�3��L\O�Z�!jx�Q�UlG�.���&m{;����x4�~��י%�+�ה_.����ޓ�s�?[iѢ��q�E��yA���F�v�(n����(_GԔ=�O���F-��q��!z�#ϹF� �����ٓ�s�ѡ�m7���=;ҙ+#�
4���*�c"��c�x쿆�҈¿͢����~�%~�@)+����k�F9��,��s�RbnGv�������>���Ъt��v�a��	�>A5����
��s��р�c99yrW��mtC�
�j��;
�_��$�"k��E��G����QRԳ����O�ax���G-Zg�Y����R�L�,B̾]Ay�Q!F'�7�t3��� Pr\�P��v��L��	Q�;3n7��iV�Poh�V;k)Qy���X�������ml]����%��xU��U!�vj��{_.�hB�r'������.�gM,�h-1YS(��Hr��'���I���g��}����w�B�ю:Xv"��ŇW[:�\���V���g.�Z9���N��-�Ӧ�E��V�y�K�ϕ�� ���T������jB#Ϡ<�62!�<�l,�G>����H4N8�^g9G:�A�E���-8,�x�[%z�=W<6���n�s���������α˚�&���]��n��_�#)��ِ�������������ڡupÓ���F�	��5c���7Ct�b4F���M]4��n�B���TzS��l�d������K���[4����� a�����HNŀ���F��Ɔ��ڶ� ����u'����e9h��$0�3������@���SA��q�lp��bxk2U[ `�~���6.&F��b��|Kx�eB��q}���DP�JC&K[��^g	&�;����{5	S}(c�r$f�IY�
�U���l}�/"��u��6,}�\��H�V5���j��dC�E+\['�`�'���-���l��Ѩ��6k&�����+�8jǦ��� �U��䲤jV�{э�f�_YY0�l �^L_֮�4v��`͚��x�� ﱡJ��K �T���E�a"�"�1�5��eM�fy����_�<���:N	�8�T݄�2D�}M���q[�)���٫&06�ш���p%u�v��7r[|�Ѻ����q���k`�%x�gL�OW�����t�Z�/���(��'u����NkR-Ҿd���a��v���3����k,�밭�p����p�Ҝۭʻ^�����8C����y|�l��d�r������I�m"0}`6b��:�Z��&�������䛙��Qe&���w?@Z885Ek�R� =��dA���1%m��zPd9dQ��z-?�+�sʪZ��+@3<�L����c�j�c�\L�gALDH�~_r��X������r��:Xߖ�p5ڕ�s���u�`����K��ǉ���[������j���X�:����dT���"u>D����p6��jE~VJ�Gj��x+�98�{��{��i@�W(�ci����y�1���W]Л����3�1�3]�������b���T�r$��	~��64���g�~)z�2{8����|�=�-���Q`�2(���;z���೘��y&�H��8��("���2��P��X���B�/JJls<M���	� ���]m�cշ���t5;����$*dZ����6��y��Ď�	�{�ʁ]�m�I�~~m�ζh�>w���J��N�t��~(���I�zf��������[��sWNϻs:{Y6F��[1��x�|�U��]�:���Mu���+�y�����r�v�w^H����9;����5�z�g������Y�%>Uȁ[����8b f��΂S���x�XŃ팭SP��4���
c��'�z����s�n����2�6f	��~{ T�[2��{�I��\Se8q�������K���;.?�T�-�>�_���6Vk��k�lT�Y�w <L��f���&�d����WR�YÂ9<�r+��L)H�Y�H��/��tLe�5U��#���[OoafPͼ� �#l�Y�UM����~l�QV��gb���W�'�!�n��ʝ�*}^����
'��]NjХU� {[NJ9�@l��.�T��WH}qџ�՝1ud���#�sT�(�ب��u��g��z��P��ۥ[w����7��3�G�e�d��-���ז�3�T��~0V� ������䀨�"�]�s�h\�Z�I�<!%Iup�˃]|��0�:Gz!a#�������˝����G�U���s�sEN�����Z�2���J�ǘ����*�7�L�� �	l ���?SgA�d�I�*~�0{\S8�qꤰak������E*��J�:��"tlk6��Da�����z��*��xb�=$�;��럮l��	b��R����U�$� �v4-��n7�͘	}��'UM�(}�
�sDÿʚ1ȶ����Rؕ��D2�.G�*��&J�B?�E�rֵ%��G���y���K��xm��-�o(v˰��ˢ�m�0E��H�f��O䞏ox,���_���t�u�ٞZK|zqv!*P�"��xrY���?&�>5�I��5"_/ɰ��<��d�������D�ͳ|z��:c<�k��r4�6o9��[-��W��Pd�|��-�K�n�)�����d�y�炞��C]�'
��U��{џ�_o�w��;L�7��T�͹�<[��Ob�R"#�%$Q�:�D�)cN���[ݳGo�#q'~ږe
����xP�86�#��^IS*��\�K��e�X�D�]GY���NȰ
�������M�	�@�
,���^�+�]��{/��f�&W��k��VR]����\h4��qJ}�j��^e�/�;�*�:=�P@"����(��M=�񍬰J��MŽ���ď{g����&����'o����`���Ĥ�\���a)�^աU~"*�����1yV��7b��_bE���~��}[L�$�{���3��0+`��������2ը^ <f`�tMġ5s}>6�6O���	[̃���d��
�O�y��k0����'s��x31�N$����3��G���u}�;|,��A� n�J�)GG�aP8iK�׍KܴL����+� �Y�P{����!�21q�{�Z��S9�%i��Ǻ��g���Q'h��l����������Hݨ�y�-J��I�.�G�	1{�'��~5��G��y*�j��a��z�`X�j�ϔ:gM��9#X(����ȧVS����Α��H�&u��A.�RY��4S%�`�>�����5��s�\G<)`����/��ۓ�ny��$�t����Wz� �?(#�?3����+g�ݚ�-��9�Oձ.7���B�	&��,�N���躻yܰQ۟�N�b�8C|��\���-Ҝl��2�6@��v�h*�p-�H/�5������,M �y��Ưa�ᣯe�V�pJ�T��vY�O�d�69
7=#$�cP��3^�%%Y0$ئ��a��*k� ��Ȃ*�����
�߄�@'�����7J���+ӡ�<���!f15[5�?��/O�	��~z�&�`�%9A�{��g;���|�Ŭ��_���ϓ�����O����W5���CΓ�hI��X��.�f7��!�6Άx�8���E�($���לi\7R;�W�P�:��8Hܺ%0���)�����[�E� �c:g�Qt�z8���)/K�U��ݣ���ڦ�nG�Y�F�o�\�R�9���	z*~DP/��65��
�F�k������u�..��������ە5�j{�혇�~#��M&����t�((�������$��k(�F���B�����-Y/�!���[ ���Dɏ�l!�#E����P�Q��N��+X^����6ҐWY�KV����v�m*�(�{vs�>�[��,Pq��͇�|/��>Z_J�&nTj(�a"��J�������rr[=@���Lu�e��p��@�����b�9Wa߯qjK�n8M��g_~X��D��t
���Ab��tC�G��<�mNۦ�k^���~d���1dR)a�XH���hҞ�RĒ~KP�}���in���x'�x��H@;�/�1�k5v���Eψ���1ŞyN���o��;�.__�L3�+�˯��[���zRΗ�:Q�7��|8�Ӹ�"���Ò�W<��)8-X�![�\���h�vC�=�pI ����^\���Ns�\����x�����-��$C���mϘ���1�*W�Y�����"|H@3�ݓ�վ*�)-�Qul��5Pq������z���  TB|�x�G�'���oSj�a�P����p�e��^hyp/��}�tvx�9}U�ٝC �;�������@���&v���y�r�5��꟰+jq���=�tW�	r��)�Q�o0�r�����xH�S�2W�5�n ��K��^z;Ī��H�,��n�8^��T����sݔ�[�!���k����2_щ]�~zL�ې���ܚh�[��k�Ź�sk+si�r�x���R��@���
����et�4�rﬦ^c�l�� $������I�AtN#��K�wNh��~Z'"��p�--�V�f(є/��X�B����������f�-��O����7�(����K��"k'�����p^C@�W]��\�Y�/�%��p�a:5�#��=�(g
!`�VF-T��M;� ��"CuÑ�F�rK�	"�t$��X�R�Wc`b؊gRiUTz�d\*F�#��x��+ilY���:I�ೳ�֫�"(����z���:�`}�m�ā�N$�]��x!�(�f�Pz!:w rc���&�9υ"��N��=��12�al�����h����>����1��Ef���9蟱�	%�W}B�q4����?���	s�����fkio�&(8lJ�hY����5[��S�˙�-*�!�A ����oxp�2��lt��T�zc�L1�O�������h�}Tsn�yM9�9ċ�ic��mhX�u����vݙI�>ǡǨs��=��]�J\�»��NB�LI>�X�J��A~�j"�o���#�ƚ���ʸ���is��r		�� ��r���FIg�xV����?d�s���u'���w�Iz��� ���q�� �S��|�]fT�=(��LQ��}m��h�4���|��COE�U��|�t\z�Fw�I<?׷M�s�Qh�`�������,S��~�*��\�1����An�}�ui�OR4^!r(���W-�n�w3a�W�B��3�&�Aw���=$�p�Y��F��D�J+��;8FD�I2���..����T��X��܏����cl�#���������=%�u��^ןrL���J�wUM�����/1{�c��p�R\_�$BC�H��M�o;,���0��XI���7�ԅ�*�(�5J:6�H_����<@�*���w��ݤ2oW��uK$}�6����]�(^���񊋞�L�)zy�v{^l��씚t�Wɠ	�Юqd��" ��81�X�ï E���飣/j`��0
@K��]�a's���X���̦�k�qN�)O��F��SkY����
�sx���qm�u��k���f�u|K��d[҅vG��7����%�P\@.~��iT�kF�.�(*�����0����铥^�n���oU>��Ⱦ��i��HS�B���ݬ�jf�����6k0�Sŕ����4HB �`PQ�0wd�ts��b��$ط�5�lPB0T�ʘ����|��mr��k;�������&Ƴ
X �d�"�ޡ����LI��p��	�����
�\ }Փ�
߇���m�	��{qn�a�i�`�X�p��'�v���aa��J�����h �B@r�j�M��ۍ""8�)�R�,��*���Rx<�����t��C�o��-�E٦@'�.Gk����@~��̧v���UK�����u�%v���V�X��ٮT��;+gw��M����@]!~�J�n��0�w��%k��ֆ�6G<�30�})�[	È�.e�\�,�K�k��T7�m�W���jRqb���64#�<0���U�.��T[kP�:����Km+d��ȗ�sd)��J��T3����� pLu8e��UT�_�����c_����_2�����t�<5v����YJ+K]zCe�UM� �]##?����e5c0�A�nibIş�gT���8/�}� �́eܾ����:6���)�*u���ԿX�DG�j��k|,����ذv�whC5G3�u� ���Z����-�@�����s�����r#�3�G�3+.�{]�V���t��e1�%�b�J����ϒ���[���(������_8�јIk��%W��wɠ_�`$j嗶��QF�1���_{N�a��`<�S�t��Z����[�2�oћc�%���6y����d�,}�E7��,��o���c3�>�7�*8�����v�TE����5�����s��"}�c�0C&����d��Jс���tV>�m8�I��ƶ�rI����M������r������t��}���"ٟ]XH��q�*�˓�
�	���,��],ױW@�̈2pxVH�U�g�ѹu,3�kD���;�L, <��㶘�.���3��Yְ���R�}x���/k���c�I��*�6x�3K(��Zp3�8b��mu�&T����I'7�֞Lu����[V.|-<~�k�����yY���Řq�݆�}�C�>fԈ��� �E����~���&��>D�j ���!R�>Ɨ\�s*��΄���0��ZyڄӨ�w�:�v�:��Q��5x����?�q+�8����"n���\R�-�l}%D궐�T��jP�"��AR�2`�R�@U �)��Ÿ�
MߒY}bAഒ-,�o�O��5�E)i�u�v��͕ڐ�'�f]`�D����ȧ�	�������,�� m��)�lr�����nshM�8�b�9-�E�ؼ�T����9{F&]�M���Ӷ>ey~���j[d�we^]��ʒ��J�W�6Zy�b �7Q�t�ʤl¸U�v�Q���E�dW��RM{�X0��w_[���dZ�c�������|����Y�Ǽ���i!��+o�mԠ�h�#��{�bA<`31y�����>~�& ���Q�%�"jF�����M"궨Vd�q�7h[�za�n7��C� @�!d�TI��B�c��YV4@@������ߗI�2%�� �o� ��G��T�b$�B�A�+s��ᰠI�9&��"E�)���f��Θ}\���z��,Ƙ�^�h� �l;`�0!ωa[��|O����G�&�޺�Ţˆ�ϯu]e-�3�"�*D��1H+��݈P�2�7$M� �\?ȸ�=":�s��_��\��zZW"K=)���}0���v���,S��7_�¸�ɩV^�8��}˘���Y��FJ�M�k���e@�{��!�	�rM�'�9�Îp���G#[/i7\�+
��Lۭ�u�;��/��޺��П֚��|*�uϔ-�<K%�m4���g
�Tn{�����+u;:q�/�Hr�Kg����6��\��`aj�Yx/_�C�����&�m@���߬i��$u�=Ͱ�y�����]T`���ڗ��s~�Ji��_ݵ�|�/^��-U��ž��͆\���2��-�4��:���?]]�j��⤷��Φ��;�>N<Y��$
T�(
9��Pg�9�r F���-bQ�c�;Boj�� M%�]K�O֞/��|���6Nm��s�}��.{G���'�J�
�S������FuO�x�(5�lgH�4>ڼ��|���S�f�N�lq+���'�G�Xi�L���������3 iaD�C�� �5-�X�(!5W�;����HP ��ջP�7�	����ߜ�����+43x��v�	(ņ�n�.B��"��@��;Q�c��?�<ĩ��#�@/��Y*�:�\�d��cj���U:�S��Vw�����R�*��3��^���v�>���Ǜb�R	ۂ��� ����R,�
�S��Vҹ�P������-.e��( <XMuj�a�7���I➵q߈�. ��Dl+@r5�K�Q���
1� e�+p4���J��Am�J�j�����t���+!����� ��K����A�E\��-�Ґ��l��'N%~FÆܓ7r��`��D�L��"-�C���b��FP��Ґ�`�Ќcl��z�q����<#+�:&�0�E	٫�{�����Ė��6Ĕ"'�VE/d���:7�B���!�"���_��ERU�/��
�GA�go��S��B�6q)�N!`��Zp���%�\C ������a6|K�M��D���(�X��~��ׂ-u�0+�zQ}O�n����PDo|X'e[Îד�n ?�A�l��������2eÊ�u��Fo4H��zW��GH��ptn��-z8�t��1��9���Y(I�<ӷog1��mRu;�fK8h��.I�Y3�ιHCr�q�H�p7E�2���|1�]39iCؔ2R﹙��ڎF�s�1�ps���p�d63�؇֩��X^}R��i��%��;�^�.H��?Y� +���χ����(jyc_��#�cO�3�v$3ξ�JlmQi��h��tD��mQ�/��ne�8���M��S�8��cM	�ރ��b!�P]��t�^`�r��'���l�>�(���	}0Î}�l3���:���!3i਑�xL���H��b��f�C	1�+X���y{�Q�Ǌ�/_��<r���I�k�R���������Plp���ȩ�"8���:(�פ���������E��3O�/��Zj˺�%u�o2E����桻	St�A�[I���i�t+4ȟ��դ�׊��w�R��Һ��Z��.:�*��l�j%�t]03�
��M&X���3��F��X}�z&��]Ǝ$I��C������iE�w>����CQk���r3�@�W��vx���$Y�4�3rd�l���P#(������b�齵��������?]	1� K�@��s�E�m���e�[�����o��^ϴ��e��z	/�ZD��x2 �&yq�A����Q=�,��u�d���7���ɲ4酭�@R���̵6���W�Ýk�o���T�7s�w4줂U��e��FLr��b͗�!����;6-����fG<'�S�}NF����Uzք�xm��� �J�e��T�i!9�t��g��rև���1W����q���?�'�	Y��Y�=���%�MG�FE���gt��>?��+��8;n�AI�W/V����nQet�s(}�~�Q�N�)��h���|�@�>�u���-i� \T�ƾ������wv���~	�X���9Ë�<l���
�+�J�~� ��P���,3�s�K\�`V,�s'x1��o�>�"Kf�
�Z��ldy�nH(�����,2�Ҵ��Ԁ�QB�
�<��� !��u��s{���¾
Sfā5���b�m"_����pM~�c�:K*���w�%7AS���Kd,B4�g�o2�k��U´�eCZ��Mo�q��RM~����c4UZ���V݃�>��[If8ɵ'9Ϧ��'��svm5�7��-��~İKͺPe{ fCcHX�s��N�F��1��e�6�Tݻ��Y��ʗ��Ew'?QP,�@čxW��[Kv�H�����C��<i��<��+j-d�)���a������\*@+�-�{T����7+4p<eYl���#�R9
Lk�G����j�Gk�z�1�Џ���;��oP�ڧbk�p�p��*$�įNS��DzOR`�$Y�>�5*""�ؿ+��p�Nm�MkX�F�9��H��,��Y9j�
(O��`u�	�c��. ��!��g	�u��}t�.zڂ�<sc$�`L�g?܅̯�%�5�~7#<B��So��,2�B�4z��Q��G��I����:�ql����6��r-������='�d$�hз�ͻ-nW����j�TyRH���i?_'}�J#������πh�b�4S��D���Մ�v*��Zm�I� ����LHZ��	�MƳ���I������Ήy���u�`"���/�V� ���`*O}���2	(��N���2��9�t���I6�u��|$����T������vJE��/bb1��ѧ��)�qv���]������o&��c>`VS�@G�6�������2}�(-'�Yf!�C�"2999=P3L�/��'=kB���[�=d�~�J`�b����Ԥo
���4*�P�dw5�dY���"|���Z����[��#*��m��p>n��	��I zx޴���5W��bְ�!�L�gbU��qW+@�ʖg��~x�^@�Ŗ�/�t�0{� 8�*Ŏ�>1��r�!Ȫ�;{s�Iď��9W�^ҬZ�@�O���_4�G�V�,�V��@�����	UFƤF�� =�]�Se�ғ�b��%��������W���LF�yH��5�,�S�gs~@8`�__2�����^�@�+�h�OU��U�_�^�@;H�Khi#��}S�{��啜��َ�Kn�7"�Ѐ��7 ��+e��
�b�%s�y�9����i[D�Kb���_�gxB�yi����(3m_1��c�ƅF��O>g�����Bv��ן;�f�6�;ad� T��s5^�ih��ҹ�Z r�����K��C,���-6`T��j������x��T��H
��D=�	#ns���� ����fIaH����~)����|�Gw��֑�G�@��<tY��ֺ�3�1sV��Z4n�
}N���m\�uU�� Z�蟳��b���?H�1{����6�0�	����UT~%:ΘF�g+R=��w��1TQ_7����� �8��LG�2�<��%�����W�|r�:�Isy��J+/Ig�j$R����l^:4�Ӷ+�ZfGdׄ���6H*̶���{}��v��z����H���A�L$��zs*�0�Wp9*n��k�Y<�:�ŀ��[8΢U%�ן��`�Ҕ:~tn�YU�$�i��.y�n{:�ۖ;bFu�����-o$z��AE(�Vx��!Q۸�0�\>)D�ˮ�T�ݦ�����w�&�3�֝�"��Z��N5k��Ҍ;�J�k�GwP�����}��	�U���8�_����g��aĴ��v��_r��&Cn��Ĺ!�P�6Se��'�[/ɣבHm_u�Tǀ�Z�Xte��Th�_�I���������;�&s4�.V]-�{�[��i��"x��h3AAܠy�J�߀������6
G.H�5���r��8X��m��͗cE��L�w�̱�Ĺ��U@�z��y���[�P=S�]R�j�K���@��m���f[�u� [����N:@ӎ��c*)��<L�i;&ׂ��C�E�ݮ�?�ӱ��A��7?@��J�1�sG�_8�����`@zs��U �r�X�����ɴ�w|�^�R�۪^��İ����n��Ӧ"��.чZ�Z(�`�~�no�Q��|�;�t~�ϹW�Q�Bګ���!�aƳ]K�YH�����s�X&�hq�0�[,Z��&K�8���+8��,�(Z��4�z��y�8�9_?���ˆ��0&Jd���Z~��#<ػ����9�#A&��X���x�W٬�s��W������'@������励�� <B��s�� �0����7�8f��l�R]J��;?� �aW�Y�r�_'FLseٯ	d�F��{R�J��'�LO�ּ�Z��8/���Wi�/{�-�5~���~}������a�Q^X��0�B�1�AI�i�/l�fSҗƟ$������L{���a���wN�<̴�����"Ĝ�<�CǱ���_��X����xzW��$w�tnd��c�xD�r�j~sD�i��f���S�*v��`�Z�y����ў[D����������a�2F��@�\�~"��A�7�P�T�I%J�5�Lʼy�OQ��S�����u	�/���ھT�'�ҹE�jAh�>�7�o~�%f^��ګ�b?5�P�)^����/��+�O��*�Y�)yj� j��HR�Uy�N]���]���tD�2���켳�<�켢�c6kU����j�����������3F~��_|I�NV��C�ጄ���Ϥ�2�ɖ����f�b�J?k���]��-XL
4W��6����_)+�k�G&Y!���z�B�1] �N����NEy=yN0��b_`�{!�n�Ĺ�$��2�A�����o�l�k���+x��ZE�F�٠��J���
1��D'5�����屫���Z�c]U��^�1��'��{<3�׳%���w0�x�X7ݥ�<PR�|���_��� (�{d�(f�a���r珀r���9y�(;��"�'��&�\��!���-v�1C�T������u�� ��P�5]�/��/7<�o�HY��bj|_���p�D	,?���,�BEI$@�J5)+Z�UgxG���:�;xYr�{ �3������Lz�O�rMH����wݒ��B�]��ɉ����:���n-��-� �!=��*ו��gw�Ѭ ����vt�}���iP��c#�Y%73�d/�  ��v%� g0$O��$��{��P��2{�����3\�*�Xr��/
������
?�xɺ��N��Cm�b��.�[L��w'����6�6�qաi~<^��<񉿞�8��\y�%/��T�Z�pk��W����=�`�����w�x���0(�,Cl>���Z'v���?B�P�G@���[c0�H�Č �5~��A!��t�b�3�8K��{�
��t7����5�}T�K�Av�i���@�D�� %�]&�@��
���}y̙K����}Fm���������x��Z���Z�v��ݦ=���� �m�sO*IEЋ�W%�`���f[Z[_�]/62�5�k�e��ۨ�Z��sU$�7I����k��!q�4�̷���J���mM��$�[�}��Ódêr���եB�����t������+��@�&iQ��ׇ���ҢP��S93*܁пb�`�J���	~2/է$,�Db�T&���J�S�}	ך��V|R�1L [{f^����_9�!���h�(P�Θ���6q�-��ia��\�'��gЀ�qR_���?��ZW�_��q��rp���������tE��Q���,P��=c6��\_$��b�����H�nGpM�=�������sQS���6x����f�a�����ç�'C����!\N���^����]H`Ɏ��݆+Y����E�����D��0EM!�O�?5^��dX�wn�&2�X��m��ڤ�9Wf�UW*9Wk�yW��+�O���2�?�a�#"�תe���X�?,e�fg�-y��I~'�b���&CgBj˷x�Nb��OΚj������ߥ�����7 �-���(���^ �^3��~A��� �-��(lc�P.�t�1tI��Ia�;�$gЅ�X�F*���t?ߦ\����D_����nE���z��%�N�K�3��A���n� �*�����gȍ��d��_�y��`�'�؁�a*�l�VR�T���O�=�S�ڀj���M�{��J�i��!8*.��ep��É��c�_��<���hghm尐^�G	A�%P�j׼O_GBۏ�������o|c��e���Y���2A9��!ǽ�h�C}u1ݹ������(����Xp���O�D�9�9+���Pϊ���r��,��"��B�۠?9�;1O��Y�����ݠ�b�5#D�5�C��ۣC�`4�a�����+?x!�J��pIW��1d���5�ψj>L����Q�����8;�z��j4�fz#��'�h@�{tQ����ῆpQ�>Q5��(#>	,������-#<˲�y��0ý�͞���Ck<����p�Fv����<�3a<�<+�9J�5�Q��`����ϙ���L�-���S1�7I����n4J�@�>���2�e��U��� ��!��1����_L��-�nIS�R�wÈ&xBB�۶��CB�$hE#mz;���#*I`g3Х�*�
��u���7v�(Vf^�?�g�N�u�$>��?����U����Y�*��Zў��>4�~��� �j:�@�9�2`�sA��%D�[F;JĤ����I�Tkq������?�9�1r5�.a
P��/�~H:�Q	Z}+������k#�ٔ�Җ#+&F�g�9�ycƜO�ީ3���:DF�86P�w�����4�'��ɬ	�~Np�G�%�x���'���y8�#���e���}eؽ�=lA �>��]�<r��z���by�Oc�i!?n��s%�W.!�;H 6z����F�d\i#7�4+ȥt-�t�|����*�aG?̰���K����7 +�0�^�Z�$'��p�}b��������)�����.K�U�w�<X��]F��|�
E����ά���t"��[��6��֬@�^�E�{q��2������3�{o�� D����BO,����h�k�6C[#�X�_!���g���:��F��䫈���"�Vm�-}-�KL.��V�ǽ8�Q�M
Q]������`E�BKLZK `�jp���a���~ˎ��b���R�i��u<�H�����WN�ޤ�O����RkN,�kۋ^!<��(�/�5׎�j*�����w ���������)�z��J{5n@C#x
y� �9��b|�8 vu�G��:�������O��ٞ��F����¯o�����zX���+�`���剔C�ֶd[Њ���b��LT��y��x�6���Uk��l���
�3Ŏ���WDd�#r&o��5�	��O��mW2��de+�U/W�#wIKR�L��=���RQSHH�U��;˧^�@��#��*YP�U��d(����J�J!n�?N�+_9�E� ���4����6�b��M�� �UR.~�բ��g�����z���aW��¤3S�?܃A���sM�;��IgeL��gܽ�����e�O;2L>��`7
��k I�On�#���ZR���)��ơ"=�c���Ru���B����:L�]1[�5�����<�r��T'9��GR��e��m��}�~e��J��G�K$?dN��[��GN'�-5�o�N��xQ~H��
L�$����u��L�cX���H���4g���a2V�T���q��t!��u��	>�?i�b��@Վ����(�]�,,I��кV8TC�$y�{�F�Le�\��.�Sr�%g4t� ښ��DUw�bt�GH�ZM�v̸D�sK�*1���I��5L�V��ؐ��b�b��ʪN�����S<���X
N��_wM�t��!�=�M�FR����d��4i���F�*C�O��!g�	�������}�+*��!)��jk��g
B���@:e���y3`����:��^9M��B��V%FD!1]ݣ���ݶP���óE��>���t�L�s�'���9��w#���*	5&�;�J�n��|4R�$zT�e���E{�h&TX�5y�Ûy������ΗȻ�8Ϟ��E.�܁���+�I����̟tb&�!��؇-6�z���9]���Lv!��"�0Z�r��qZ�-%�/v��Qz��aI��3������4F��f��|4��+$���*"��N�`��½��R���*��L��'�
�$·i<�#1V�� D���xB#C��lrh��}���Y���w��[f��1,��o��$����h� �p�n���*� Ay���v�(�����u�;��N��7��"T��j�{@�*;]v����N��5�^��~Y���uYc�(��V����*�:���i*��������
��D�w��$x���i�wc����2��_�\�R���P[&fξ�((�2m�P�s�3�L}.����~��!���i�'S�X!����H:��mHG�,�n��s�C �"n2�#2�5���p�e�]��x�b�����,[v�{��t��v38:�Y�F�@��Q�,����r���C33H�ǹn1�� �s�/�#�5u}'5A�v�3��%�L
�U"������D+�hn���;�Y'8L)T�?a-�y�]�X��n���?n�gw|�.D��|N9���Ƒ�9C�`5O�QFVf���kNUl�!s#A5�F]�����qY+����&͒���o�8�2��e�.���ʟy� oQcĢ��V:���2�jX�~Ή�W��]l�%Vɨ�nb�����GI�(ى��hZ�|?�byTM��qHN,�hy.RB\Y"���s�� o�P�ߦ�4 �o��	�mx��PR%qE7�K�غۅGN3���b`�WE�E�z�z�إ(��S���]9��#��Zm6���<��	��<}���+K 
�H=6�D_�� �b��=xl`s���k�G܍(��}O��dڐŃuE?�EԂ��9w{*{*\=C�֐��RQ>TNzu6�^���4 4#�;�W��ވM�ak�1��
�
�&~��ݞ1�:^h��Wf3�����������g�c�r,��+��]�J�.�䟐%�W$����֒�J��i�]��ҿ��ɚ�*6�����q� �s�X��BP��7'W)�^�ll�t�u��ng��^��2�����P1ѡ:^6�>m�B!Z-����[+$�j4���j����.mqWh7��uN�`b'���]D��g��TQ���33�Z. ���W�3�%�#A����oK�3�	h��y�:ٴ�[�.���ê�o���v����6�`F���mƽ�:R�����VK0ᜧ�v,�Ҁ��U�vr�?T"�f�� �e��q*�!�u��K(3�j}����
����9v���¼�����Î��b�[�V�T�
s͹�ӜS��b��L˭�p���w)ip��(���7i��`"���L�X��n��OL`/�M?x;���Y��3�0�f�H�����sM't6�jn�Q,��i?@�y���sB�cg�����p���bj�lSJ�X����)��}�M=7�Id��<��f�5��~S����[����c�̆"�̫U�`aI>�_��QL�Yu�:�F}fl�#��8���F�%T�����n��Bw����֞��7VCAUNs�"����~�]���dY!|�d�����5�=�:�����u��������Bb%><�^�����
0J�o<����mW�~��b��W����� x��M�z[ت�k�d�Ԇ��c[�}J0ͮ�
�t�%@K�ૹ3�j��V�.G�͖���Ƭ���o�D��-������O�IM)�d3xD���l�0p��}@p��5��Q`&6b<X@29a"��"xH�/�D�����5��ǟ<�����=�n�����8�X��hi�C`!+v:������~m�	U�I1H^7jd�?0����od�b\WH<">��7�F$�
�3�x���%�r�*�᭝�/bڲ��Z��W��M��������\�����[ow4��� /a�l��5�����5W�}':�%�8(>.A��'D�\Fs�޳<$X&����W�r�J����~��YI������D������eI�If�P޶� �x�E6��G���x)p��(�#����*�%���K�2�Jm�T:�F���*���+�=rD�$P�#�U�:�#��a��<D���=ˢ�,�(��+��go�w���?G2'�U���2��f6�J�|�m����G�!&3����D`h�N�0�O@�57�Ck]J�C}�}�~�t����CI�v��T� ���]?	��&�Ek�:���R�:2�-�qe�X���ڪ�Dq�wa5��6�M�c�