��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛC-�b�4�l�]u�Ih{L�a�u`dL��������]v5o�3�,-L� ~3�g10B� xW��Pnc)��US�W�6����0̎)ے����$�XŚ����PŎ���I������+آ.G籥i��Abz�D������h,ఉu;-{[��*u:�DV��i��X�?T�L�� Td������׳��k�1f/�C�Z��Dp��x��]�l�$���(�����9��{�]=���֦�֮*)N�np�g�9q󝼛�<8�0E@+���m	�]�RH��Ӗ!|�}?d�;~��hJ��$���d�)^V��@#��C�� z?�&��h<��?4��=E=}F�^+��b�_�h<�X�[�Z��n���9V����pN����q�7�����$��� �"917��q�B�7���W��I��5��c?���pF햓
ӕ�eV��Q��kD�:��,���׍���6ik-Ĝ���"��	Z�)�>q���7���Q�F,y�5����^7�aH��7��ʐ0�P�Pa�3/��\����YOߌ����V���cѢ�m��yS�N��#z�lW9aI�2�!�yq���͡ޞ�د�%GW[�t�ͺ,l�g6Hz�1��wx�D���!�u��f�ќ7����W�y6���H���a_5Y���h��P��.N��׎o![�B=��o8�5��7⣞�b�}��%D����J3�iUC������Z���ף��y(Y텽b풌��Z<F&=jRS*y
�4"���li��X*�  �%���?5���,M=Ӹ�0 �>5d[�H̍*�h��t��E���d��b�h�3�"e���π ��(B%����)��v�>;_(�(����<$�Es�g)�PQ��{�6U9��hn�A��B*�j��j��9��xF~�dD��o?oN��҇I�o�e.�m�l�~���x��C8˫cW�خ<�!�z��G2+�**R�%`��Rmњ~����l�qF��k���U�}�����6�M改;�(����+z�Χ��W<�pw�J�b�:�6��8e�-���3dܦ^On�3-+.�	��o&C�#nF�x��c:��,�߅M��i�@�>�A%R�%��k�i���@�v��B�}��J�h����6�=>��u0����([����&EۊƤP2Y���o���훻��*}F�\
���aK�{G��s�*.��`���T� `�m`��!�vE��{)�&9p�u��~�%�7lȣ�B!�����X�@b���ߺ|��V�`���_Q9	w�e�8����|��_>/K�\R}y��P<�{V��^tq������7EG9ɽ��r���ۘ�i�$�x#Rx��[+���V7�AEYpp�$�[�l#R|��C��-���%�L��G���u��}�w��+��&(�u�n��+1kvY����P���2O$~6���pw��c`���꛸�Ȟ�f��|����,7��8̃Sof�&��v̐�֓���3��ޝC+9h�#���\��D)���6خ��%!�U1�̏�K��o�<�0AKA?j(�X4�C��!�m�ώ�oC_DO=;�¯�|cԁ^��(V%��qM0|/��aCx�is�ĳ�hDK��(�/EF~�Y֕.�̈�b�7[��Gd^��'g�>�D��	>����rI��> 2�'�k<�s���>�g1��iLD3�P(�~����x� ͭ�G�|�����~�5�\����%^3s��;I
:����@H�HH��Y9*�� ����0~�m��"�BD�Tv���uG�b0;!;�-�e/�S�b�� Y�ߣ��{�� 9
�He3�4�W���U����au�XY�7�$%^�,�fewsGрl\���er��
���|AP�����'O�	�Ɂ���B&�H���NY�a�>�g��:��.+Xu��A��<i+1�G�.�j�A|��YKD�e��TAƋ��-�4j���|�[�� �ҕ��@zT/#�$ �,<%���v1���û^������VW���H�+M��u�A���#^�[���0m-\����?�_M�)
���3�d�_u-�PS]�]:��r����V�D-ٟ�(]9� ����@cϐ��R��`>-�p�����ND�A$�����KCr:��"����d��8���w_P�s�p��P�`��"��*i+�4ɪ���=evJ#�w�z�%"�f[^փ�-|�Vcӎ2��ؿ��(�����K�X�	�+ȑ�w��~�L:�h<6m�߸(4����D����Q}��(|*:�&�	H�w]�?�@1�5��%<)2���זm��~f:C�6���z�U�.f-�pxh�F��P�/[��e$���62Vq��)�Y�N�^�ߊ�Tt�k@6��UlU����R�����r(��Vf��{ q�#�HՄ��]P�~��d^\��{s�yᗶ&�]��>�n�˘s��m�H��P%�׭.g7�n %˘�o��jE��m�K�Y�y\p�Þ��S_5�xd���9�b�<��2�:+�m0s����q��H�$ ��?�?P�ֺ����%�m����5�hO�n�̃'U��:�v�[�|Gl>2�-M����؈W���d���mb���h�M��L��6(��P��~��V��4�1t[k�:�s��dy/�ofy3����
�-�n9��~_v��IP���G*�>�%��@1�>�)��9�Ʋё��S��$GP����^���'�z��_�X�v�S�젙Du�[���x����ҵ5�s9H#�6��E��9`qN⬴{�*I�ff�-[q�/�한�e�=�$��sj݌T(8��
�h��ň~�N���^>��D)�8m��*]��d">u?�4B��!g�W�%�6��r-|w��/�
L(+ʷ_&J�"q�s����_I6�y�]$l�'��'�E꿗�uy�b>����Z4���VryI�m�8������ʰ	� ��PF��ʪ������;� �w����_�0ʊ���L34�7��p�(��ܢ�\�m4�K��i�(�c�B�]z��F� ct��7d!���P���2��Fk�$`oa��Sj)��hyJXv�<�k�2*$
aUi޵1��G+�a\<[;�AP/j�$cHM� �otJ#��2V��T`�%�!��,�z�� s}7%�P�_͆�{Dn#R�D�̠�m9��Uݧ� �S�u�	"��1Iй���CΑth��`����
+q���d_����j��0���wZEU��	�`9x%^|Y����V��՗}�_��cj=f_֎1rj��=-/���p��9�G��8J_�7\`V���*��/�����q���vf�U#�/�+�ӆ�zp��F�$8d�� �݁~	w!,�$sl���Oa4���*��QcC���� �r@t���� ��ڛ���5+}�k��z*�2�	���������x2%���C0�� ��'c��~Etǥ���W�k܆bjf��x��� *=w:�-'�bhW0�#�X}z�D��!�l��>�k��u�R�	l���K�,��8�j���XTl��HY�^ �ҝ
I#VQ8�P�ՊÍԗ�B�0d,�~����4P6ٵ�ҹ|s�p ���ۗeF�F3�ݞe��@����p0Ӗ#�F+SC�Is?y���b����@��i�FOSr	*c�_���I��ʡj/�K/8����y�~n��L(D��s%�E��䠋�~*c�\��F�e����4{ ��(�g2��1��ܡ�o�:o�w$��	�D������h8s����f�#v�sx奪���M�ȏ�=F��8=D�o��!~��9q9���C��2� ��^��n���IQ ���� ��zv��.��Bu�.$���x�Zې�*y���G�;.�zn`s��2{1��T9��L3O��v�qڼ�\hqn}i�8g�q��2��<�>�
���׊G�C~{I��O���P�P�R�2�w����\mh��]��(�
D"�(��"5C	��J4ZKh�t\㫵l$��c������@�hı�\������k7�"H|H��.��P�#�@���J�Z�o&���[��4j<)>��ɬ��.��ՓN.��\�*�d}�(���i84�
��)e�B6^4b�eV=P������{~q>��N]K&�SP�]]:T�C����τ��#=�:�=�V����6�aob^FZ��y)��0ĕB�2gN�tSaH��~D�[��\�ڧ�]c�#c�?���6ws���`kW��v�|`uڅ8Q af&�2J���Y2�*����pv�YP��$WLt�)	���o�f	��>���v#E����b�Ô�Tp��$�b�~�����%6��A���^�3G%F���~�i��q�Qd��,X �hP�3�hy�X��z�d�yo��9�S
�H ��E���A���+��g\���Nּ�9f ��!aLTr猳�x��4l�b ����� ۨZ̊�M� B�H��/V �j��
:���`�(
��l6U��D;���XIx�I�y����+�{hs0����p�_�v��,�[�� �d^rP��n��v�w��"�����#܆�h��L�t����i�HK��~S�����V�IO�r��*��h�"^�8kK3]�|]�=�xhi��ÌF��p> qc��O@N���� u�f>j����b�NCC�����(
�ϊ�s7i�j�������Q}*0ƪyx-gR�V�%ʟ#ã�~�y��Ղ~��0.���ߒm�*L��㫁$*�pn���!��F�0���Ά��3�F�@Klz�1l�ȧ���Xv�uwD�z���H���]_Q����R\���\Pk�Zq���*)�:�3�*�8�~���
��/f��J/���go*��D%�U�����[��$r�r@MC!m�$�͜�4���M�q.傛_�~�'�P7~�G��M�o�F��v�烫�Ye��?��d �����������Z�z��n�8��%����-H	�r�1����"Q �b`G^@���x���C�P�%��;��w�L�f	���8ׯ����0BP�ʍZl�ſ��yp���|!VP5S�ӊJ�����I�'���\����ધ�FξkMz��+L��� ���1���1�ž1ADUx� �a��H��8rܜ�+u#�{\��TF."����=�x�|Mň<�"�w5��
n�|�Y�'��ȍ���������9.XM��KT��@�_%��ub�.\�(���`�n���U�I�Ҕ�R��`x���O/����P��s�E#� �r����[��!\S\�o؝�~����8s´���x��.kԃ�p�x��eG	$L�/�+u�*���0�ݱ�x)���!�����.b��~�	�O�!�3���x��ӛ�T�'�PԿ����_/�75K��fH��$���������8�4�'����9	��h\����E��E''�ۋq�$����IZ�J��4=m���o��HN����Yh�i�a�	�~�a�!2�����6��u�,��lg�z)elnj�l����[A���a��-,?�C���b��'�7`�?�U��4MkX�
v-�~�q�N���#���TB�aˎ�Z���+��Zkv7�ʶ�	Nn;�(�.��yi>%�I��#�QS�\���v�k.�"gIt���8g{k��"�Z�˲�Q�k4���~U�[��e�_Ұ��}/k��2��#��erl^��Y*�Y��n4�*��U���������r�ӕk��M"�4p����M��&G�6�,V���?�I�A��[����?�S\W�y�l���)	F�b��b`�z��)}���c}������E�<�0������N�H��{h�v��L�}pl�]_G1�s�]z����\2G��g��'�[P�K����И�	.I|�ۇ�|����`�4�JV6����Ts�>X�EE^Yn7cF��M��r/a���j���A�ꕂ�</�^�G)��{�cq��^�p����Y~�"��Wi"�b�CS�d�4e�a���33bP�@�b��m�zW��ma���oy��w|�2��u^ƶ�g�b+�ե�uN�U�{�)�G�2�+�/�M�����ĳZB4.�_�������ю�t����B�
�0(�3Q\�[/=1g��"E-Itݸ-.��`���)�-h.���p���/P�m ~�#��
�<�u`Q�*�O>�!�h��`���>H&�5��$��E>�7��/H:���U�9� �&�K"����4���ʅ��;
�Ա�0��D�9�jGvx|�G5j�:l�LO9��lsD��	���A�	ÿ��
�]�ra�<i��~SYr�d��*i|Ņ�"��JƵˈ�?(����E,_�;GM�(u��8� f���m�TtD���AR ����9�Fɗ��[+�#����G�� i X��+�$i���dv��z����x�pU�r�.z��nh=�
�&t��5������D{Ļn+��I��$�᷼%v۪�A
z���f�1��)����-
k�?4N��Ds�߂����{&\e1�͆�5˖&��x�O���^���x$55��e�+g�y�_��!���?��̨\Z��DX���U#�U��f�<PsW��h�٧G�q�*[�d�Z�/O����8laY΋��>^��y�0nʔx�^�N��1NРur�T�������~�$��s{���G�e;�]bd�J�kP�`�T�qc��ά��yk�3��c�����آ�r�����n��������I�lQD�h� #i�����K�bDro �b��8y���zR[[����5�U{܂C�K>
Yb����ܮ�-1e_.�����F�B��!7&�����)m��V��4Y��A�@7������������ai��.ӗs������b/Y�L
��"�V���;8hPS��KW�2
Τ�$E	�E��e���N�f��㗩�F��hz�Iֽo�R������HQ��tl� ���SY,�&��z:3Q��O�3;Bx� ��Ǳ�m�8'ɾJ�I�B����~/]��|rv<8��y�����T��1ZF�	��1��=dc_[�5��-��n)�4G�oQ���y:A�'jj��g+h�dGC_'K
d0)���_��N(��;Z��@B~ʘb�k��R��Y2��
c����@�^��jF�w�
�*��M$�2QT��R5�<4w��4O��I>W�&�MK���]��eRx/P\�������%n�Zj�\Y?d&��؈Y3,$�<
>�s��X�V�d�I鱢v�cZ������>~�1����;�4[��(ާw\�a�4SC�ӏ�Y��!����@\ ���gg}�q�c���Ѓw�n?:F�q��F\o�ɠ�<7�PN�%>��)a@M��i�P�S�Y�T#���>R\��?}uF�M)&f�#��&�����+ܞB���z���i�Wn3�a�Iش��vѹ[�(�˔�ܿ@|R�A�w'�lV��wI�s�WO���Fn�/o��J�l-�z�������Q��g>^:x[L)�PqU�W�ד	f�5��?�R�F�X����b��'ײ�o�ƣ��Dxi'5����;�i�w�s����7�D���/!�"o�A�9��,x:=S�.팞ȭt���NV<�� ~.r/�\��?�,KX���:�P!�P��Ep��eu��o�V��ٟ��-�%�@�IS�3��n} Anv���FأG-���{���3�ws��N���ǃkɓ��"��5� \��.bM�wK�.,<�/LM��EY�H���ӈ1z#'żue�N�h�N�w^���:o��3�.��=7��vЯ��	v�]^�5S���^o�K��G@�X��N��V�����)T]]�W3��k��3ٔTAM��av��{:���2��p��������Cu齩3���]����]A����W��k�6(Ki�v�J�L�C��0�gu��UZ��S"|�~��'[o�<�6�%�E����w <��ek-�Az���o5;��A��F��|���{H���8��	�eQ���=!d'��R�	�Oa�����	��h���U���&ּn4#js;~�]_�(��<_��[_ú�A�1�ƟX�r�]yȘˉ���($,�W����u�V��d���Q��(�3�	���q<g�y��3/A���2Yd}�ju�i.Յ�n���5n>��گv{u����M�x�'&�S�r?�/���d��h���;�nho�I��o�#A�V���~�c4������t��:�M��e���8�!-^�xܣ�Ҷ�q�t?y^�5�!����w��ooQ�G�\N&�����%LL4��Г�L%8����#��&۾�Ԕ%5��٥��!�&nP[�՘(�4�=��vy��J��K#�)�1�%�8��X>�	J(��gQL�v`�1�m�$fH{���;�_�*N:fƅ�0g1����.I�-�t�zg�v�Y��l�@�}���(ӛ�u�$L
 ~���-@��Mn���O�E��r*8����F����T���BHEd-7d����I[�d)9k�a�/S����m-[-��4�8��?�q��5�He�!�Ȳ�/��j�0Cniy��p���IW�P�%+����D=�T���	L9���Es˿'�jQk��/.d�G�{�������
�����?�A)�XD��έ��ԭ�0��,����?P{E&�C�վQ�#�c5Z���"oYA�
s����G#q�rּE�A��3J��#z(���2��st9j�p���)��("&X/�aD�nJ֛Ѻ��+s�y��v�[�0n�M�fw �M�*��������k�ӽ��"�D
OX��'΀B ��e_���+N���4�^�
�(5]��a���ρ�Eh������*?Ϲu�?�l�'��z;� ��F�1�s0�Z'�Xp<����,�����og���S9�'�Vv:�Q)0�ɐjp�n��J�Uɶ0~I�EE!ěC��2�R�x�rU�d���])IM/��@�=��m�S�j��R<�0ND�k�	N���4�4��N��&e�_�&է�#�9w��)`ZX�2y��ΙE�g�e �߀��&��� ���.�M�� �3�����1�C5A}�aU\���$���S�����6I���,�XoN� c���jh�i��J�M�f��������2�C�}�Jʳ|�R���<0����_�~5���֞j��/#��ׂ�y
	l�j�CWMtSGE��(����׶��!t-��絛a�������T(��>7��X��c2E��>e-�7�j�׹M��9D՟:qC}+��f�p}��g�0+���8�֙�'M^�	b��>
�8�4�4�Ńz�lU�\�)��:��I3>�2(��2ɹ촳ʹ��>��o=�ւ�<�Tu�'e˰�Z����v�y���.T����m�N��t6��Oc
���T��3{+u�I*��|�P1K���s��1�Vȏ�W ʹ�����i�@��r�}J����c������%`�[�Heҝ(�CϺTj�����C�hT:���|�}��Hz��<���j�\����g}O�� OP���������PIwWTP�\�^4@�}��O�P�c� �Jn���Ķ��"���eǎ��־�$Oq=OL2�����S/������(�'A���:gnnYP^��&�yo��;$?*gڊ>C`��Җ��X^�vIF���>�"�=2���7��h t$��� �ԥ�.�W��s�RX����
]"e�Sn(��v*���IJ��6����Ji�����yU�yVRG��p��\y+?{�*���4eS�7���[�	�E*i��� �C��a�W��|�Ց$��"@����>-=���}�>_���Jg�J��F'ݣ��9ĭ��I�~h�f�����l��ۭ���B�x�@�F*~0r���N���HŁcs[ȼ�s���,�����C�f�v�ǫ����W.���.�R�j��z���0�������N����~�i(�V+�~4V'��Ok�#&``�W��a^���8j˹����C����U
�^pa���{��:�X�X��9sR(���� �K��'2���Z�F�^¹�����z.��YY���B���	[=���T@���V�\pg�F7'����y���0��O�B�ʂ	�%u�qV?Gk�R\�JCVj�+
�����xq���XRO�!�3�'ѹV�p��+� ���[���]�9B�G8=�2؏��Ӕߍ_йl��]�v��Ư��z����i.��u�ɠH��+8�� �����1�b���ܷ����&�O[ӎ��4@���w���)�)��G�	)�BZ
8X�Y�o�0��p�y�Ov��KH!�ʄZ	�h8�.W�?J�����p�_%����Q�TM�W��;u�}�w�å�6�o�%�1��ƒ������_3�{>;��C�I\�$��Ҙ0}�˸�q��h۱$��u���߽�N�UWރH"j�_�-��ח�C���L��n-�
z�9 =�$<g��*�ڴ�(��AeJ]�tR�:2CU���N���k0@5�`�)��]�K�s� �������SJ�Ϳ��8v���ƅ����R���'C�	�`����؍w�\2�������g3�*r�19,��5\D?Iw.� ci��QƻؕCu4Sf_:ud�#K<	D�S�N�
1��&wQܲY����=%Eal�$M~FdT�s�O|��	7z���?���F�e�xWW f\l(aA�<ş��7�"R�S�C3��6ԃ��t�4�͘e����Z�c��>���"E�}�����ԧ��K�Es9L�Gг��:<��K*����v�qb�f��;dU���"����ڇ��1߀ J qg�7b^{�I�%&,v���FQe�z���6�����S��,&&��H�{ϓz܇}t�f�[���bg�3è��m+,
]�N"�-����is�)t �%x����
�h)��%Q~���<����/ŗ�w�2��,����;�2De.󛕦}f�^\6�)-�قO1j	��Ka�w**y�%�xr��3R�|țL#��(\x��q E{tfE*�ܕܜ|�Y�H��_%	Al�NG�h%���B��x��+��iV��G���
?��_=��"�<6��a�!ή,��)��@�S j=Ւ�<XP���؞�B�wL~_�7Ͱ'Q���">~1B�l� �n�S�AAW�f�?�X�t�/���&ŷ�7����6q��ӚHjB1-eP�e�0���hi�*'��.��3� �BI����͐r5���76ٶ�<v�C��r�d��GS����t!���x���{^M�\�K�%UA�7}6��s�tV�.4���u�ϴ�# ��-32ѕ���i��|�Rz@�Hӿ/��Q�֫����O#rҰ�*ʛ�ʲ�}��L��o��s���2��e+aΊޢ���Yd�2qN�s?�����(��$�yC�)�l̀��#��/����O���H-,���n�P�3�f��:��rY�g���յ��{@)�"+41M�1e��j�V��� vp8�9,�%_��~��PƙR�q߶N��}�&һ4��4m�[.��y >�.�IO��Lvۀ�Od�Qד�9��,FNc�	b�Cl�~ Tx0Mҋ�>� ) ��Ԏl�"���/�J{�:��K��X��:L$9T�S��;;O@Y�����*���Z@��"��Qw�оNA�~,ߑ޼H�����C[N3)U�A���A>Q4��'PY��(
N�b�ez��H8z�A�r/ɝ�V�%�/+n�v��� 9��Ru��,�0 b0��'^q[a9��  w�ٺ,�_pB`� �~�(���zŝGE�f����Ǜ��_����av���
e,�ڞ�Vx��[�BL'lڲ/���������J>|��8~aچw9ެ@g���]���>�r沟�.	���D����ɀ��4�J{��tK.�����1&Tꉎf�M�8�_ Nx�=�C�$���q� ��e6�y�_��}�E���p� �R�����MSf�E�-S���d_�;H���c�Z��B��[��0�݄�O�(��w�Z �ti{�ЯI�m>�M�u�Ats`a|)15��_����y��x�hm�D��:���H����p��� �A�@k� ���Y�'��_�FQ�8�`.�������}8��闝`DԊXk4p�9��,�]�=��t�(��7:$��neӝ9�k�뙭rdp���# +�m���H�P�Prmf3�C$6�� ֧-��xR�؄�9Fz�T�h��~3�}��w������F��N�C�5��wT��4qB�28�/rU�<�Z�!�ɛ}q܏Tvɓ�����e˙���(��5#joj@�r�y�Q���/�-����K�-\`���G���_Ү�1[�O���Z���f�*�!��p�T�U^�;�"w˯^Zm;�kg�K�ʤ����w/b���h@��iڕS�Z�S\�D�6��OXg}��ؗ�cנGn4b�3ҕ���#����\��[�H��8�"�|�s���_ۇT�l��_�S62�	�Ǉ�xJ�Ѿ�|[S��_,�.W���A����6]0��S�-]n���H �}Zu�.P�k2$8�q�����.eS�(���+D�Ғd��/r?���#�����fG$�24�?"�eA�J)���Gs��y�?�m�dgo��	5"OQ�i472�!��Y���Dyf�C�j5����'� ���-K�P�\c)�<E�̙��x����GF�'�Ҳ!{�]�2�G(ɓ�)f6������z�U,'�/�(qa�W�N�ux|a�|;ţ7C@��(�3U��u?AkƱ�V�"$㕖�$s��$������;-<C�F�B��]]�d�w�q�V1��MW��I}&N�ӂ�65yc�O͟�At�.�G�M���Gm
�F��<q�F��i�v�e;��6[��?�%��I E4a���L��G�w��G;BX�O���^�v(XtK�7��j�q0�QA؉Zؿ��Պ-ԾZ0��ޤƪ��aT���S�m�Fj]V:l��&��m��
b�1�B���/C^��� �;��6�
*�����o�B�w+��U��-���b�mX�p���.���N�=���3���fւX�]�B�x[+A�h�25��o�8�j���ϳyK�w�AF�WV���L�+�E��pU��آQ��]}
uU������l��E��0�lP+��C��6S����W�����%�l/� ����B��o�O}��.�W��踂1&�>jk�4}��6W�y��V�)�{�H�3CD��f���! 2�*���a�������g(�-Ia3���A?l*���n@�E�l�����I����e���#_�&L�&C�R	��LD7�3�QͶ ��^}2,j� '}Nm%a\���D�҉ J�K&�DK]�W�`�a�//����sa��D����h��;��q�0�����Q[�E��S��}N�/�������Y9q<��0V��K=6%.�\��N{RPn1ڧ߂�T��͐i��
 �YϷ��,�p��� ����\>y�TD��%&"Z6�<]r\6�0v��_#�T��'��MB!��Z�}|F��ݑ�p�7c��ӱ&S�+C\4�FQ�|!�v�C��̹o�nT�5��B$���=SlF4�GC9'&�}��z��ChHX���K���>��S����/p+�8S�� hBQ5y�k��k�̌��n-`-:E���	����ö�i��<3?ǅa�xp���s'rs��X��Y�<,3;�)��k\����Ri,�%I9��L�3f��ueGE��0N4��v��lz�=���c�Āf�E?�d�gX�W���\֍��ڕu㳿��n��*E�ư��{���q�s��kJ��;����|Qn�ӧ�(#������v�4�Q�H�PP4y�08���v^P�k&"P�jB�e��N`zj3v̵�c�}I��|�].3���K��
N�4f$+e�F�"-�J2�Sh#��{��[n-[(��B#���7tp�c���D��E��Կ� ��J�3?%(s M�m,Ki]�Cܱ��&��ʅ�z��_!T�*zH�*К�LpV�͘\�u�AM�e�{�t�	]��GG�A�c��g �ě���4���?�O�ׁh|�17+Zڛ�W8��dڐ,P1�����H��F�^��!ӥ����{�U2Yd��v�>��,H�w��Io��:��+��!^Q��}.
H޶,��~YX5h<�#;����>Ϳ�g�X!W+�9�i��aXq�F���k��тObD��D�ފ�N����FCBv�{̪� �M��y�՞�f�J�t�d���=�(D�����}���5��N��x]�~��.�U˴��`h��*�G��?3���WЙ�ad�!A� w戓)��a=j��"2N�L�[��]^�9�M�;�k6�u�ff�ڕ�(�;ID#��:�a�\EiO�67qW?K9��9���$OVݴ������ ߤO��1*t@ko3�~��k�~��(��]��nt�_���3"�T��E�j�d�qx/$�EW|β}5N:R��"�2��R%���q|q�(��~����Pi� ��&���ϫ�M��@^}/�:�A��n���Dߣp�$�'�Z�^c������vȠ��F�{�ZCB	�z�D�:��K�OY�L
�i����i4�%��O��4�~�쬭�Z�<6<@J!�.,6��{!X�˚;��AK֫�چ�|\�� ��$>��GL�Z�~��Cv$�r[�q����6�� ��9�u�pJGD���������q�`|2t�"� �h��f�����#�e�?������H���p��4-+}���
����l:�N2�j��'��n95���8���	ڧ�@Q4э��.G'��rk^%��P�I2�XL&�cz��R���)N�A��0����R���b�����J��BAdX�O�OȖ�F(�Y�
\(��e���Y`�bAϸ�T����������U�y˥с���޳�}ZF�/ B�p�4x��͏���56L���~�ٟ��X�YX�b+� {����8�`�� զ�  �,�0e�������l2"aFy�?������>�gi�K�w�;�D����]>��f��Id�R��h_]��[}jF�b+�X�?1F�ݦ��T���=�\�M���*��!	���&���'h���?L�ض7Ʋጹ&�Yo�����\.FB*!��Y��6��C@�F1hx~≶-o,��|%�ZM�duH_��i{��#�"o� ��ڋ>����8:	<$�k�R�h��J�5���$iI�ԋ�B���.͞��gff� g#��
%KC�0"v �4�2N�*�x3�V�~��X�g�WF��d��;�p��Ay��O��R�jqE0)K��]�/��qH�o�c���l�p�����v���=�B��u�ݛk�I͏r��]�:�p�m� M乶QCp��r���-�������3�X�kD��0_	;���o��ƺ/` \`a_��n�1ջB%�u����XA�xNJ�Bx@�(�F$�b< 
S�g1��|�{e��e>�j�:�}[���Ρ���:� @���A�X�:LC ��ή�-0\��k{�¡�8�M�	�{NQ�68`}~&�頀
��
uO5�y���i�C����/�Ö� h���f"���IwԬ���#�Ǜ�s)����J�
9�a�:1#xSU�����'�я$r��'�$����⸁x�޴Z�/�IK�k���#��d3�A��`MCN"^W�e�2�w �)��^��J�^��|��¶G��?�%��k�������h��uօ,�|kw��-�����"�/�=U�O�����ΗVT܎1~�3�����v����b�to����MF��Fo}zvY�i׫j�L)=���Ad��3�@�`S}@?
3�9��u(6������2�z�Jn4j1��bO����>"i��-'�xxr)����.�l�����F����w�w�Uxb�4RP�)Ja��L�!vN��=���-�B��H��o*�?�ɩʌ��~e��f�"N���$�TĂ�A�º�Hܲ��\w�W�����w۹�}=%f������c�c4��av���φk�i�F�G�AL�+�8���r�F���4 ��\B���gj��C��?87X.ӓ3pTs �W�G��z*��m�:�M��'������pi!�^2O���X�Hn�%j��$�Joؒ�J3bbg?*���o������2� v|����.3���V,���nU(c���2����?e�,��e��ܩ}�k-nfV핰�qD�Ϟ��4�Yle��%8��Q
Y�o����֚��d92]Gg�jA
��⹤L�@�e��~�������H2U.�z�/U^����Za���A��*��O
���i��^�*�ӹ�ں-{��n�!�|�@t큀A��"܉���z{YT����C�.-�W�͆�����jf%�Kx��%������_�!��ZwZ� e�} 0�&�n֘a^��]�����oe�[	��$k~ ����:���j�d\��{���S�ߥ�X�Ĕ4�Lh~�L=R(_2Q���,����䍬)&i�5���*�;�Q�|<���ejm��Ŝɻ^��n�+8�.l�"#�� �.�'
��+��|Oޑ%��Z�𣶍Z��^V��kkF�G�Z���^g2��:�qqF8$aaOU7��>u�!�	�D����%{*~?^u���Ҽ��h7���;-�fje�N��c�����%Qt@PXu$6��HAی��,���}�}�[d�Y%�<�� �<��Z��j�^��r�ip�_��4��|"<Y2�g� ����Zx����?�k��pk�W��P�Z�����h���ЂcM�ƚNR�� 0�dR� J�S�$���(��k���H��pt��ɧ��:j�7����j�~�8����'����C�9Uh)89�[���׃4�}�p�2�û�TApD ��߀�,�*OϹ,Y�q�V�.���#w��g��I}��&��l�%���6��C:�Q#p��J[h�Ȇ j�f�t�������Uxc�J?,��	��_�pO�c)�T԰�r�V��p!��ғ����V�G�Ũ߮��`��[����N�(�ba�	�c���u�9P�C�11a)�t�a�۰��� �� ׷���4hMA��}j�� �k�H����!�_[����ŋf`�=(u��m�����2�Q�QhHϠ������Cĳ'��-�j@fDMt�|�X���k2�,�gH "̌9�U�چ�AsDc��HҞ�d���]��Ѓ
=`�6�ޗ�c��L�����D��b�����BTp���x�]g+�鲞V�<�3�m�*��9��S�����|�;B�"�x��ZV�bS��{dCɫc��+�vvd1��&��y�;�?�}�|�oS�b�����6��9V�Sx	��y⩜+�/,��=�z��(�����6$�d��$Y]oZ�Y?J��C-<3��"���X��Zf�~�j<�T�3��R��B�=��joT��?w�?�y��^+�m�t���#�Ɉ�e�ȭSQ��ў�z�<'N��O�A��N�?R�p9~��I��ϰ=��%B����X�О�����)�I������ŉ/&�i�XQFInQ�4f	飪��A����̐��Yr����M[d*���tӢ�P����zw��&<�t���Cyq����vz$2/��5\���	�MK8�����F���?���N��!�C�0x��B��\���A�R �s����g�P��@{��6���i-s�\�BT��L����N�H��_�5�\�1�VAH5�)3�z�;۔�9Y%�H���c�	]�(I�x(�j���ZA3�<<�F�	ѹ���H�Ú'5�1�	X"P���w�ea/UzGx�P?SE�>(?�a��a�|*����
|�4�) @�^�y��c���0���=�C�����.�wW���M���]�Mg�Pb�Lt����	�%:��c��8��k)}?���g�"��Rx�X�)�"		����Ø�L�U�Z ��-���`!�t�/���>�2�&�d��rz�a���P_�#�%��cCA�	�������`�v/4�i�M���)f������Ac6�h�^	���m�Ҿ�|w���ka�� ;�놵¢������ H%y��<d�	��������x�G�a򘪮�% k� � �X�j,��?Ebǚ�9�p�{���]�ȮO�+ �E�5x����9��$p�������um9��"|�P(��7P��C���LEB�6~Z/�ᇰY�F�'��V
 v�z3�͑2����;��U��I�YY=���8(6!����.��~`�������+��YҦ��>�GBF��.���떨:�M��Ҡ���*jQ]屁j+�^�5����>�0�"�����u[?��(:���%��p�o��L~s������S��˲Uu'i~>Do��Ô�
4�;�H�K�\1������ro?뛏^}�����y�����2n����{6=�Ӯ��Cf��ը��h�;����@�*OR��|A�]�Z�i&$6�\KA��B�M+_-������̜~*<�ʜ���jy��o����d�t�)(u�� \�G��4i@�)o蝥/�H�ɞXVtiw����V�b����5�N��l��E��6@a=`�q�Gb��|��t�!qL��|�4^;��N�t���Q���|,W9���8�8�{}_,�bӿ�2��x|�.!���t�OU����@��\��a����zb6l��O�a�x�3`�YJIWſ&�vR�� Sj�6&Ù<��[�_��Uh3�iS/14�\�[;�W�����-�J�����VҀ�Y���3x]�k��C����Iad�;ƋjĨ��KFq�}9���/���؝b�i��+����P	�l�e��Th��o���b;y]�n�WG�p�Y%��e��3��Ŋ�bs*�8o�T-�ͯk�Qa�Q��?�O��?�>�_��dw1��?��N���� Ѐ�<5`�~SO���4�R�D�����(��m�蒡T��Y2t�� 5D!J�6�W%�U�X	��O�<��g���sb'8��)�����Yl@�T�fYT�S�Q�6X
y8P6���ɿk|ŇJ�[ �� J[%�u��Z����#��RS�QE܉��fC�G٨�r2�{�'4�'��������x�K'�Z̂9@|�r�_���.���˃�ל9E<��?�s�z���:�qSP��B�įB�M�x�w�R����m�4���B���_�6���)c4"�7;'�f�◤�דt��	���+���y{�����2�t�
b5S��HK�ajz8U�Ya�DA;ޣ�Ho���[�;����(����� �#�w I������!Y�D=����I�J��!O���͕�b�Z��>��V�H������u�I���v����|!A��o�ˎ`���/eV�[��S�A*S5�6�[
�Z�e�:/�5��]N��^Gd,^�[�ݴJ)ܖb2�gà5y�nB���6	0
0m��仐G��2ՌgC�h�9l,S���A�F��g݁{�HϼG��S.џEl۬Xؗ����/p'0GϿ����ԕگgm�Zh1U|�I���Z}�Ϡ�������E���J���6ؒCn�M,�-n���7����_��j��
��1���,w�0@���d �/42M����	]�ޟdB��);�C�Is���䝉�d9���'���~�aN񔞿��hG�gW�������ו>S׼@�1��Z|�Y(^��-8-z�AEˌ�^*��,����Pⓩ�/ ���a�����;=�xB�������J3�X���Y�~�7�ae!1���m��<�RNK��:J��?������w�Ң�L���#�Mw��+Y�!�B7������И��Fȧ/�O�a<���+��2Visߥh�!"QB6�_J�]���g�C�:���3���&��{��M�u|�Y'������{���s�Rk���r���5�h�������v��v�v~�����2	�R�&\�^�E�Ǿ��$��D���"1W�q�q��+ e&���-Q��p%�	b;��[�Oio�&��ÿ���Oj�X�@<d�P����G��K�F���I�����ܲ��&T��.��[�Z�e�h�DOO6l({��u.�m�K\=��~
����;+�swqRE�ϵ�)f��d��yq��7�U	8|��U�"dR���lgP�7(�e�~��?��[��ܗ��]�}ݭ�-�8s��
ƃq{��ˮ�I
�It_[%���6�coW٨�R���PS5�x@�^Տ���d�JVY����i��y�TO:s����%�)MG�ƙc<��vH��e�dPXP�k�?�&	����!8��6��۱Q6�O8@ˍ{�Ū��N�|êݝ@X�����!>�l[���7�04�O�����.�
xk��ѝ����H$#V!�A�T�Ӵ��TW���E24�b�P�yHb�o�4j���o�4{ۺ���,�UG��8�rS従4��\C��E�u��/��4x�)��7�(P�۵Ha�}.�b��dNv{V�Hu�DW���t�S\)8vF�`���(�R@q\�� �|A	ȩZG.��`�&J?II�@A(&:2!�M%�آ�}��:���=U�( :��� �1��m\�'�?:��� �&�a!62��'����Z���:L�Oȥ%ﮣ��Ԝg�_PGnȁ��`}\�켴��+<� ��HˑIt�n�Y���h�u�Ĥ��'�c' `�i��s�ݿG�؊�m�V������<��u���#�KxIq?ځ�oR~^F�b���/��7�����4���r��Ey6��xHP�M��5�����[��i1j[`i�ߓ�!���?*���,�a1��}��g���Z���֔�b��uJ-t�4�9����jk�����N��,�h�t&���ՠ��9�m�/"�����	�������{��/���z@l�����(��gm&?ፒr��6�����&I���'��k�^+�*�=��h���~����]�(�v�*�@�f�\5�����`F<��$4b�T��l�&ci�/�&t;P$��(WdH�InW�7�p�DDיɫ�.���Z&�f�>FլxO�}�԰�t�g(������]����
�O3�9�N�B���.>�}?�16(i���I���Zv���B��h��\��'�q��7|OM�k��с���K6��@C���l�~��.G����;I�躌lW�R'xG���+`�1軃܇�D�<���d�9#��O:��A�ElQ�N`c2	{��-�\a{�L4��S�n��ʧ&��[�/�=]'8S�.1�AM�N�Ad6�\���sԖ�z�I�z.qrc�yy�Q�a��j��r������Pt�:.���\��xl�3��P���0F�GF���o�w\!+���0.�4b�A�^�@��:����Ǣ�# ,�a�;�yr�!԰;Ð���#�V~S'�J�&Ur�c��{���sBp�^��@�L*g7���Bq���6=��g��J��'g�`/�����A2�H�1��\S�G�g����D�(��EC��5du$ ����g
m�5-�
"^���	�K������Ds�����&9{n�/d�H+�%�~آ����~���l���D/a��G���P|��_�>h�����q��Ojj�5�w���u�6?��%Z��<X1OLj~}���7�~�h���:a+��,�&a��N!��62�u� E���UU��J�jQ�NT�T�
s�E;�d�o30Up��(�l���.V��2k�Yj?C^oT�G5@̃��40B��C�� ������L�" -Y�ƹ5�yV������t>���ϥ��������=N��!����*>U���y2��.�� K}��j��1E���I��|����i��_zH,G��jd��ݑq���>f���9�Ys؆����8N&������F	�z���LAE��0����	�S�߰��,`��=/?y�t�N�p���"����q�;{ʁ=5�:C���P텎:��-DI��-� ���W�y'��#�h�� �9Q��mU�Ze�A�%�#�������x�]W�K��)4.���g�y6�^��g�򬚟�� 2k���;'��_���ߟ�4���U!�:P:7��ڀ�����n������X�9���%�5v�]�DN��;�
�JB���*'L��S�&O��պ�J��A��h�]�I�)��5/i��r���P�5��A�7w���/l�x��K����؅��+�d��Y�^(��A�d#�w��m?/P�o�E�g��.ե> �������ۥ r�B��(/��h̇�#f�ˀ�J�TW7?$����u��u=.W�B�&��&�Cd����H���4h�z$Fdm�Z�p��W�w�&��W��3t͡pR�n��(�	:_���MŬ���h��~4���2�*���)b>(YR�|��������#���:�5f�mO���i6��Uۜ$NC�{1���(�7/�y�(L��!�\G����{��A�m����D�%�R�.�r���?F�QS_�Q�l�ޑ|�D�EDdq3�\�؞9�g�_y\�ۼpp�*� y�gb^��_R����\���M���Yq/zhލa��;�'�f�gXe6O�I�x7�<x'h�H��I��g*�p6�o53��	Z	�;=�单~˃��,*�\j�� �\��� %���_ي~�~�4�ގ����H�AE�J>8Yq�l����,4Tp2\F/5�(6" �E1�`,���ò5�;���a�kQ� /�U5^Hw槜(S�sy>�V<c�N�yN8ƾ�f��3Y#
�sc<>(���h�o��X!�܀$������jB	�.u�@f�5my#t�͋�gW�����1%	K3�=��%��`n��H�M'�R���dݶ2��~�Q����Jߐ��|<�UK`ș��Xmh���^�C�o�9�q.�	��mI|y|�d �k�<��8`<ކ���vU�x~�0�I�.W�����R`+V2�K�E?�a	�S��t*�@gN��\9LO�hF�h�b�����'7�^�B�n�M�.0��tH� �۪��?5މ&�p�����=�B^���o��B�z�?K<��~5߂�(����$vr�BFQ�Y�0\�IoGu(��,��+JA'C��[ݷFw�|Lzg˗�eX�y����BK't1��K�ښE/E[�S�3�\���S���]rnvµ|9�.�w��ܩ]Z��U���ͣ?�u\��z5UY��XЕ�:�l�v�$�"$�����TX���h,$3;2(����e �z�`��F�S~�-
$*�<0���^]�u@|�4����H���d��'����w���G�KB)��D˱H�J���ܨ�BȔ�Ԙ�z��l3ݱ��&��a*`r�#�^y�%�S��b�ѯ��p�j�.�� �d"�:--�	�l��>ܿ��#|5[��jS�#�[���Cۘ�@��@�p����6���('�xbH؟�0��t؏��{.��Hͺ/������S{�Ö8�HNl:����#s9�^a���b0p"V���q����xN2e�\��z� Ҩ�Oڳ��Q��S5������E>��O��j'��c( s��|s�Oӓ(�p�rIjx3'�(:�e)DǤR�o"8�L���L���k2�:��k���
�܉C��\}1V��u.�j#-��BWh�G�)d�p|:��޷�s-�Q��D�R�G�fG&����b�e�g����\��R�� ��5���7(����������z�����;�O^� ڀ�υ��qE/?�sr�'�^?�u��Y�\��q�|�٪����"�V�����DT+�57��J��/����sq�)7)�Z:1b����Ւ�A�٦��(��<Wղ$b:�����a>	�_ƃ�+u9�UY����|��k>_����,�z2� ��-?�-ӡ>%Ɓr�	��d�4�ŗr\�c��ME��/ʶ7h�2N`���RdV�́������C��R'3zW����E����o?��j�儦K���t�x��a^��q�h�����qՈk��;��Zh��`��{>����h� �����`Uٹ�R�R�秎E2.b�Vb�$z/I�m�:��>�N S�6"S��U�6рr��aʯ-��
O��AUc�� ��Q!��m�qi��}����i����.$ml ��s�����Ta���o����~U�X|p��