��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�����'<��;��A�%�Eo�e�pggᡍ"U-������'o����4�1�$A���ǭǖn�q5�.�Z��e7+X7��u��]��1lN^4�w�Bɿ��{˳�YY�Qz��E�D�����(������'�e����QX*���dȐ���G�ݐ����ϗ.�-����U����Y������.d1]�t��?1�YH��wҖ0w�t�Ǻ���_V��>�!�؈�����hC�w�K�H.�q�Z�i��lQgJ�U����������l��`?�R�����tے�7pj�oPp�K��J!�3���"
�iT�[WQ&����ΐo�S{Q�/{�y_6�wJ��;����3�xO�W;�J)�%�>w	��X�b��%J)~���g�%E���"�KA��P�8�we�m�:@�e;�����	��J����)�7�@�-�#rٽ�[.{�??0,����m������Zϙ�Ԇ�;#�5���6lf�����Ӄ�~�_w�&+#0rS�RSё��~O���O�����k��C�{/��u1���4w=
��4y-�3��{)�k����rm@+�ڬޛQKUa{�&��:�ʦ^�DA�t�Z�14t�|�Whh��36���~NS0(K�`�o�k?u33H����ܤɱ�� �K�ce88�5��~G����V�������~ޗ��Y�Խ��I0k��3��Y���ߧj��Ͳ�My(5T��l�a8|��:.!5��q���m�ɤ�n8U�.Pf]�v���U|9�(���"�O,v�R(����L�w忁�^*�������bg�A�V��H_�^KS��~�����"��&F�e��T���H�'�3�B_�a!��N�*%�^�=Yvtf�?�ϰ�_9խ֥d�S/PIp��6���K=s�g��݃:CGhRP�Ji�]�mF2{q~�'"��U�$����}�s��F��zap�+ '�틷���5xB�0��;Qz����#r3QC���6�"F��d؋�V�\<HW��F�-���������yL3��8�����;֣[���F���kU�F����Y௙h5Kps-��vð�����093�G�¹7�o|QA).�TϚ��ʮU����.�4)}������%,��{�y
�s�Cr��Y�aQ(d�X��o�����3�@�>`
I+1�4MR�]0( vS���q�T
:� ��M������o��uOM�j1��e�N��;����P�pgeoS��I�	MrkI����Y��^���E(��:K�5��%�}/:K�s�ѿ�;���X�r���9{��?׆\ϙ�&�ӈ��%�Y� 0�pȼH'Q)��>K�
ֳX*�~��(9�g�,C�HA�ƅ^O�+�h=`n�X���pU�b��|��Bv�/DhN���'��ׂ��V@e���*`�8VJ���f��+�*ѕ�6�T��'�@ic��G�H�<�A^����D�e������n�����6�l5Ӭ�Z�����e������A���G�,*J��`��m&��zoSW��^�^�6G��͢�L����WLg��fd��u���<��C����?bTS�ó@������1ES��P{�2�X+)[ 8������x�&@��$7�DL*|���tb�+T"co��d�@*���/w}D��cŜI�^ٗ���*'!>��u�Xm@V�����1%8<�*W�T�M�O�ת@R�ǏG��T�2CqX�t�Q�^8,d8�z��p��ݭh'򯨖,qtqf}��k)q���'�!Mw��_]>8u�RПÙ�"�X��@��V��=u������9�MB��lc��T����aC����M��y��&Q�BLn��k�?o��3��G� {��޼z+IT����̦j@i�&,TKPUoFj����5�_����Vm'9N���OK�l<��w�3�~+�lL�`���
��W9hu�r�����S�*5I�4��i+��<��V�$��TU���Ǉ>�����L+�c���{[�1���%��!G��V�#`�&���#O�u���HN����b6(L^��a���������T��N�0���)���~�̚1)IV�[�hy�_$u5D�'����+��(�?�\6����>�82f���ng;K�'���P ��yπ�vn�or�R���]>����zeH��TZ�I����-�	�?�Ț��}��XX��CK�*K:��|���I�z�s"�TVxM�;-{�߰���s���&՟��XD7�8�Ȳ�w!!B�Yl 8��穼������j�k��kHɀ�����fC�.�^j���n-brݨ��Su{�B������q��8��.�%���y�t�a�*��a�ۚ�"H��uO߁/G#'=q���������DaY��]�9�1e*3z�:Y z�C�����>���q{�;�~��m�Sg��W�G��rz��^��*,+q�%w���]�4��͗����<�f]��0��#�q$h�׊���
�M�Q�b���g� Bk�dm�,��~�?�Ɗ� n�*Y�4Q�iq?�8 M���:�fWܺF/=�э�(�e�ZayYٜ���!�I���rd\а��m�6��p�1=�����­0���C?�����FY�����7Y".�!�C{�{��d��� ���.p1TƄ� �ڼ�z�M66�2e���.s �'��^큫5)�9�XA�BXC+��K
�Y]������E�ٛ��:\;I�{dQG
>�8YiO�&�"Y�GU�	��p��8W�UHq�E� �s�E/@d�N�bO�M���њϘ�B+9e����)�{,B��?�֗�d����Ɖ=��TIi"�T�����n/`�x�)�!����Ȝ����6�j�%������������_�8QM��%���� �!;�e�}c�8�C�1~��Ϙٮ���%��*o���:c��P�\��^��uBK,�����l����t4�&�?z�h�C�a`�܅1�o�#fdk��pe��v��IG< z���S��:S�P�;"S#B�,[�NK8>��9ȹ[���Cv�e'��f���*D"�
17�Ѩ4�-i(���N�a4������ȉ!��FkW��L�� _7�474]\6"�R���/y�z���,���kZ��+%cK2肫b*�D��X��k[���0��p�:�}>!���EN���]r*����͢/b���,ne-䵺�vH����ܼ�<��^h�g��:�������	��_�Y�Z��� ��Y(��̤�yzc�^o�nt��_�R���~X��of�E������釀�����o�BA��;���0�Jњ��E��)��r3�к���-<��Y P�,���$K���Ys�X��i�{k9��t���gc-5�B�m�)BC��C�tg&4�m޺����!�6���
�p�	������8��9�w뗬bf�D����`��=n�BI��xaɿҽ�����&@G��HV����X��e��:`��J�N\���V@������>5�X����/���mL������񍠼9IZ�5��d��V�=�}�J�,a_��Q����,o���|��*4وz�y6 �۴��)EeL���œ����� �`>Q؝��S��P���E	���a�
��.�B/G�
#Kc��m���J)�8� �NPճ�%���*[�/A�������
,�T���H'z�W������x�6�L$*fkG���X,�pi���v�]wxf���7b�>��SZk���h�ce{D��'�fݗ�M�W�5I7��9�J�繿s�	���߭�z�+u�OJ)�
s��
�����)�f�k=H/Y�2�������+��O=�+'���d&%��G͇����/��.�]{!����.[��s�^V,� ɫ��f
�VRn_}��/Q)���zj��cY����k���ܾ]b)��/��Lr.�A������ԫ*�z�j;n�_er�L�d�����H?V����e�f�(�
y��0�����)nŗ)��}��h�wK<�G����zQ{���+���$ZAXĒ�2йoI�cv'ֵdy�=�!o�!����(zP���V
��1���x�yw�f�]o�9T����D)D��S��>�e�W[�`��y/�p>4�^��r4��s�������*}�	0��I����/j���2O�Χ��OT����g+�K�Q�̇��P1�&�v�R4��Xٿ4�f~���*�6����M�G���P����q��q�k/u�C#Ћ��ZP�j�ѝ�c�ŕ�;��X���+��S�3�86��+U��S�:`�料ߌ������)O�(�:E�Uei9�1��==�e�%�������e0U_ڒ��g�1F��<�u���f����!�k���r��:��� ��X��>T@��c�������
��y�"!�3l�`{���믵1�AE�[
�H���2� 7�.j��N�[�Z"t"�-�U�[>��$��H\{+��Lؗ�`�?�hk����N$\���%�H�:�,���ѹ�3���*�t�Xe`��xFU��I���8�@c��u\{�������2hN�v`��IF�3If%gQ�}h̉�W.2���H���s2���}���J��Ʋ/�4g���6Z�5p ��[�7s�sR��}�0���m�>iUz���+:I�4e�Q��A�H����99�Mr�f�F-��,]P���oP�h��p��=>��8	��S�K\�{�x_WG�H� b���e۳�^�p�%����ѭ�|��ѕ���5u	��F���bF���O�䰊����m!�a����{��ڂ���:����SƟ�w�<puiז���>:���\�z�%���O2��5MT�2
V�/��<s6r�p�<�g�Nۧ&�9��\��ʿ�>�un�:K��&�� �߼��~��0��}k5�k�� ����B`%HM�I�$��{��x�3ˏ�5�G�7]���`B�� ��/ ��JN�8��\&���ˠ9������HvL�`�n�_+�ʟ{�#��Z����S�s|���^�+���o�������%�k��Ђ�]��_������&�pX���/�_Ͻ!��8���q��~n�Bx�J��~&C���� �O'N�L������C��5��,y�-��!�E�"��n�ˌSQr��b�P �P��˕� LĥuP>@���'eı�"J?�<�����8?�?EM[8#GRM�`&�s,K�mV��.m�zJ�y1��{�����3R���'k�A=�$�h��]�D6�P��h��!o�y���E}��������N��k
���
�r>qc���2Ӽ�!�'F��F����m�7�_��uY��Gp\�49E�Rf�g�v�b�+����a� ����Ό	˃UY<˷L6�-�]��=G��z��j꧆l����	`��hg#���s�f�Κ��ߋ�0=��6�+
���¸d�S�������k�S����������;a��w2��EW�:x)d�Y��L��zh~��z5������?����Ns�=X�<�vz%�!-��������q���!>{��h�0�v��+9jE�%���>g�N�M�Af��;턻 �=�Z��)\�����iV:ŸI���,om���A�
���\�>����h���=B�S�z���a� < �}�I	�!�f�i��5<���W�7��R6Q@6�����Q��yg)b��Q���I�RE��VD�Y�j��$$��y*��Y�����}D܃V��xIC�q�vgG�5�@�H�����Q�sȣz�[�U.N�a>nȼHgr�W��p�Cq����]h�@$��1�s��l�ݱ��/�����+��,��aH~",����T7V��<��~8G���W����7:Q�[�m@>�L m��o�|큑4g�L}7:
�=��hؐV��k
;�ȭ�?wp�tbvԜ+�a�a<��R#�Rʆ��������V���?���)��21Ъٻ�}��� ��uI�c�y�+�O� �V2--%�B�e|�����TVRi��� �_u��@�*�Wc�"o����Q���|�i���-��6A�d�T�/���%$�����+�/L_M�f3�՜5^�fe��ʸ�i�}�]+��jt��p��bD�%�d��#���Onn�m~�궩��7�a��p�(���
5π��=	2�*��{��uSZG(��ο����,e4����A�[Ӈ�u ����z�,���n�铞�θ�Y������ͷ�O��B�^v9����@��c��	R���(��-�j����l>�?���L�T��(��B�yo����l]WZp:5���>#A�N(م�O��D0��b��\�#���\|,Z�^W1�Pkꁷ�|�u��gc�/������!���(��g��4��#�9փ��;��l��Aݨ��_ ܑ���Q 2��Ϗ���q76$/0����G"f0hպx9��T�^ڰ�-7��l�91d�۹V������U�ڎ�,"ڳ_Q���:K�a�d�{`�p6��צ�$��e���e�75hZ�ٙU$�;&�On-�m����;�O}o7���C$w�Eq!�e�4a	��v�_D6�V��+��*���Y9��gR	7��S���J\7r ��6�
�`|O"{��8����U���WC���.�GZ>F1����p�R����[���?�����/�1�����@G�C�s�Ϝ���3��n�Zօ�������{��d����~��u1� ���hB2��N��5�L-��)����)q|C���	�Qٯ@,$6�JC8+]�<�^/���a�9�)�r�M�x���*�mX�a�9������rӢ�a�&%�>z3.��]�cN/s_�Б��7ea�%A�� �� ��bysԹW�^����Y�lXx�S�����V���c3�&"�.����AR';UM���ˌ�-��+e�jt��\���t�i(z�E�]U0�֔}�q2�PTKU9�Pjl�u,JD�2�c�b��3���_+��E���y�8�T1�����q�A����޳��
�מZ�xhKF
���p���Q��E�>�Pȴ0_�N���Z����q	Y�?(�$!]�4a�0B\%� �p6��x��Z���c���g^�ۯ4�.-"
���t�Nb.
ש4,��?�a>'�[�;�� �N�����NcOq�z����୲DM�6�|9�*�Yx{��fL���� f�"#�^ʏ�Q��ۦY
d��Y>LT��b����N���H����k����ue�Sr>M�\왂�8�/]�ƞ�YX7q�Gp�	���c]���f��K�Э��L�D��c�u|��յ��ǞDB�o�=�PVU���R6���L������D��hƪa包1�y�,���`�����,����
Ѓo��̷�m3��xE���_���UVՐ�����N['��]@�1��5�|�Fxt�[}Mu��`p�"�QI�FJ'U�R�ˈ������|�tA���:�}QtǾ���F�Gf�A�jpP��*�"/�x^/3�m[��!���
;��Ȑ��l��$Ni���H�_��柺h���!U^�p�[���r��?�.ϰ(�َ�kZ��}�<�;k�Z�$ԎQ���~+�c����Z����q .+CD2�mCQ��v���^�I� �R�L�^�E����߇��#!��Kml��戝g��$��r!',h�RD��ˢ������_�}�.��6J�]/Èp��K����r�[TJ��\��K�٩��'`b�uKi�IVk�y���9g��5*��T�q��B��)��vQ� !�|�O����Dڳ�B�z�Fץ����(��=�7;Z���4O�@��&�W�w�$R��.����H-��<4�V�8��v����+2�4��>5���/ ��~`ETdٔ$ua��s�ڡ�D���x{4�9��h�"@$p����n�-�u�+��mB�Qr2u4K��2��}Q�LOsh걩�@[����9�
�����"��7 �����V���|K�v`�Yw�Q�r�2|����:���{���ކ�\!�Z��>�gsP���o- @��h#^N�g�@K4f�w�gJ�nѱM��x�!�!�8������������>K���D���_d����	��u6�Fߤ��ZV_�1�Ix�Nu��6ix� ����n�W\�?;�z�N!��b ����t��<��a'<�<_�ݶ� �q-"[�F��������oSd8uҸ?�*F�oEC�3GЮ �n�r����
Y��|�V�{��Qvo��~�yq�z ��8�����.���n���Fm��H��s����%�s���$ �����{��a �s�7�n;Si�hzHjS��"�Μ��:����*�~�S#��;P1SU�X��r������%M)X�����0|4m�MO-yDM���y-`6-�u�Zcy'�5�F~���n���,iK��>H�P5#�J����*\��:{L�Q��?qZ�X��%H	��%?Ȩ`|Oʦ���:mFy[Q�5X2�Za��w�@g�+�U\��]3$r̒K|�D���^��N%ԥ���4�%��~�p(>ͳi�
�Q(�=�u� �E*hϹ����nK%��0k�Vj��$D��I-n�@�0��[�����= s"R�4�hٷ�*�4t��/ǻ�[>�Pk/}�_v��"D�N����)��U�w��;���$()d�:��7bd�cӾn�s��4����z��z�7QD%��c"�ĲDr+�'$!�tR'Ê��������`��;b�ܗ��G�R��	���{w�mI�/d�(�@��1�wT�)4�4�?��]����b�)(dH�2��\���"�g[���BH\���#��L��D��y#��Xr��m��(�@h8y?w����_��@��>��ˤ�]�.M{��a?[���ҕFxk�����i� ���v�l8����3K'��&b7����=�I�Z"<��z��2�kؑ�4�&ŀyEQIU ��i<O!�������D,a�����p~Wo�i������8�(֕%�W�YhN%����܇�cĜS�����ő�oH�d�΢g���;`��6� �TjH��Ԏ�62/<g�L��7����RK�t�"�\x��5G�cb#�2O�B����x��0�\R��f<�(`�^�&�[2�n��~���� �lX���&
�04��=o4�.��^9�=����s�qi�l��@%ѹ	��)���u(�MʫޥT[=,{�D�@߆���Yc��W����@��Vj)I�
�/?
����T(rVȱ��'�.��&�0����րF��}*�a�1"�ػxi���������V�[G�LHpt�,�Dp�qq[AT9�_ȚRԸo�s���$e�B�.e�΢��T���o��G}o���x�����[dA�j_�\L�^=���M�X2�%׿��w֪,9-8��c䯫?�����lr���:� �C�S�&��"�C@���aYS�0�A�f�!u��rj�G��Qm�ʓ@��I�� �j�~���`�T�N�_�����d>�=�\_�oy�k���C�����T$�"��Ӿ�0���4��N�١q��r�"��R��k1�{e�ޭ2s?����g(�����`��V��T{Tɏ}�;�\�^��
���O���B�d���ol�=��;��*�����!�8&'��8��͍��`[�l#�	�&�0�{=5R�Dz$�N�-�y�)+�8���G]L��$�1�D���0_������i611mQ�0K��9JZrUО�)��d$+�0��X�[���}Ժun!��}]kf{�~�-8M
�Lr����J��L���Ӳ���Lf�<�%��o���w˙d�A��Y.W�)e>�&Υ�^0
��>gX{�-'�%ߤ�i�n+v��(�e��{�'��ߓ�}ls�6��!����UߙW��� ��A#�(��1�"��v���&����P�C���v٥��9���5^\�+X�Υ�D��\�v���%����@hw�K��Mz�ޢr�8�`&�p[2+H�뿋�G�`��*�����"�B�c2<	���I���V|�_2@4�Hצ��Ea�)�i[yv�i#G㏯�Ob��4j��:����`ˬ�IH��D%Kjg���M�H7FzG?X�a�3Zs3k�����O�4@Ue�R%��O�Α ����R�=���6���̰�{B������c�(1��nlB�Α��`�UM�!�&��;{�M�du��f�75����ti��9�2�PH�J|�@y�g�pX#��A&tZ�9�l(���X"�m�D��!�,��I��2I�~���0��Wg�����x��п���7˦��-�>,�LP�CG��T��������K)��_���N�ݫ�~}O\�?��Ņs�T�jz�ݾ���{�u>�k"�VwN���^!��~U\Y�[?Vu�����θ�
�u�C��O���I!�2H��?G�͘�6q����e��_�H�1ԓ`��Q����Si��O�p˟UW��Fdz�Ӻ��euO�L�_>v ��{!�m�mz�Y������p8h~~f< m�r�G�A" �#耑�n�_�����̖!�2@ǿ>i����Wl���rOa㡸��)/�1���R`R��t�U���h�Ҳ�:��i�u��j1�Z��Dȷ.1Ħ�����&��%U�w��\�������v�{��STP�z�˕m%tc`'��
�, G�H��6���`���Zy���1%�k �F-�x�6�T��ۉ��7;�mLG]�t�U�B`��Uc�����j���b}�p�FX�u�����E�[��7FA���)�����QD�3~�SI�l͓�D�΍.���F���#�㇑�F�/��I+ɌXt�bN���8ހ���4'�5@�L\�yMw6��m4nT;ۀe�����M��kp��A����F�-4�}9��T��D�!�]k?����z�O�V�o�z�������B5�VJ���&J{� �B�ee��3��]НǊ�}����9+[#4�2�Ѵኦ\7(�b1�ȹ���`��7����
Pԥ��hc; ���h�]o\b��y�7��N��aTx�F1�w�K�6�~E�y��^+б1�3^���� Ƚ��8�ޜ�@�ʵN֯§�;��`�IDP����t�o��8�[�:A1����۽��2�
���p���
�@�f�"fg�8	����Y��M,�r������	B�T�c��(�&?7��*���� ���\�07�Р���C���`o*����uMM��k?;:?��ŧR�e��Y��!��(J���IgdԒLFmcL�?L�N���P��1�V��E��#�/������%8�����h����� rOs9�����.��I��d"M��n��Ä��P7��jw�`(xP�*7B�/8�1auS�Ŏ��	%�|H�q�հ|^� �S.8A���Ԏ�U}���.�00�YJ?=|*�D��PH����*��|��U�`y� �6#�R�,� ]��S��� ��-��N���*���ɞ9�Ve��Q4W��S�b��;Q�=�,�աz�֕��=�� #v�7�	���*�'(�@�˔�5Իj��(��x���%L�Z���(����¿=��ctO�P?!���=����o!�8�hVm���҈L�I���	�E.�y���ؐ2�}���B&A��8(�e�9;u
n�4 خJaeV��T� s�2��ρ�^΢�QIN�����a��_�8��,qg��-|���ew*C� �_/s�xrS1�j����M�'��	l��R$N��i��Q�N��K�_/����G>�Gh%��ETK�Σ	�+_�͵h|b�J#_����}�A���8��7��&!�]�����0-� k�¨S��]Mb@�~�&���l$��3��m|�	�/n!͢�Q� ��;)_N�u��D��R���q�eL X�5��%�WE� =���V��0���r��T�/7��[�* P��SZ_������ou�{h���H�!�ac�i����И����Y?��/w��q���I���i�2��.p.���ӥ��ݹ$��ճ��*�HPA��<�s�4ԓ��a*'Py������|�uj<)ީL}o�� B��a`/��,)��$dw -��Ƭ�o	��G�\�7%��q��ӎ��p��8v�H7��:��% d�V�ͷ)�2	n�M+-瑲I�/��imJ��rl�9>���Wp*nz ��i�N�Q%O�f+u�H�I�z�����} �eO��9�J-���2��-l���W��{� �Lw-o�w�o,1�r��)M|�
N�_6���)Is�|I#��{EU�
,b�z/���8W���n�Ҙ�):��}�6Vr��٦����i�Su]���US:e���֯+��銏b
���~9?�,.�G7�x�̱r�C���n����M��/?��2~�&�^������
��_/�}Z��ָ۫��H\��	��{�N�����&O�$���%"��˫Vû�:�C��@�p����Rf�&��{P�8�v��kT��ց��e��b��[�D������x�f�vo��Nm$�$(`c���~>�pF)űwTs5y#F'8�t�[]{�Y�T�O��Y��/t5���߮�q�5.�
�
����tl�7�;t<6�}?íM�j:|0Ŧ_�+��E DæF䵺8��z�r�`�*VN1$�>=*LF(ȥ$pa&}�=� �� �����4ʚč+�
WB����8������2\
�]<qi�7��>�sY�D�_"}Pc,M���e_�ON�	F`S���?���?���y�����oыZ�4�@�Kr�A�����Ն�lmj�¬)�����UI嚽0��(U�o-р$�X����~`�7Ü.X�w��a����L?�
#J*#�^x^"��f�<8��
e��j����z])9A#K��My��ح7S\L��P��c��f��#I]fS�'���eW�,����i*j>�jG���Ik��A��[V7�n#6����9��nA�?�zF��D�Uc=�֔�%=�>'$�gA;S��`(v�
Dy���!t��G,�j#{y(��@��W���b��DL�r��՝ehL�+��^��#N%�[��}R�Z�F�7�<]�����ԄOi�����o}���}Ȳ��/!�Ћ�[l��6q��#8��W�yA:.Arϲ	B`ߟE���`���T��E���P�h3�hܠ@ ũ&sF2�_Q�tu*���Sa�� �Sr,�~�iX%���m�*Z��t�jg^���O�(�\,����!\�{���P�Y5�$�/F�7��_�G�>�j{i�_�^���>�Y�DX��<�y{ܩ����)��p���w4�vC��v�\��^��S�./���/Me���s��Sʸ����X����L�X����� �bS��Y~)#?�>#b���WX��W��0�.�N��=��q!�R�	�_8HZ�%�Y����*#\g�^��R[�L��i�'8�Ѵ-��* �/���Y3"^W��g���ɛQ��Hz��F]�dB��f�Omnm#4��U�{́��콩0C�29	�pk�]k�&����oFN�^j����i�.�F�͹R�����	���mz:��[}X@��!_�uÑ�6$��m�)�lJ�n�k��L�p��w�,[����Y_6��"���K��~d��~G`����l3�j��+���M���q
V;��/0��"��'C8~�o�k}u_XA,�AO�yRW����e� ��jF�G��˵[�� o�e�A��n�q&���D6y[�m�άC�G��}'�?�b��z@�.�t>��9&�@����4ņ���&��+�5	��J��!����>�r�i��x$L��-i�t�I��KZc�^;q�F3i��U5�����h� ;V5�w�8�A��R�h�!"P�^�TO0�3�����i1v���j`��/���Y�Η��.�`�"�/d��>\%������Ti���	�,f-Ϥ���-f�As��4�ElVf��'Pu�^,u&N3;���yq��~����Imv\�^�:B_��RJ��%��;�\�UF����R�G��
��~��[V�%W}�@�v�R$r�r���OgN���惴4 s�� �p/JgZ�0�V��B::�v���(�h�R#/�;�ج�PX�r5��W������t��!$?�I.;1E��*�hݤ������&mn�q����J�r<@Ͱ���bj�Mp�4�����YU
���>�]3���ER����í6 �jW#?��Sw��T#Z��_�{؈�����R��E@يl(s=�J�vsM���@��}�sOm5���U���츶a�w���ӂ�0�l�	k����Un]!~���ΐ�ps��U��LH������?]D�pr�ա�2��m��=�Z��ɽs'E��(}T�d�U��osݞ+�ve�����c�v�����a�������Q��7��w�@�����H�֘���G��x/�n%�fC��2a�� E�(Ϊ�+��8%7Iɛ0!v�.�N�R.��>�ϼ��������<e���0��U���_���Y�R%l�R���������9&� �j�p�t�E�$O��Ak��̦ӎ�a2m�7d֨�%Z+4��i��hw��٧&JLk��ˣ�(W���5�I0T|ױ����j��^w�l!�ZP�H͉Ȃ���g��� ����Pm�:��x��Y�㢩��˯��7Ǟ��9e�lM�
xi��a�8^⒚tU�Q�S�D~��[�朌�y�9�kB贴J>�bG�@.�U�j�hj.��פtZGPW���}O���UbY����v*�a-����$"/�ʸ��e����
��уRr拰��ebdn���j���;_4H�S���"�0���a�����Zx�~dG�R�JbrB&��Z
	��5�xe��N��#{n�=� ;ce��?/�����yDT}��ERln]��j��"w>pe�ޖp�z�;��p�:�R� ��s�ʃ3>�������V|�#��b����?;eX���르6�s:-�T�
�oH�3A�L5Z�s	��p"�q���_^A+hwצ�Br!>��|��l�-�?��0�3�}%�4p�ů�����M����*���L��/Q�ʖ�G��X?=�:E@\��@�Ի�	���@�'���ҡ�v�I���+�q��w���2M�	��ѣ$Ɔܹ��J�9�,������r���f��W���$���?�C[�0��i��Ar�o���r�$h2�#��'\,B�?�+��=�w �Rj����@�_q95gkR�����Z��l�d��������po+�Í8��&�,t�|�pk���n��r`��x�ҙu�J�����;_����������>��jᥱk��I��mm��l�?��k��be?��0�ђ\��ۤ��kJ�i�P4�_�Y�><H���)��vv��C�׋0�E�Y ��@;5��UE��'X�
αN/)�X�>�0�K��|tg��V�����[��T&	y�7d���/��3�ɽPt��m�R�$CP�my�0#��i��S���c��R��qh��n7�]�Jd�.c����:υMu��1�\�u�