��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛD�))`�!�����h�7L���Xyu�& �`�ա���+�X��i��o��+�|� �CwZ�bot`0���;��3"f]J�,_�D�(/l怾"[-F|�t"�êZ+�P�� 3�ט�4�yx�u����4IA�&����v���b��a�J�uWmٛ�ސ��	���<ڶHX||��,�D�#�%��f�C��/ڐ?�{̔�%��Q��vP�D�
s�חdK�Z�d����bĘ�/~Q�]�o�����ki�+����κ�A�MZF?�Ye�ŁU
�F��ecg�|.4��\�~C�.�َ�~/�$�����1�g,�T�����c�͏�~���p���^�+UR�?$�9%x)�ќ\� �þ躇���N�f����y�h1���w0�N	��O�aŽl[%���}��ܹ}�l�t��	r�~��y���a.b�۹I,�����ޯ���.k�^%��r�,=��lZz�~]�����#C�:�
��_K-��ِ�e�c�f���py�T���*�5�Ï�G�
ւ~��<�7}�<#O}ڡ��N [4����Ѫ��x�x6��H:�P�o� �]���r,��z1	�ǜ��^���K��~Z��f������ ��h47��M;y�=jͥxب��N����[r����2���L$M��z�@.���8�Ws�T����M�X���R�Di
·3zɀ�F�j� 7HI���j\�t�G��U�l
�2OB-\*Ty��L�ǈN׹kh5*�r�J��B��U~h�����|��$0Jg̢[�K.K�#�*���
hT|�}�B�
s6��5^�0����	d�H4n��t���9�+.�t﷤UF�`G�͌��۱���he�����vFf��&'�(�yV�v8�O�-hD*���ܨ��;�9}�G��Ux� ��L�v��瀹�Bʕ3��"X���tjX�2�#"�Ž/0��i��D���>��2\��ހk����/��^����{3�1�P�L��Kc�-)����R���~5��`��(���n<Ma�����-E���:W��E'd�p��z��7�2=n�|����L�i�I-U�T�,ԟ>�Õ,'�x��WyC/ZR�M;�ۓ6ﮝ�I�~��P��>���Hz��Qt�F�؊ǵ��@8��d��y�Z┒!M�UB�����j��<o�-��qX/�{��US��y��eOO����4#�I���g�'��%8~g$ⷲ���ܗ,}˽�?���v(�/��R�Pz��r�d�l2QI��i��s�.g�oH͖h	��*�ބ��~�Y������(7��ق�~�(8&���w<y#��W�؆�����q�F�Y�)��2��O+a!)rZ.e��L[���4%e$�_�7�����D��ޡ0�|�L*��_�2%��iL������>�~��l4�M0�� M�͕���0�̛�RDa@�k�kAN��.��	=�"ʎɡ���P#����V���E��0`ԚPT��C0�PE�L���1�WCm�cJI�B6�DA#��;��u�#���N]�a�z����awwT�Rz ��Z����,�$����������ܕ��NmM��Lm[�L �9�P1vp��ee�q[����Y���@�C	��Q���n�.6��J�JEHg��.W�����:���G�������;��苁'g�F{����|�!�ȡ�@s��F���8c j�*��(��x�m��2?���E���!S���R�*�J��xC�bb|%���E��h+�%p�l�B�A� ���	e[p��qg]�"��8$Q�)����D��V������c%�	)��D��{���kSpQ��dX}��"(�㋩�E��}�'K3�x�!K�XT� ��.#��8���C|4$#U���km=����tx���!�ˍc��I��|��`���_d�aI��2��n-k�w�]�Xz�h�����P��Lj(q���bv�{*�{kl�d�=�m,���98g+���D{4�TE�4f�e_�1�q9'�T��d1�L1^�j���F�ׁ�x����Ը�l���q�w�.*d�bH� �t�sem�'Έq��>���yJ�R2�@QF~h��n�¶��4�+n	k��]tM?5�Av�}��g��q=ºf?0b�^[��'���4Y)�d�%��������ș2�2W�LД��aF����'��f�F�yHRI��x	�,�W�qj1u%:b(�د����ګ����Gm�U�~ڜ�Y ��]�����k�ə�EU�ן!,�b�1[be����}�V�]1pC���R
��][���,��C���-1a1�f��:�D�w�Q��������!�Kx.g���l�T���:R�$ �덚�0��PΖ��`�eW��I� ������<������Q�^�O:دz��kr�K=�5�!�����Ab��o�-�j�TS�s�I}3XU�,kI���B(�p�e���`��]�挦7�$3��ZI���T���,�X,����v�������S�_�t��K~%x�8���/ղt��(�j�^����Ч��|PA���kF!/��7��ALW�[2� �mV�F<�Ep�@%bH���D�ܰ�md�`��̂�;��F@[m��B�#F�( u��מ��'��B���a�?��(�%rSRP��~ϓ�F3�%As�������8F�"�e�+YC��:��j�P��6�*�f�׋a��%�N��C:�෣��
����	eGL#��˚_]��r��h��O�2gM*5sR*v<.�����CZ7���U�ajKq#zt<x�)�����r2=S޽��
	z_g��������I�tPcT���j����?<�J҈($9��)�N"@Z���21�t�r輧�a���ogO�Dziv�D(�pŻ5`n���;p ��_�mDv]�Ӧ��"c���v��?�T%2�Q��8��h��3��2SnCn�u{9�E2�m�9$D�ǥyKHQ����0�8�M�5w[]����*��0�%��-�}���W3�mE�(���l{��"��N�E�o.��X��� :�0���/���н�U>픢J���#Vh�רE�L�"	����X�mݶ!Q�'�k�(�uC�ӣ+�v��bbƍ5ҙ��#�hx����9|GG��QK���1|��!v��w=;⭼����fh������*��|�R~�xq�Cj��L�i_7s��2S���w0�p�eҙ[�<|�(.�{I��q���j�L�ߪj�CO��@���͖Ƙ6oد���[T�p4�M�w�o\+�9.�7�0���;���ڸa� �~W^�D-@H~�L���DMNL�T����I�ݧ�=���s�gQ��3&�"Xe��iLL�L��X�Y�j���'��Fe�|�=����k����C��ԗ7���Dβ�`��&��+��Y�zn�K��J�{-8+��>i$�l����=e�tN����mNP��|M������ٛ�B��ֳ0H�"��Qf��9�}�7X>�ڍO�V�^b��IT�ˍo���6�~C�=P�ñ���ŸO �5�d
lۿkz���v#����lt����^S�u�'�-̉���XH�4$�ݲt_�~u�r��w��T���M�Ǐ&n~�噽����4�~I9R�[���7�ǤX�l��i��Ƣˉi��g��&զ
���75�ɬ�ܖ)%k4Mh!�w�'�CЪ��)VS3H��o�6�@���cV�;7bi�u+�$�2���9��T�$|1�����դ)Nh9�	Z��""�O��Aa�}��Y3D�{>u_;.���{A��Ki)Z&��a�)1���^��׋�4(��.,���\��%)��ֆ�p��{�^O�E7ذ��*�v�@H"�7Ov�q�w��j��h�w�hB�j_u.���E�1ʮ�l<L@~v����s�p���^ܽh�L7�Դ���z��N	�B?e(��+��/�/�Q�`�F�v����T�� s����vY�T�	��EG�	�+�K�f�CV�s������a����!����zC��hИ�1����F��kX�,��9��U�&#�Ėx�g5���p���Jm�g���|&q�^��_���}{�,N��|nŃ���y���.y<��������"}�+a*S'��H^�x^p{�](h!�ʠ��n�P��*��l�ަ�;�M택��,Fh`������\�{I�̎S�}��m�?:e�o\ �T�{H4=�s|{�����#�mp�ǣ���XM�B��J|[�����k�B�����*x�.���]#B����΁�b�Z��ӕ��Og�Y����Zmv���=�W�yNʹ�@ԫI^����4�S]��Mٕ�U�KO~�o��T?;7�H�J�����#yO�q���������kkq�����'�z��j�/b��d摡�q��wt�H&~��=�hv�D�\y�>�j�ޒKp��/��F��t�����_��^�`�g�@UamH,t0j��}���2���O���R (h}yE�V�w��wW,���:h͍�G�Xm;W�G
UR��nX4�?�Gr@~o�>�;���6<�>5h���;�$�A���_�j��lT^��yBu�_wu���-��l�)!;�c@��Y�5w	��]���R�|-?��l�|�;���^r��+������!�ǥR�]\������\7�4�E{�s�	m�,~�5�Lt?�
`���4w�dS5{]s��O<�tzx'-��6sr[�#Τ)�9o����wܜ~��l�����b�J�pI|�r�g�M �^Hp���[:��J 7�h ����:xሷ��!-
i���ӻ�؈�!����W��V��}�|�_���y?�ϥ�����)�!U-c��~�<���z�䆛yEY���b�!b������b���A�1;�E�4�$�x�t��p|:��Q�h�^4��>PC��_:DoGcVA4�Y��c���;���/�`�H����m��9�k��Qصz�,W�0<@�p�+L�ؒ�Q�(��c�Q�����%�p�3~I3|{�0�3S8��M ��8�ʰ����Cb�2cq�@8Щ�� byHd�1Z�큋��I�1&��?�b� ���L:�#�I5h��2Ͱ5F��ع+ ��T��V׸�V
f����'�.���d����OŐ���HoV�Ґt�M[�dI���-�A��%�����bࠧ�&T��K^P(���!U�i+
���g�6]%���u�v,+���F���H}�&�ƓDi0�I-#���Ṍ�����������Z�x�m�����&���HD� _8-g%�{VJ�Vc]��s~�ދC��nا�Vtq2�`0��y�����H��_�yu/χ��tM�1�ZT�� �Y�G	];R���H�r(�_n4��mӂ��m�������0�S��: ��pC�huW'&��U��?{��"�������4��'�:2����6{�� b��'�V�|в��/
!%��o��R�~�{�/�:w����ϸӟ��/"��M�x�2?}1Z��Ĩ���:k��7��-��VK�\�x�}m��1�������f��#�c_@����O������L�9���A���9�g����$܍D�8(�v�e.��
�|g�[�Y�k	��Ǵu݅$�c�k��- ����'�˯��%�	;LP}��WWfH�[�;~����Hz2Y��Z�$��k5�o� Xْ�{�Q��L���S�R�TT�X�&�u�)���u�O�{�}m3g��0:J��[��p��W! -�I���lwM(��ZM��`5ߢi�Uy0���w�b���R%:8��|{�