��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6o���Vyȃ��I�L��2_�v�%��=m��zwfq�[����ɸ��E�����'g:��F�	���Na/U���Qj}ć��{���b��I�5m�/�W��7{!95Pn(�LRO#���$��U���+�r=� ;�.�����_�T�u<?$o?��HH0�P��vڡxg"�*̅�{��I2Q�nQ7�m��]�Q �� �'�?�S�i�����|I�������rM�� �
<J�e��u�.\B]�>D6�'�.D|�;l`J�FVZM��~Q�3�6+I|<��.�{��қ��f��;�'f�T��j���`˿s�
����������M�R�u1��q�U�����hF׍��4�=Y"�ձ�_Ÿ́ۙW�KT �/��Oݔ�k��}�T��	�V�v�Rxu���F�����8��n\c"�d�F�+�����3i����01�p�+*�2�uu�&/Ŀ�L꼷���_/�}L�܁�6��ID�&2(��n��|���r�'Fŭ���h8��(�7^ч0BZ��P�N��g�w'G�7�dNo�:J�:���0��cC3�ѿ|G���Cz�W�*���(�.d�����G�NyVU].��^�x����.y�FɞJ��p��)K��V����xJ^I
Xg��rz)0rH����AY����-��C���P��M ̏�8��;�j�����_�D6�a��� ڪ�y�j�~3j�� �����$�/��z^�9��(������������CC/F�(��]��K�RT�p �<���AΕ+�k�\�����7c�+Aһ%��1��q��q�,����4z
�֘�j��тa�������ȕ �l�7�h{�4�k}O�(<t�-	"ޯ��������S�춛e�+��M���'wN�,�x��A)�˸���}X�XbT^489�^s�V��8��Kpm�N-$C�;j�l㦝���R' a��4���ҾF�Ô��.���{9g��a��wY#FC�%謼P�w@|���ٵ���X�ļ��x��a��_�X�	'd�e��3t�BC���O�E�q�m���@���cn�!��Y9�g��U���N������R^|��@�k�3�W�p�:�����&��2Y�0�E�O�R��ygjJY�}��K�~�)��Rd�^��A9�lŒ
������T3y��lЏ����3���O����"�K&��/�����Jy��0A�`�c�f7�Q�ƚ�Hu�1&�A/��@o�v(��?�E7���R/��k<���NqSE�	g���{��� ��4�	"O|PM���3y`G�X��o��b��KP,�m��T�wɢ֔��b���~^��wCo�6�E@�r�J'���U������!%r|V��{�����(�[�X��J:"O6����h�0��#�?M������ֆ�n��V({&M�T���=�nR�~�w�oC�҅q�˹F7��r.$!Է#�qT���1L�Lu�U��K5W�솧I�Bڸ�[��J��䷙_j-����+��}lUԢ�{SUZ\��H�Rx���d���l^i���K專8UI�
��B�����s��#DP��}G������1�������0j����#�0w���3l(ˑ}Q��"��Zj�a]�aM?���x�4���-W(t����j�z�׮/(n���͘�P`Q�u�v�)��@��������nw�L��B����	���Gy���)���:���"<j�㝪K��gl�~o���&N�i~k���73�bn_��A�˄���q;�5zA�����'�-?Z�����V?W����$��$�	���l�y)�|U)��X"�6ɵ7B�M�I��QP=��vQ=H����K��39��$�=?[�� �֗�#4>�vc���fɻ�s��DJ����i	�p8��`��0'��D[�@:uV���/��L|.���ϘSl�96O	X�R	ϼJ��WmD=9j`��P����<2��k [x�L�	�&���
f{gqrmmW��B�QUϦt��N�w�Ȃ�/�%���!ED��0��
)��_��m
���YL�5R��y���x]�˼(��dɐ!�տ��t�d��RL�)�S����<篾��VT���E����hДb����Y��-�	/<��ڣ�pō���{%��6#~`��@�;��Տ'�����\"��C鐫��tpz���(ww�Ro��a:��#b��ls��|SJBxi
����]�#t�lKM�e�`�-	��9C�"�v�����`H�S�i�k���@hl��>�$'4�JVj����&U�B�&Z�On��CS�Y	��Ճa#�a�F�4���X]j�áQCw8.H�\L�*ܬa {���Я���=����f"��������B�!��r�xs�Z�ہ�P;K��Z"M�!|����(�ڲ>��O��IB'�(h��ѥ��w#ZX=#�9g6�ҋP�f����zg�	(��w�T�U�n:p]��>� >��jhv�ʉ�X;����>��2˒	7*���X����H6�m��G��,�eP&&��V�ؐa��;%��fj `鞭bVV�C�n��4���8} �9�F���j}�g�^����+�k
�,T�����A��~��K�9xM��M�k"v��"���Q�9������V NC��Zb^y�6~,sJY4gJ�%{��Z���Q�&r;#9?
��$�18ml�7��G����,r.Ƥ�I񄩤0�z'�S��o�X3�_=K�� �=��W2U|5����H�ۦ��K�L���7W�[����P�)_@I�>��kI1����V�����IȕY�%e«��Ir����V����Ϧ��Ie��T�"�Yd��MM���fn����ߣ��/W��KL��/�(_��,�qx�B>�2��j��p�����X;/��j3fQ���Tͻ�~���Ɵ��8O���R4�
��Ag4�.��8��$�����s��ڑb}�����K�)]�bK�?S��X�
�pp�VM���;�83ͫ�m,)���ŴsZ"%��$.tV���P,���~��z�b�X���q�.}� iib�� ͕��z��=���Mw� �#�F���?�/}�>�D�?�e3S\���"5��=7���B'�=u5����!6��ߓ����:�媑/�"��9kS ��H�J&��$?�kpδ�Rl �Qhd��ҽ�r>��ې����j����I#����+US$2!��LQ%v�n\L�=�^�h�n�,m
�A���a!��}�.��8-.�F[3��/��]�i"c��Ɇ��b ʩ�R굝iu�z��cS�Q�(�9� �G�|#��ѢJ�3"�r����֥�iю�e�L�F��޳��hzG�R�l�����$���׫pW!�q�e��a���T���a�P���1pe�<0g�x�edO*�7�G�e��m���ݿh_�n��H�1�vҸ��>-�ؿ�վ��.[�L���@��i�����-hT@!������	
�bCx��$�E�&g��`�Ȥ�Y����"�ǹ������J�郊e�po� :��1�2�do�O�y�ŗ��562�(P~��0�K �i��1�����f����*���)��[���3E����t��m4���Y��6Ҳ�JG�e��;�\68RЊ�Ў����_�$�hK�(pA�ϕ��n��5[�'^�6���
�B���K�D�̍͆io��zJ����,��~��k��fe���D?]�>�x��ZO��~�B	�G�P���VzC�)]绵�{@Z�~n8������(�?	юa�pZD�`v�A�1�^6�@��篅 ��U�k�珯\�4jT;G�0�4���K혪���(널[Cs���,[����@bء��ڐn�y����i���B�5�:|�X�o�0��0��.A���~�8ٳo=��E��U�3.���P��*���}do������nf�3 #|�W���eF#g��
�z�o6�!ȯ+�:���X��2�M���
F�3�
�~%�q8�\FMo�hY��Z��C;�gV(����ѲB��%Ey��C4�2<9%����9RQ�Rߢ�8xqʣ[�Z
�����U�vZ<%�΀��*�g��?U���9}�V������$��WU�\_�0���'�yB�a�2�tx���	5":��`��~m�������_Ӽ�0�m��|߇�͗�*�y��&����5��0#�C�/�J��:����ZW��-����`ɡ�[��	H��
w�d��M)�� �(�]s����F�eL�H�|���k9M��2���خ���=,�ɓQar� �]����G�)^/\����(�Ţ}V�w!�Z�\��:3r9f;(:sn���7�v ���o]L2��0g�eFd�F��W�ֲ�3ebr��I����_e�pN�!3��\E�&���'c��얾�c��n*���77����Y�(U�u?YlA�4÷�u,K�����7α���40/4Q��Iahp��<���K��F�2X#tۋJR9���f��Z���Hhj�
�]ҫ�<G�PC���=�4k�S$���l-�mx�pM��� �F4�����
�#�s=�5ڹ����C��w��SV��0a�)s.$]&�ϧ}ǚ�(�%����]�N$�@��R�9o�d�7.6�FX�n��s2�?fZ�A1'k&K�����'�<�����d������c	ԣ"�VA��m٣��<�U.9�8US��k^�Ɯ[^��q��j%��]�hԎ�-�� ���������UҜT�9�	�tBN�������`�6?	�:�8�Z���:gv%��E�������t��3�@��%]�5��hN�7�}�)LK2��(� �� �D�������ʩ���r���6�㕵�9�[ 4k��ɘ�l������
�� 8g|eh-�K� ��6q8�z�CH�Ӓ��E6}�<��i��R���y~À3d"۰�_x�]���\��h,��jE����6��z7��ޠ���#�_�J�0�u��{B�����  �Y����#��NhFf��v��; �nG��Ưp���	")�F���1������(靲��|́k�F(��l�l���i�)M�:����Y)=^�/��� }�sE��U��3��r�!��������I����Qj�T�2.����Gu��N��Q@��1��k��Z���X�s��/��ձޑ��ա�LSX���Ѫ��%�i�	]ز�6� }�+�G���-]'�
�N�O:�ZM�6o��θ�z�4TD}������W�*��Rwy�<��¡z�>FZCP->��Ւ\*���VX��m����5@��O�b�e+����Z� %1�E=��4����-7(��	����b@�?Y_��aR��b�=�]kϏ��1g�A/�o1���޴9?g���!k�����k�(�#�>z�16��a���,>Z�3��p�l������h��2���/n8��Vu��xS��R���)�_N4@�ע(�D�!�h�jJR�z������F�DZ%'7��8��x�����ʷ8�ۅ��  x���μ?�ǭ�MT;�WZ!
���W��D�x�dh_���+-��|����e�D8���t5��k`�vCٰ����u��(��A��Ч����.��DRpU�3�=��4�̹��t�ɤ���x�*�]/���BUYp�/�&��O��\��e1���#�l��d�h��'��?���4:��!y�8�<�'�e���F;s���H�WOCq�%�d�ɓ�_}�
֕�;�.;d�d,�`�w�b[ؓ�Iͨ��t�Z��(�t���# �4S��ԍ���g�k�tݟ�.��@�?1P���qC������&�[�h?�� �>��!�5�T��d@_=Jԯc�-V��I��&��Ԏ�zV�y���+l#��t�VR~P�>Dz�j˭��b���@v!��N��+��9o����դ\�hLԩLG���D��j B ����P�����q�I�SD&[-q�[5�:�4��]�,�&�珔$n�7��p�&�:��vp?�/ch.�{����N'WQ���{hG�5ӊ�֨�\J�^���S��j��7*P͈���?���ؑ�m�!�łb�k/����Ne���ZƉ뉂ճR«����tz�(t��K�o:*H����'�x���ܢ�Aէ���1��FX�0�),�yy؄����Q0���p�!m��: J��T [�	7���P�� �71��[� 4na�o��ݖ.Nv�1��袀i�����Z�[�?�Q�Үڐ�7Q�_��9aQ䋝���(6�{ӵ>��?�=X�v�>���x}����(�"P�D�_�.n��j��q���eqK���6���-�EZ���$tpH�2�B�R�$t���|\����\A|�R�/��B-���ev���F�f�zx@a���{IAsTbDqC�M�nO	�����u���L���JL��?���Aj�3��\v�Xx}�N0c�-&���4(��-��J�Q�����bl<�@j}�+#�"1��l��ǀٿ��@�7�q=��_��@-�[���Nr^99�d�	3H>ԡ��%/�h��8U�ܹ�bm�/+2�7��N���Q*3�'��ҥ�F���������eg\]�,	�?g��e�`n9!�d����էy�\-ԔA�;�%��:joet���/���6����`�����*��;��Ƿ�e��^ā��A�ܶ��P�i����ïC�,��x�!�K.[�B�<��}�A�z7@�˜��9*�C}�c��󵌜6<1�M'�P�nEk����A]C�-�di�����^4�� 3�v�([V(6�
�ɝ����+�`�-�L�ἅro����w�>$ЖS���N���x3I^<b�=3��U��Z�7�6i�r��([\:���H��+/�+�,K�hzTA���"�:�<��H�"S(�A��U���"��]�;Һx^D�G�Nq� ~�[Иs��ϗ2���y9<v�����W�	�U˫V,*����Brz�~4����%#򗯮r�ZGaE��양����˖�_q������b��|N�e�v1�������AhE��,��a�-O��b�,UL]�+;�J��2dNH��&ӆ�s�7%��	�{���A�\s$��Q$���va�fn���cjBԓ̜�=#$��k��[�M?u�]`lpF ���2�wL����8U �?��Cw<o�D�[7���u�7h��_�iUIR,��;��F��NG���D��3Xȟ�tJ�4J.% ��2�Flk*���N���h�^�'Y:��C���n���,��"�X�]��_Q�-�wlQ�W{dc�m.�8���pka���e~��>��V�oaI�[^N���p�Ip킧��b�|^Fn�H�m��	
G3���Ͳ`�
T�.��cI=\\7�p�([d\�`T?�lQ�t��群땑�5�4��Ug䲅�DvJ?�z �8��S���0��z����r�c!�~�v��&��r��s ��`~��!~M��%�5��&sm��W����[��!���-?�4��TO\�)���w���c�g�F�tn�����+K3�5���hCT�Q�gO�Zv;�a{�]�V`���$����ӸM[p$EբPP�/�>ѽ�Խ�[����)��3|��=��]�y�IĎ �֔&e�b�=c��v�~���ʔ߶�d�&L��}JSڝ���^�2�H3?r��lDs��i�JíW��Cp�l|=%�_�1#��x���7z?�;܌Ġ��7˪�n6���UK�dJ�� ,�vv��9	tT�P/W�.�
v�Ҩ�=��|���"TY����h�=��S۰ڔ��%P��3�^wQ��� к�#&�U��n!��`λYJ�}XC��d�'��N۲�������o?�gw֊9�6�D`/{M��J�x�|@X:������w��z����Lq�
�,�/�T��� ��ڋ���(�i�o(���垮�^��t���bD����O0z�G��K�Ò�'����/��M���C����1��8�'��7eU�1%T�SH'�"2�vc�+�?�=6\S��ic~Nar��+�����v~�I�q��i9N8����B^)W
�_L/R���k����6+��}���q���Xq�/�<~���vNv<�	P,�H�
�og%
Ǽf���Բ1w[xg��Ç݌�����F8����+�����+ѴL��"KaV͞Q~��������_Y�f�s�?E�+Yܪ�k����v��A���c��?���$EVX���]�z�>�I�d�kM?܏�ӛ/A��!�ʧ�"|p�y��s�4~������/S�����Ը��_��r��"�`�s�3!�k�Q� �=�o=���6�Rͯ�wN�Y��A���et
X���X�Ja/�a�V���yiC�4.����V������-�w�S��+�}�a��~�%�{B����d���%6����~p�����T2́r�h1�U���l�g��"(!)���n�PͩM���4��bQ�V���K�-�Oo 8Q�0�I3a��������E�Љ{�U�X�����l�l�!&tS�Y@�W � ������Ȃ�+{�_�]�'��1Y�ݨ��;�{�쇁\�;����tϧ��)/3�2���p���iZ�Ї�i���wQp/�xm�L!� A�:�fO�9q�( j�^IC!�}7��CE��n�	�!656��q���C�F§��K��q����Ⱥ Lע�hb����+����^�V�ٮ����`7+T72��=���[�;�Z�6���bP��2[��G��Դ������*G�c@N�R.>�VbKp���/S��q>���da� ř湔�;OWn� |E�g���b\0��ҷ��H�L0nfy���\o<9�/��_To:3�^�ŮE�}/�?߷ۦ^B�u�o�}�W�8ꈁg�k=�#
k��x���W���x��~��p�����O�`0	��Z��	��A/��7�+a��� ���s��Zt�΅D��_���C����2��P"�
��\+��%e�a����=��D��)b��I���@��`�@�M�_�]�'�d�&�;sj��}�4�Ë��+��c�~�:����p��u�i��j�W�wO�BA�g�ƍ��p�1��CK��bV6ș]�#�;t?1�q�طå"d#(
#���))�(���w���$��ѧ�X�����8�F`_�}��T�	\��p= 
��V���O��M�7
l����m����$n���J�xb]���h�ԙ�n
�wV����-�q��,.X������趽�Aŏ�����/�8�ӗ�@�(�{�����p0��.i{Z���o{&hI�=2���Og��0�Լ]A�V�x�_?�Mw�4�A��\'h�]��yw�7p(�!�1�3�����q�i��`������Ӛ8���C� ϐ�^ �T�!�C�f1���g�p��p�tV��&x�Ͽ�)mgX�I:ȻL��
m@S��d�����,��J�����>Qv��.Ӟ����`%�J��G0�Y=�z�X@�	���[�^��	���^�nT�fb�����7�Eå ��Ԕ��I��^�B�r�̍�9-���F �y����ނ��Ƥ*'����T��!��kS@��D";ES�E ��6<���Ô��£%uc2q5�M��^;<�X��7L�t@b�)1����Z��g~~�_R�'�����������q���m��\�YZg�`'��|=ԥch��h�v��$,��-�<3%|%2�5b�@��(@�����=~@$*��Tǝ��g��{ d'�+��PE��'|Z���:�o�\�L�v��js~U�+�G>���--x�F=�
0�
h�hI<e^x	�4A����dz��]n/4�P�K;}���y�X�u��#��ܡ�(hI�!����6��ö$9|�#\��+m�C��Z{���I�liQ�� �]OU��1�@��:Dh��^�Mz4�-���	�(��>��T����)I�ųa7�b��.q�/���ƶ�_��l�g�#�h�p{I�I[���b�Aw\I)��Dɦ��O�E��}]�a��C	f���>w%�C�	�� �	�Q�D���ഗN$v��:F�;����;+p!/2�*5LH���:�oz"��vy�����6����gtP�3V_hd��FRf���ω[z�ĎS�ۑq�
�b��ػ���x�m�vhV[!�*#A� n�ˁ�.Ds�y�R3P��,ZJی��\�%�%S�2x��8� �2�A �&B���}T1:I\�>�~h���?v��%�҄�)\�-k��>�������ȃ�W�7%��?k��I �:��B~�@��G2�3Kr.�"�ƁB��Pg���5>+`��y��x��*KC�?xvRA|8�JR�]��Ɲ�N�r�}B�T�&�h�R@��n���H�8�,u���~���Ʃ2�f�OXZ!1茩�}KP��i�r��4�<}M*BP��^��01����������9�y�g(�p�1�&��7��;K/�=pU�"�V�h4Y�At!^��:;��u�FPf��K��7�瀓��Uw���;�}�������΃�#���#����~獷��l�+i� �pK��� ε���78� 7*뻨,��\�}�BB��0�[T�id_���3��U~8�) p�h���tص�tۜ�M~�㱙Ɛ�`�C��٬���Q��o$v>���9��zhD(�Dr~�FJ��id���� P��YXg!&�n7��������B-��U.�����A5�l��ʨ�<$UMHd��s��(5��m��'0by��ߞQR!e�x�u��wU�G�ꊶ��?2��� �Ӑ�AQCVm	�"�t���������1���2�(�)I4�Ի�xf`='�MqR�P+�x�����:������^%���i����ƽ&��;I���&��Q{�m^�dē�^��WE��}u����{����NN:]`��M4��B8>�dQ��{ܶ���+eBXyr�鋐��JdaPJ.�&�86KyY��E�Y��a�ޱ��?e�3�ٲk� ���B��_I�\Q��|1�����Xk@����}���Ǻ��B��3`�J|&���)ΡO��DBwv��kX���=G�l|o�IOY;�w��V)�1���T�p���‫����K�t�Nv������tT�t<���HF>5�5AgI�+#v�0>��#���b�p��: �����S�:lc���D�j��(��oa�A'�mz����$0:�]�:+�����!�u��%�X����:���l#l�������)))?�-V;�[\y�\فÈ�d�;敘�Z�e�VϦ���(�r@_;�r:m��U�H��-�b�|ߧ�W�r�e�wE:���2�d�֜(/I1O���5A)�Ԁ��ئ������̙${:�L��sˤ�D��A��d�l �klĝ7T�e�2�ѷ����8gӳAb�\Ӧ7�ek���q2e�<�~B>�Rw��x�	�HI/���[_V���Q�hg�j,s�-�ܽ�wUaz˰�p��cA��7�2��A�{7�(_�EVř���T���O
ŷP�����e��}M�p�����E�$=��>�{r����;�|G�����l4�D��%ѥ�6����kg�H��e�P���5K���꒑�JO�TS�ǜp���J�]a	Oݜh��AQ��:�g��� iYC�Wp��(�j߀�le��։��������X��\*�r�Y��yC
�ʪ�:YW���cL��z+���C5_4nr�+#6[�A[��_p&�KϫBi8�a�؝��k1�J�:���*OצEE4��s�Mc���1�8t��v����_G�t��-d���k[�vC�wp�����ۺm��K�~��[jvG��*�~fA
9*����p����k�$k^�#��v��[����n�=�WV�3�t&%93ȱDt�$�5�߷�p�@L7�\
�2�T�9[iQw�C.`(�s}�����Y��#���u��Q d���5����F���r�����]݌�e�8�АRnΠ՚|��1�1Q최- ��c-�.�k���t��ڥs�ˮ^�n�s�8q8s���B훗=n��GJx��NaP��
G��cQ���W3���yn%�'�k��q��:��2%�H큋��<O��<"���{� ���:��
�@w�'�ؿCK~ѐ֊�� S���Vl�S��R��kLϙ��4�}�y3gMhh��o	��YW���^e��,t�����U�7�8�3�>렳'eY�7=�@4>��5?�{�uT���-����G�4xx�w�z��
��n�0����
$�,����� 1/�x�w6z�^�QY�~6Q�"�� 5ԫ�A�&ǔ��n�pdPW���#��pNuv/v�K
��O �l&0�+XL-�'�u�΄�!+�nOW���
����!@�aI@�e�(��K0@R����b9$�F=���1W� ;I�6y�����s����-.`3RoӝB@�{�l� TȷLܦ3��m���m�~��l|}�^RQ���ȶ7HF4����2��#���ɡ�DE��13T�R�#"aP�EA&%��"	�4�v��0��%N��g����&p%mB�G�� ��B��-�jP����gFu�L&�B1t��
���|�S�KlJ#C�tV��{tG1>������w�;�m�L0����(�#��b�$��q�yq�f�^7"�o����R��!���D4�o>�o��o����[�{�|ݐ�|�pwec!��DY�L�y%�{i���cٗʐ�yN��������W�M94�6������/gX�bJ_�����l�|�$6?�@}�	[�B�s��p��뱍�t��U�r\>�)�p����]��RU珍�d~�E��d���wpj� ��v}����Mvh��S��c������:6<8�^e�0Q�H#H�/��̀e�L��{ʌ�2�����y��7""�&�_*�y�H�7�Uy�t'�G���*�f�
D��*�Wc��^z�U�ܣ(�Q�K�e�3��b�Rǡ�l!p��#Mv��+C�ڿ4m�(���1ukTtX� ���fKU�0x%���D�t>ִ�������i8d�a#��=���S$�1�K�p�Ә������Ι&ε��]V.E�Ʈq�iՅ� ����w�v�e�e� ���W�w�����g_3(��wQg�U��3�ښsu(qq�Q�!Oh|/�Y*B$$A	�(�I8��v)b�\~�#����SW���r���W�������_�b��+�:p���{G)��\A(q6�uM�>���5N���H:�D��@��*��;!s%�@s�sn���
s���эᎽϳL�l.�8�	cfV �|H��)!��v��^�l��@97��{u��S�jZY������ه�U�q�W˔m�[m����'��*ǯ����*,��^ƙ�<��>ݞ�(�:F��tu�1��}���b�Ə�R�%/q,(~�x���㥧��{�r.ZՃ�o��Y�m��H��p�-�yU���2��Jp;��	oï�� ��ǵr�L�`q��kC8����鋆�I;*���ѺnMU�L��o0I?3a<S�C���8\<�p�?_U���T"^#Q�~YѺQ������!/t�P;���c>�4�gW���^O�l����xu��/H�ֽߠv�����pU]��VQ�H�z5��-5GK�8,,�b�Iُn[Ԯ꼈�j�]Fw/y�V�ㆱ��*�{�_��K�FFH�.a��0le����?�72��^�$�4����_2��p��7������y�,�Ձz��٩`����.BS��h�*�s];<���uZ�!�>���~�c��k\���2MI
�y�S"O��&'���
2�cj�讅sV�/�Q��	O*8}*���KaY�/���ǜ���.r��?>}1����U�m�Q=�tڸ�ƽ�UX�jگX���&َ�>wg+�H��>�y�2e�6vP�<^�Z2\��-1��	�ꅵ㿍ztc�o���W[[���9�?�F~;�>�X�D���y�B��Hh�v�'6/�M��m)ڲn�t��Ը<����hX&ߕ����/�8�=v���̺=�+	�؏�փP�X��"s���m�tF�+����贍�d�S;C��H��0¥�nl_�١����;��Q��6�r��uU�s_�sN�q��H���#������aҪO�|d�E-_�,^�c������-G�Q��|��J\�-Q�@���'ܖ�v�A���?
��r�T7/<5�ԏ�ŨH;E��X	�H���C���\�{�;�;	�	�]1�hT��x��Ҡ�>��yQN+�'k��� �ܸPr[.wg���?Q� [�W� ��/�<,�Ơ��h.)^hO4�>����<��; Ԁ��&^�eD��jT� 5��J�����΍���/�o��y��ӝ&��r�(i8�n(~k��Z���W𔪑O��8�͸��y�� �;��ޯ<�'n�:�f9,��Z@<Ocs��2{�C�S~B9J�6���>��	<=�O�^D7��T:GRXIo��_�����.��ȝ-=BD�cp���#��[E��O^�L��p���e�ū�fU�
u(݅P��{ ��^?_�������Mnvۜm���}�q]x�jW��g�;���k.�;M��&�C��u\�w�
*B�&P�7 ���҄�v��j���!����Dh�R<��h�"rW���p�J�Ǖ�	�.?���6h���W��i��5�7?>k�C�ꊽ��^��=B� թt4�w)��
|��R�7'�����J���e�Yju;��O�sS�#�ΡP0���Xq����<RSw4��h��b��!�r�k.�T Ύt�����PbAݐջPʩ[B�
(?ľ݋��"]K�`�2I
�ͪ;. ��%��w�I��vIj�_�-��4~>�G�o@�������O����T�A����pdǅ��Gdp�4@)�gY�h	��<S��x��v�?��X��������&0q�1E�p�%�+��s��P݋�9KX�)<����m���_�����ͨ���JA�-o����S��Y<T��p���=��v؈�h�0z�8*�v��h��zN���x\+��gH�sӦ���4��n�͡Wb�K����щ�_#{g�l('��W�*d�/�&���Ҷ�O�~>~��l��u�I*��.�nX'x�ha'I�U_�G|�
+ v�d��3_��LwK�m�c�g���ƭ���E�$�J[�gHUj�A�s���N_���u�M����[E=u�v��1�ʋ��!�S`�+G��
?v�������CH�?������g�z��7�"�|��A\t�����Ԡ�ұ��~��ؙZ��(��]��rH�^�L��@��6����՜Z���p�����m��2�u�߫D���ɱ��hC^����l>o-�h�<""�.�1
J�G�X~�|�{����T��X5�I��V���8S�=���
=�R�(�'�w(��D�� ,��M^d�26�7!�[�������������.�I��b������ѕ<k}�ѫ���:⛥�r�®s��#��2���B~�ƴ���C"���,�I\�s]Kb��پ��K�㹳�����BkSN2(��}kS1[%�g��փޥb��p���jC��g�ޜjH`ˇ�h��Wv'jyUh ,�(E���&�!p���be�j�C�r0��J#�귓%�8 H&��_�2~�r�C94��P�n��!]Mł�3ץb<'��Ś
Vm��X%�h�w���h�2 3 h^������CƝq��l����Y�pЕO�,=!�WT�e�/b�#��Χ���R����(2��z�5p�k��tl#����X1��N^�L�42��i���;L
���8�g'��p�8���*�%��}���8��ޒ��2?�O���٢/o!=���C�#U��$�_��z?��ФC�r��&1�Ձ&���s���b�)yj�^��RG��d���g~ߒ��ݜ��h*�8 ��()3>{.�����(	 �`J�}�g&Z�P���j"�-��f�ۗ?�ZW��=ß�i���~�C�k���ےB�c��ʾ)4��t�:�-���	7Џ������T���u�5�?b���-r6=�88a��e�ɰ����8q�"J�O^_�P�7o\��p�0)y����M2��X�as�&�,��Lҕm��?=)�@�~5���ɼ\I�6�bi��	�:���>�i[��}�Y�ɓ��]R�u=I�o�hX��"�"^J�T��N�i�]��*�2
4�� z�!�@�E�^���}=��Qm_�x�A1V����� �@D�
h�K�M�
gD��e��z1����E�Z�b�^h��D���Ʋ$��E5k�My5��������F0��F\C3�&� +,֓K��^���ܾ��
,��2>� �%Ŗ�����Su�^�ÇX�}��j�9g�J�<D�̨ռi�u�e�U!�^�m�C ���R{��8[��+D��(d�H�F��v�GM�Q�W�;Q&��C0���.(kwS����q�:L��H����m�g-�k���ܶGkL?�+C��Z?�	�z�Z��N�@ĖW��@�dK|X���X��k#A��Ȟ��lYP6hX>��y���,�|�`+�����̆������yG� �a�[�C���Z�`��J^�C¦�*�6�}��Zq�
� ���O�JԲ�KI�7\���μ��(�g7?-.��C�x�Y��n�Ib@%�U�����G��7��1~4|�5��=#Ù:H��nE�p,gu�TeH���kSB��h���`LԾ.���������QNȧsZ	�v�Py�jb\�gT0��]R�fK�Zh��f�1s��[��Q��	b�R0^ L9�p���'*n��|�v��� (� )�}4���)�V�\lP�~_�T��w���{;���GQf!�n�#�!���*w^�HL�V
���u!� �\�.I<���հ:$<�Z��Tӝ9b囵Q��Zd�z ��'�,/>~��h�F���]K; ��^��L�?���5)m�,%��[��|�J8XV���a�gV?�U�7���_ ���ߧQ��� Ue��k��*��$�a.�,�r���������w�K��N>>ȇ�Ü[�m��o	w�v����� 2���b�
'�c�L;�w:�t�1s�̻��nu	lj��8�Z���bN:�ݽ�(uru�ka �J���^-���馭u���V3�g�A��[]��G�D+�ݴ`�mnf�� �$��7��s]�x͒{F??t�j"�'e�C� �#��d�3�z �]�����7�o���H��Q��a�#q^�Tz�ж2CD0�\Ty�c<Ҏ����)R�4=��3	��;�(���9B��]D�y6��{=V�L�^��E�XT5�S�B�s�rc�F�P'�`�����c?����(f�Vsj����ͮ����DĂ*I:e<(AJPP��p��m�*nC)j�s���� �4��$�ߴ���}Z�@�῵+Oì}��IO�2�fs��\�>�&��M�ʯ�v���r���v��}��_����q(��M_vQ�٣����У�{��m)���<[+�TW����u�[�f2����;�\?��T�5��jʺU}K�C��S�=�]��
�a:_^HS��\;���8��!t��_�K:�0�7��\G���&,�%.�)^"8�'���g�+����U�%�����i�1����j�9�Zm�ʃ�s6!������Z�z�}��^M��L,�~sX?�&h=��,	d�+���rz%���2e)�0�0�d��INፂ)���"��{AboJ�<B�Uq�1�,�*�l��G�x�b8 �`Y��������f�<_Ҍ�I�6��=U��9�C�0w ��_��+Üe�S3j�!$�}D|Ap)x[�c�"8��@��R��xJ屛��cE�|E�쳄�}:�vq�c(�T��[@}̧Lb�&�W�<�\��%R?BKNaEn��n�����:w��i_Y���N�D�c'W�5"(9�&İQ��q z9wC fL͟�}DH �����3��7��\D\֣��eE���Q��m8����"q���%)���v�Ya��d��k.*K�2�NEN�S�\�2�E/�HAG��B�;��m�+�,��oq�q���d��9f�D&�K�=�塘��`�-�s��yuaK}#|d�*�d����c��eȪ���P��
i�d���vCw�.�jT	���O)�Am�bSl�2�0�Ƈ�\O���"�&I�fd��L�{j;�}�Tt�ɜ��h�������ԥ�߻�,�
�wъ��{D|��퟊-�?ȡ��C��&n9">�֪�����}q7H_VՇ�U�~�քf�fD�U�5D���*������)�������^�����B!�����P��pBP|I������#�K�c����(��T%�6�{k�nC���bE�oe�}΁q��\�U���~��~#��pNRÝ�N�?4�*�Ja`�N݁oc%�q��F]i����1�l��f��pi�?*%.�_X/3ce�r-� a�J\�7�4D}�D��t�*-�Y�[[X��0B�����tH^�ʑ��{?��T��g��')�
^�;��C��Tk�٣��%J%���u���O��ܪK�;*�*QמS�@��]��i\9���/B<+Y�a�y"�e�Qr�g��PJQ	�wy�z}Un6�k�y�:if��#�~�ܭ���O	�V����iލ	=%f�!��]�2�h\Z��9!�l�9�kLsv���h��	Q�@�y_�r��[��G���+�$��fކ�yP2JAT�ܤ�fG���J���v�WF�������O���ݳ������(����z�H������6�y0�Sd�h�'OK%#2����`(FFY����Xh8�\��/`��ածA�`i,��3�@Y��An��&��3����=���F&�o�v���K=�������g<�(��jGZ6�U�_��� �T���ٔ��9�ih%X�X��H �S W�l����q��XJ3��d�#��Q�Ѡ΄5�2AL���a�0"ύ1�V��]�̴e8���`�^���v͉2zk�u�\���vVi�]���(�U�3���G�L��[��� �<�a��gj��l�.b��g\aюr/��92���m
�D+�fκ�u���-ԝ�<=�V��<D=C���x��O0���,����$A���ak
k)�o<��G?w�����j^h����nON������ۑB��Q<��曡8b��Re|0�D�5�(@\o�M0�?��9��2�����b#���C$<�|
��,�/CF6�ˠt.�hx�)݌��Mi�3̵�tb���[K3xBMzߝ���{����'fnNX�7���~���h��)3w텓p����㶧^���^����}㐸'g]>��Q�mV�8 �ە�A�I���� |4�nK/Tt�w�� P����m%���L<�x랸�hɉO�Yt���f!Ѥc�/B�+��3ƽӮgz@kCE�C�,6۩#�	�N���_5W��G;�I��"�u*�Sl�+����Db�:5R��ב�{S�Sp2�7�	�p f&�r6 :,w|���" {�:��=#X����Ƣ�?�6�]��d=]Y�:FJNO/��vs������	�[%��]����է%k��d���!C�وM�����{��xhC
�B����0�����B�q�޽�u9cZ���v�C;����e;ɜ�����G�n��3�����m�[�涯��Qa��M̀鐉e�2[%ZR>�Ԥ!S�cn�M=�y�k�6`������?���a�l�Uv��^��̣�j���P.7��{�q<)9G*�(�uw��i�k��xorIN��N�%���ӭ��'s�D�)�v��,zK��FC�ua�]vg��".����Y֝c�f��2��prn��7���%i~P�����+r {A0�*?�e���ODֹJ�ؽulVU䋯ß�'oK�d��6���r��kD�:�i��y��ڔ�OrMM��o3$]k��,@D3�"*�	�����a��t�ag�t� �7��!�2����s^2܌ؙ]]aJ��|��b)IC��n�a�NT��E�yE�X�h7��ڧ�����vy�9/�De�7�M���4c�΄�F�`�.D��t�4ҍ'��N����^�8F�^���{Rc�-�j�$�y@�5�B��Ȫ��h5�"
@rv<Υ�b����,�$�ѷ�6B�:�.G�2a�6.�]�(Dy�c�؆a��>�q堩�{:3���<[�1�6"�?�S���"1ÀEQ�����ݪJ�l���|��J_����5 v�%�91�ws��N�!iU���5#Ij�b�-�ȶ�|�h�u��?B�A{����%=-�0B6A�dV[d���c�?Ye��#�`+��!�	ME2����`����ً�'1�@�%`;G�� 5}8:����yB}����Qp��e��ډr����䱊V�Y��M=H!�Ʉ���P\��DuM�)�,�d�W��G�,>��	5�d����A�4��DG�wW��^9�ׅ݂a����Vg����˩~�p�Ux��˃|H�k�U�^��1z~�>�(���<�~���B����c��ͨC*��8��nT[�1�YP��V���,�`
G'�a��Q?C��)�(VChX�R���s��Z$�"m�ȯ ���d�R/�jo����c 7���$�m-�N:wɉ��_pA�Ӷ9/޶��n��i5����@�gժ��u`��A4�`T�"ȵ���eI-����U��#��qEZ6itp���u���X~�7S���_��<�Ʃ�vڪX}R
o��:�f ��%��S�h���'f,n'����pӓ�T�ߛ}�ڐ�LP��'`�l&��\�T���J���K�7�W]�~jeJ\AN�0�q0�����z�2n
��Al��O�?�`!x�-�/Ե�P�-nJw�F0p��-���2�|�6܌�)(ڃv@����M�Ϫ�$��GZi�g��Xk+!�<��G����5��9�_�B��l �i��p-��Uz���?tU�r7��*km�UQ��1�p�wF�\�XJ�ڒ���5o$��t��ƴ��G�f����$��w�3ÁV!�gI�71v�Ą��ۡ�kJ��?Y4d4Jm�f+m��c���qI��-Yp�!��;���Mғ} TP�u�����MhM5xE$�.�
QI	p����Ү��t�zV���,�?���AA���,���D��,e��Q�Z{�I��H�w�	�N�Q�g�r��mz%'�����*��$.G]"v��ś�G�~�����#�[+6Go�(�(]Rd���$�&
��L#yҕ�š�B<�
:'�;4�u��w<�Y��bI�U��S`W��re*c ��`�	� N�w�
����*�r�����#��qU�X�)�ytaP�V�ߦJ��oMN��w�r#ѠD,�y��ɳ��v�Y��#~e���6�ؒϖ}� ��R��pK��?M��KH�,A8u�,R��64�E1�D�b�*�#��;Un-��>I44;��ycR�$z���ɚ;P��U�h��i�/�2U*����r剟_<3��8���^~m�o3p'9H�$�G�R]c��/�B�#�;�����
�8�)LR$�TTb�@lox�o%[c6�~��q��jr u��u����6��:"� @p��g�*=�ۊ ��cg莙}M�_=�����o��9B�&��o����������H�e �A�X>?����M��!�M�n람�r7u*h��A������P���1��j�� >����Ц�}!��bǪ���ZeQ�4̴���Ύ:Mj[�;#��TymCk��\�/HE+����H,� ��)\�#�ISM�����?b��TbY�uW��n��kCH�w�6��eaJ��oJ	�R�-|�n6|���/�K{���pEݾW�?��X̆P �恬�<[q�9復�׆�n����
�Ijt?���x\�uO�yE��c��\e�_�bsW+gc�K�^�/�L�0X�o�o�{�97 B���CI�fha�3��a\,~�ʈ]��	H/��xOnP;>ROnn�U�y��D1��i���A�|�ᅗ,���E)��#C�F�基���q��-^0�h���~f۔�6���Vެ+�v�S���Цu!�7A���rƺ|h�7�c��M��B�yq�
�ƴ�<���� ��jKv%�\��K2c�"y�� d�厳��T����(��En<�o�\�V�M���!t�_�z�7T�8jn��6A�*PcZw͸��{��vZ?|��	��%��"/ܲ�x(�1���~��X@ ���~��z�}[��sG���X��y>]����g2�h��N��_q�5|�ׁEw�\�U�5����R�X�+$���<�+���mA���Ƃ��N���Eh��^_z�Î��y2Յ]v�D2T�0��.Qk�>��z���UB��tNC��|Wr�+��}�ylP?A�����V?9,p��̌���yQ2�!6�T���!�H���'j3�*�B$�:�{1�$���������&��{;7RFN�t�*�T�
��i#�h��_��z��84�5�vŬFD0�A���
�F�$�V �|�]�)�$~�;����mw�0�_e�R��<�]ޗ�ˈ�lch��6-��?������f/!M�j~�����1��x�39����O-��D�^�6�/�k.^��1�dڷ˪�=��&�W^�HiԬU`$_)�zǱ�b�䳨Vy��lR=�
�92S���	4��<�r(紹�%�ᴪ�lU��VZ	�bЀ��W��7Øqv>Oq����R �rU­�(i�^�h`��qr�b��u�K��`�B��wj{S��q��"���O�\�����?e(}�+�p���Y*8ZI�8/=x(�������Q�HZn)%���ϫ�3��g��ʦ��Ec�H��KI�hr`r]����Ty�Ƴ���)�Lj���S����(���PQ�����ydw�?�QZ��=}�a%�.c�fy!�x�H��R�C!���|:wV���[��(�k�B�xz{��DJ��,�>e�e<S�_��O��~�4m.Y/ �����C&3���.�v3^��X�99}����l�z�����G^��]/c_����ţ�D�L�S0�%�Y��]�?�}4�������|�G����iC�l�氖�t\�	~ɞGm��&����γѤ��T��L'��Z1/�v��g�#@�6\Y�҉�Ʉ,惛���`g��7�3�H<���Ԓ���?0w�m��L#�:���(M�d�����<��l0�x�h�A.gN6T�M����^�-���)�V�<`5u�#Ŗ�q�w��Yw��!*��ܬ�31���a���_W�z��M]w��W�G��wrČ6�"�>�ش78���,;���r�qUG�x��W/FKW OP���U_�Pq 7/���ˉ]�%��+^�HaA��pD�{�s�izR��t����;x��:)�)���5~�Ӑ��"�$��,�GQ�UO�����Η���~������[�Si�������+��?1�{߅��ϡK���oKW���8��x�r�)��pA�D���?e�r{YK9����� =h����,��0�Y�� �t.e��
�-K7�x������(U�I8�篼!�J:�_�|�B��-5��3x����KW�U)�B�M�V�z�����Bll,�����B�ThN�M�%I� ��̜|)����g�AR�R�hEB~�[~\T,Ь&6�w\�bq;]Ź��T�ږb���s� Y������k ���â�a�u�=��,��6i�鳮�ͱ����jY� �+�8S_7���퉿 [;����h3\��Jou��>8��K1�n?[�ω���"��J1����)�Z�^C�x�XP*����
-��S.����zXn�"�#K���, ک���V�ݧ(^��e&�[OG��V�6 �� �XikC��a$�%���8j���=��{��U��}@��,�%��E%
�8)1�0&tW�t]^�1(�zM�w�V���i?[��J~�w���2A��Nd:�:ELO��R2Ar�6vĸ`��	�U�HnX۞���E]�	|/(}Xc�׍�P��g��n_c���Ȓ/=q٣TI�1]SU��4����G�� #����?E�ίV:ʹӍd�
�y�'�Οz+���&�4�g�zPܷpE����(`t �6��I�
���;\,m���(�
�ܓ�B\��һ�`��97��z@@��B�_#@����&M�rP����"�G�"j%���
 q�1�fyaiw���?��A[���X�^�Ͳ�����$G��m���"��L������N��0�M�Rrjd�FtT���z�R��:�|�1���E����gm����~����q>�Ԅ�F�I��HhWAl��TeǥԿ���Fs�� ��2�f�yx��ߓ�i<�v���b��)��@���Q�)����[�B�Z@s�+�!�·�z"��aDF\Ҵ�k���`�~ ��d�e�7��߈�%��h�uK3�&<�j4�d��Þ@� �c�ӢNEI?X��@��e��$xRM�ۘ�S�zi��T	��y��\�7IÔ!s�:ǔy�u-ͮ{A�׊\k�����|�	���g6�����T6��	 �cͪc��/7G�+0.�3KwpnJ'��i��xIFA Y��Ex��n�,�A��ŧ���0��R��y���|�_�g�Q������T��-:�*�#�o��[��F���.�)z���˴J�~}�\�К����I��w*���U5�������ǛIS��=��u�y��o���������^��'�kƺ��!=Z�G���(gP/�"�9�z��H��}y�C}FS��_:��O$��1�����L2PQSUB������=�o��s-fǘ���-��O��sJ�A�be�Y�^H���s��,�c6���ʯq��
N�"@X{�j_��e�/���|�ID�|L�C�6��.}
A�1X�5��L��N-q����{D]��_񲜗�uK���i�G_�v�8q�qb	��h\;=�7	Z��tO��z�\����`��&�����S �>�3���Pc U�{�ͻ�I�ɻd��v[���pkG�݄��Ƃ�F���܆	C��}O����� �H@�$��ĉ4I"�� ~W�/w��n����f�=���)p�n�k��ֽ�ؙ�@|	Q�N����L�����$�_����/NH���1�锪�v���|S	����<�c�I�9%W~�s1��-+�����B��
=�Lmr�(O�S;GG��z�+��)鹵�9K)���p���+3�N�W'8mɒ`��ҧ�
Lz1Dc���?��ݸq�@ݪk2<��M���8\t��ͳYE���k ��[�9��ʈ�'<�7�E=E��oQw�#�b|i�3�F�x�����1,�qьXyz8īK���]���G}�o�a���?�Yr'.Bጡ	�0��?�{��,��"ëf�,�_��y�)_T.��I���V�aE���;;ٜM���O�<8�b���[C���
����>4�������~R����o�Z�Jؖ@]_��;1��W�IYc%�->P-۔S�=��נ�%u琱�=�755�Z�3�xc�*�h�iH�e�0i�>��iw�V����C36Hj�E���ֱ�2E"@���jls�HI0ns�L^���`��g���hAK%S(J0����Z���Q��uo�Ҩ�b-�q��p��EH%��(,����S
�W�LGJn�J�S�}���LK����"�Z8�Y�C�|�E��O�Ȳ�wq�,6c4��� �j[�����w��P\ʆ�H�9k)/d��������>��|X���e#2���������
x����%��F�ڼ�wM�4�f����J�V���4*��|�J�-��t����c��/x�}��g�]���2pg��j�'`{�Ji�֗����N�E�ځ����B���0^!��h�Iu�	�1AϹ�~5;�{��������~��t���=F�}� ��p+#YG��EV�f��-�� �`n�^��_ta&�k��f���D*�0���҈�V<o  ��Ȕ�&G&�D�'s��4�2��>��>91N$+���%M�PLЄ|�$e�������&���0HEus4#'3}U�v?�g�?`�W��m� ���O'�2�{���0�J�}��0-�(�\�x��L��9e|�/I���trp�6�i-�~���-r��r�V�y�����Á�����l��jy�W�U+X�:"����f�`�v��M�����G&�y />G���7~�S��3qYن������ph#�QLmŜ���
u[ݾ�9^.�wk�|a�QFTB���"�S��kÈ-��zD/�̯΅��5�ط�l_;��C����5ꦹz�A��s
���4�A��z��aL�'�y2ޥ��4����Zr^zR�r�*�ϙU��	;D� vG�oK�{����%�`�C��<�l�y��{y-%�?��x��q�[�fan�(i"7	8��}XӃ9\$F��.{	��*��P�S�Yl�	�j�v���H[���� X��Oű�����x�
EW.�.H��]Yg��1o���  g�����h�]R��N��hzP9.��\o��D���.�&�k,W�1{R��N���?����S!���
�y,��Md��^��J�.�6`YU�sk��	�ll{Ļ8~m��ؖ��5��r&�1��<�e�n����5ƾ�=�3E�Z��TwzS�
�9���S��V���.щ�bs����b��&W�^mÄ��S�Ȧo�!b;!C�3$�D�)� �P���L
�J��ݼ|f�������B�8/9�s:9�37N�D��Q�F�Ə]�>J�w-�i���_cV�#�/�J�/1G�e�y�?N{���U,�����R�4�����Ssu�7�]���f�Ou��4�)ܻ�d|���?�bE�[��jB��O��MX�%�&�ii�	t�25�W�q��M3C�]5���<+�|��sD�:`�2��O3H�YEH5�s���gp����(��!(�+ˢT���1u��R�y�.E��u���(6}�G�8��l��V&�7h�VW<*���&j/��w����y2������ݾ���L�m� ���,������lyt�\%�;A�0��BYs�g��HG�m��c�%�֤V�!
��ְۭh�g�� �G�;okzT޷r\�^N*�������iȿ1�/-����)5[�޹����O�]��^p@����LE}��i��>�����r��2����ë���Z�<(���tw�ض��N�Õ"u�j2�ev�2M��G�2�m�_�D5�_�W�<�=a�l�������ǡ2(�K8�D3?�aUn�G���9��������E|�J0��P=߰TrԽ���Yo�A����=Ӿ�$�W��F�@��Ì�P"���P�'��R��ou�˰o�ͽ���Q��a%\B=n�6�/�M'W���3�a|G�`�g�vXsm�&4L�2j�+F��B�p��V,��5׏�a��bB�'��OF���765�)�^��̾=�^��os��KC�3[�}��~��/�)��R��1$�k�=!B�;���G�{$R�9L�.1]v�y(��5����@ʣ����n��)?%p���5�Q�y�]�,���šo���ޙ9�1 ������	����6g_��Ĳ�C#��)���a�J]��`���!���X���� P}�P>�Aޥ����2��,��1<i���H�C����>��U B�� (�r��$��k�����]�2���ʤ�ű�les�5{�G�߶�U<�ׅ��5���4�a~��ɶ�
�C��R�b�F�@\:ՄűSة��[�8X��r��72O!�������$�{#���UTwq!'ʪ�H����ŧ�4k�GY�{>�vx`3��E���&xW���H0�3�+�Xs{��v�����Z.�I~���\�T�P'hyL�pj�k�;š��Ґ�1��Ǥng�� OR[���9��)�����	>tT�䈕��9w��������9]�"{�J��\�Rqg[#X8h��q*��KU�;⒡�OP�.؆*�7����Iýiu�����2M!la���Tm�ea�eӗ���Ln_�3�,��UM��0�sC�`�W�:���m�Z�#phS�ɣM�B}siO�J;#->\�2*����a,�|�9lg�쨱Zk7� ��w�*2 �ug�:a$3�<��O&��y��IyV�NZ��Z9)�˿����䄍sȹ����g�&���c?50����v9���h��T �+�F�;0؛��O�s�3�f����JK��,qbFU]�h�n2w-3~��q��i���
�,�s��:�X�lc��Pp-"���Iv�?�n��Oh�yE<�eH{�,��� P3�g�������q� R��������L�؏�?�O�{E���XH��N��^u�~�j1�R�6��x���h<�jP2R"�]@�t�d 唗׮������-@�����=�;Δ)��c3���wGE>���b=������q&�41l��/�:Ԙ��)��"Z_���g������z��/������ �&:ұ�%+#�fO��4?���cD�̠Z ;i�R	�𥉗�Ï�[E�C��0��6�,&C�"��Y2RP��ȡ\
���?G�Y ����r�sl�VVa �
�ީ�UDyy�2O�1?"�uW5�F�854�y>\r�%�Qp��b�ϟ�M��>�Y�B;�N�r��x�?�g�u�����|�C�������>�gaX��-��CI�E��b�����d5���@�q���������/[���#�x�P=%H'T�=��'dS�\�Y�#�
g�hk7N��!(8i�N�vL^y��Xb���<ܵ�G��d��'�-��,��1��������Z&�F\�I�e/N�[KL"��u�Q���&@���3�K->�u0}��Ozh�&0i�6�~t)H�����I��rx=*;�}��M��!J���n��Ytvizd�R���#��b���$Z�h]���ϷkL�
I�V&�Y��uDl=v�w�Ñ�y��YY����m����E\.z��Աrhxo�Bg!Mg?VrB2��Pٺd�e�xl�摏W �8�d�PΥ;ê\��ߪb��8�x���¢�:�P�YN�9���W7w#͏$9^�V�t�Dmk�T�$��f.�x�JI��T�,"g�A��q^J)�5�1��*�Yi�qE_a)p��)S��\8��%3_��ܛ�.rs?ԟ1Q6�yٟ'�ė�c/��=���D�+�������ټsI��`E���%uVO���ZS5ݍw݆��x�)��Gx��x�v\!bӸMK,�/,�S���虢q#�o|����o�6�RO =�D6�%���z�;�fY�@VBZ�[�Gs�x�#7"N~�С�S�Q�t�D�|��	s�柜C"6.r�q��G�Fax�d<���v,����@B�[�s��H�-[�{90;����x����p�8J���$ݙ�_�ks�Lmd�_Z+?�#�Y�����T{<��N��J�8M�h�5,�oB�oͥ�7�@��X,�?���q;�)������^ŗ��`JRB�l_�?�V�X�j,@g$_��J2b�i> T0U�"��>��\Rk���
aþ����[�hR��}=���q�wQBkd���u�f�@�v�$gL�n���3�s"�|��[E�fZg ��h��vG[�݂տ�݄9�� ²ʀ��%�-TK�5�ewq��e��fϋ|���b��9qA��M6��&�[<���_`�7Y��
N��o[�MEޡ��y=����D��bv|����V�Oh���W��g��X��_���� �k���ڶP��]��6�;�`�4s���,�$UO�����������!����y�vԇ��(u�p���E�m���PUmB��+GmA{D�+^E1hT7�2_��������u�Tz�Вi����8x�Eb���I�	�,	Ɏdp�'��P�l�dU��Jv9u`c��D�*PJ�q9{��b4��$�)�s���V�N�������9 ��5\)�F�܎R���J�%�cړ�Š�����(��y��$lW�(�h�,CGU80�'gˉ�,r�D&4�Jw�?��G�5�F�𥳐�'���|��sǸ�5��KR�]�] ~����X�?Ƹ��G�X`�E}��1�D�N�3�.��<���s����~���Im�@.[��׈	J��O.6JӃ�|�y<�B8��9�[��1.���M�J嵢v�v:��O��*bM��Z�!N�#��e��F�T��h�Uk5�{���Ji1��.O�k���V������O�Dn�|n�J�{���f�%S�D�q��v�a{����N��>��&��s)'$��J�[���b���ϝ��'�����ꨑ/�>�ݿ��^�����Ũ�<)UkIe�6	+�"�BX�����V_�l���0ٞ=���ZE�M�۪��i�/��[Ѯ��;�_$���rC<���e�p��N\�U6p�Nj��^�p�߯��0�~�˄���B��c�r�JD��p�x:��lΐM�=q0F?A�����@8�^+���٬%�>������T�#��kޗ?=�.�gfS�����%!�y����W+2���p�5�94c���˔ȳ���Q?��*�$Gv�^���jݨy�Ә+���Q�I�U`�4ޮ.Uɀ����8W�\��V�0�F��M,�i�c��I%�����x���"-�� g�!&��� Y�\���'>s�H!;WB6�4��Z�,T��;�T-��{h�4��G:���m�p�5��pR��n�_wko�A���,e�l��vD���Q���{�՚��`�1!��5����`9{�(R�w!���u)�̎��a�3��k=��t���s��EJ�*;=���kH�������O�� �6�&G��J,�� �������0�� EX�l�Q�lr 08'���\ְ�&�5K����.[��t	i����d��I�"ئn�
�(�%�y��})A�'�/K�P���|�NеPӴ�Ǌ��4���s�H�� �\_[r}�b�h�ei�g�U��W���٥��e��=��1�0�Q(�����p�;i��X���´��.ȿ5�Q���p�#B�wm)��(D
˵9���I2�9��Q" S�=�w	����L�Y��J��{U�c6�Stt�� "r��ٺ"�x�;]���7 �聭9z���;�4�gdF��j�.�{�6�٨�F0��b��H���D���C�h�P�u��Wq�(J�+p���`"oN���B���i�z��2奱/�ک���5ү ����|�֨�T����CP�޵�Jb� ڡ^����T�L�VVۭ�K/O�1�z�r���E�t�-��āց ����QA- L�z�&�^�B���-�:V��rA�WgcS�U��I�F�>��m���9��.��3�ġ��3�E��%8�2d\\~@��cQjߛ&b�ցwь��:_X��>lr(|� [5�f>3[��tArz"0S����eDǣ�3�G��v_n!�2���b >�No��G����R>�8(���7�F`��c�Ǫ���DDcƃ3;ӑ �"t�������c�f��7�]0��4���_��������7tz�!8uǐ#��)C�;��"�����z����X��7mqӑ��aF�-�|]���j��T���P��q�� �j�L���*�j�)T1����On�/`6�V����oZ�O�nA^N���O{�C���
o�eDQ��A�N��9C%���UL�350�IpZ�l�J{��[)H?_'�J�c��KI��jM��H���{�*-�7Bc�XV�d�ζ^��&���D�\<��$�U�F7Y��p�pW8�1	^ع@���E�ɸ~XL�D��Ȓ�:[]��岑]!��K�p��H2TCf��kr:����*a�N���0sK��@����'�4���13	�Q��y�����h#
yd�Æ�h��`���u.���x���{���@ff���zz�3�2K��%�S��f
�J�I�"B{����S��L���<��!d�TU9݃x�ѽ��b6���&+�1(
��\\|�J�~0x<������t�fm y�u��������I�X�&n�Ћ��ċʈ����c�f�2E����Iky]����X`��-�����D�1��ݓ�0�˼���=�ȦO'вÊ
��K��I��������l����=�p�h��Kim��g��m>��F��	�����g|6y�{��5�xf|�=e������Ыǜ�'�BX�A��(�
�$������ٱ��3(�0?�e%�DK�S�@��mH�6�o��"�1yW�ED�z�ɵ��M�}��ƾ�x9`@-~���dXy���;B������.\����~[��d4~�T�E�lZii�W�w��cUctt��Y��Xۯ[��<�ް��
���@|K��V�C�|�P?�9���<Z<�Ca���S�o6w��r�q����0S2_��;	���q��2�\��"�����Íp6�K�*�^�	~����&��O����.%�����"��N���sJO0�c��m9�'�O��!��&��������B�w�|f顐���/+kk��a?��_@���JE��j8��۞�R2cgz#8N���
C��L�$��:����>���>3�s�Bq�.����9,��/�|��i䁏5nP���/��q���sU��vy�̼��,1_J�:�ЂR�/H�L�;S�"r�]CKH�xOv����xNf-�e���X���]���w>�`�>sp/Mp�>�5�s���N�Vc�ǵI�-�����F�p�L�y���������쭉H��O�M��ܣ�D���&�(�to�#ْR��8	)P��y8:���j3�/�sl';~)x�,�V�74��`��������\ƍtQ�d;�QM}��؎��ś
.$��he��b�*F"�W����/�����Ij�J�tj�ǜս+"I��O�����-�=�`E����������˳ƗNIt�³R�x� ����o-�FN���I�k��%t*�m�H�xؐ�����`�����D)T�:M���ԥ$��L�`8�����s�[K�gv�<���t��ԩ�y���g߯�#0ʱ>���Nl-���j�1��GaU2�g$ҍnL�I�/i���s��Ê0�~�%c�>|>�"\�r���o��0#��M����{j��a~�����{W�J���t�.lhnY��r�̏��F�Ԇ�B1��ܤn	_�[[�ib��Y���u���d�h)�_a�h����B�����+X1`υS�1(J!S�q�5�_9���Xk��#7h$����_�`!~�=�B_�%Y�S2�l媶f6X�k�s-��~�"��p���)��E�>�h����6���	��E��X�����P��p5:��PFi�I�w�p�RJ/G�N����F$x_d��3ށ��2@?	��V�^s���P@0|N�l��WhK��{b�LI�'�Ib�4�3����tJg-��3a�g� �� �l
4ԈꕃI��ZPNo���j��4�1���D��^D�I��[�T���'�#����d����;�c�(�0��8��P��m������K��)r�U�P2�"�%��qL)�WL��y��$���A�9�(Z����eU�<{�a��x�v4,[� ���ġ�4�8�R��������cp<AK�R�!�;=>��DӍ����4� -E�
v�*	�Z`%�d�����F��G4���̂s�y�ĘbS�F�5n�B��^'��L~��$|��x�\�=)5�=�R������O���u�����ˡ+� ��l�U��ݓ�����_�c�^}�}�������I�I_�>`�������Ɏ�>w^�]���cd"�g2�=3~e'o��S�[���_Z��K���VL��4/\�^.�o'�r��qb|�Þ�=k�����wh��~�*�A�T���1��W��թ��>��h�vtk�Z�#G��+ա��O�U��9Vl�9H�KD��)<x\�Ȅ$��;4��ENn�œqz���gTy`���k��B��,��M"��L��\H㞕B0Vϵ(�m���ȴJ�Up̻��9��!ٺ��*�A3g��s�!�!�����MP�c�ξ����e7bq�hR+�7V��I����"��l�}^�9��kc�f�@��%HJ^BV;�k��������	������D�:aW�3_J����Jc�K�8ɡ�7����4>q#,z���T��PhPP8��ƙ_Ԏ	��L2�i�?�V�4�T�4�-y�V�uiTTװ��2�{@�1MLߔ����lk�Md�N�W���y�FrȖ�y��QNI�jc��}fI��O���;�Y#T{{���8��U�>���[�!z�\���I� ��1���݀(��gSYG,9���;���p"ÊV{ ���p��*Tp~��R��{�a
�@��S4�����/�D���ȭ �b���5�aE����G%�Ԝ�=tJ,���|�ek:aj�j�5�ܸ����>�Á�2�Pt��=8��]���E�8���S6 r�"<}���r���H�{O�b��E��]��"���ZR��O���z��ý�nznT_kD!�	�����)�E���h[�tQh�]�ՅK�7a�	�Y
��3�����e�g ,k���G�{P"F��Iܦ�+��KM���ǯYZJ�S��:S�:oM�5�b|#�>ƫy{�ǎF{@_�$	��Z2寙 ���%�x<��X<ݻ�p�i'��l���`s����h�O/O�!AZ��f]#qp>[�Vb�̅*���÷�p��4���3>+q�Ի�0����O#p�~�$��}�ΠL�
=�l��|"����H�h���W��ɔ�.n��VZuy�����l1�&�M9p�e�z��x��@�jO:0���VJ���@qD�/;՛�18bg"��{���D�|PM��k$ײ:�����o�U��ǻ4�1�E��6�D ?�ξ�C׻�C�V�$N�L@�r����`fL;��-�"j�K��mpn�`2�eT����jWI�Ч���Pe�ӊĈp�u��3��ݯ�0ݗ��<���D#���@�z;&�7��&�N�	��
4��b�H�
�~N��CR��^i��gx��4��Z��X�>1ٹ�P�}�P,����{�#KȄ�B��� �[�_:��te#�?O��=@[��l1Ԅ�Cw�(R�{_���6���xJܘ��[c���z��!�5�j�Yr��i~��¶ᐽ���Ȏ�h���E��[�B��0_��Hz�X�`O`-���j���˻D�m�	�T��L#��,��/�l��PȘ��#��!�S�iH
)#�m�u�`C�Vab?�������6�ga��k�V�F!ꎯ����oA�@ݖ -p�G/"]��@/�`��){��O��ϻ�7�1A�C�Tڡ���:|l�ܺha�!CT4>�Q����" �� D�k�����$�13'5����h�i�%���E�T�;ҍcy��?�0S�~X��ÑH�S@�'������Xx2�晫5������B��>:o~u����X�j��]�|��ۇ��%y0漡�5J��;Gq�)�������a�#��(�P��@I���o��s�"�}d%)�|�xh�N��,ig������#A��ɵ���� ߮�U=�dm��s�4��z�Ҕ� ��8e����KMdʣ6E��	�R����:����o�����' .��,�������z��_��`�������@�o�3g�u��ky5 �$����5K�ь�!q��|��h�p������U�z����QT����,o�a��Z�Q��v�Ү���3���u'z��"_r�B�k�p7�)�p8/5�_�/�U>Jh��?�'=��f܂�����%NǱb_�U(n�v�*�j�HK%��5���̬d_��3{�1��kM��U���[�OERq)W�s�K���bV�9ڑ���{U,�.Dծ��DXZ��odb�����H(` ����a�u#�P��r��H�\�䇘G&oդ�eʕx�C{we����*���TRG%�]Z���1mo��nw�m!�	Vl���O��p4����BXJ�6��	'$�0ñ�c�H�#Q�Z�&���f�+���@��p���T���:5�H��귖yMoc���++xؚ�<� 1��B��3�_/9ջ���E֗�gnC�))=�	��^�^S(�b�h��$�ER`iL�v"+r��V=��d��=�*!��)��ȗ���sχ�MçCu�h��������Yn�EtH�e#9QR�Gu�-R�H��8�s�*�,�ئ1q����Na@j��j���v��R��f�����)N����V�^?�nzA*y��
��F�r��g�nY ʹǮ��$6�s���Ov<����5P�g�)$b2M�g'��VZ����$K�VK��adG���v u"b�Wm�oO%�
��M��7W}���:�,5���0Y��_���gP�22׈b���G_�fu���+���|:Yb�A��I)�G셆��j���w��5��m�R3��߇T+t��i���=|�e��{ң�O�s��{����[35S�4�E~k�t�vx�N�.���o��� �qfz�:�m<���i����bN#r�>Y��59�7 �NK�$�)`�����;���E�z�����$�G�<��x�Z���Q���~~�ܜ�6� V�O��������'�mԋ���!����v�_X/tR�,���G�a`����ir�6�8�H[��Y��%p�QkO��Td�n�
����`�rj�@>�|>��H�ܐ ܀9va߸/�;Ov+��O+	����!��)�_'S������!�ʮz<�o?֢TW�v�͊Z�v��=�S���� ﷵSj��]U���x6��!X:�(���XQx��V�f� �E��k��x�����r�uP����F#'gX�j����MV+g��'�ȓh40���J�x�g�x��u�'���
�L���?|����œ|q�Eȳ���]B}����m�|�M�5��-c�Lyy^<B �ИHg������ŋ��ܙV�چ6���o��vm8rV�枢�vIj:4�VEB�P[z�����U������)�ҩ8c㔼�YǺ��!��9�~_�� ���J�3�&'#����#�?&_6�d��h����jl�_N�p|>����3s*��v�����ݒ��[-���<��ۛ)�#J��>��o&��T��R	���p��3�dZ+<�d��i��6���la��C�PjT�r?�`�<V����	7q�k�=�������I���N��;���z	��XC�[2�<��Z�S�?]S��a�}�e6�:�-�}z���lFZK��C߾��d헤P7z�]C�ZR=��,��h���n>N-�����nP��1BN�^��>�`�*r�ina���-��O��˥Z�%��AIJ��k��?v(<���~bT�jc�;���L��|m49m(;�|8����[�.��!��/��q�m��/��m�Y�%$�
�ʎ�`$(<��d���g��%|V2:�*D�RzC�_z��^����q-� �!T�pE���v��Ij���!�x0Q�|�3�FɈd&�Ů�����v��]뭖�<$�?n�z���o�R$�0����/�o�j��ƕu���zO.%�sX��&����Ͼ���D�w*h5E���f���r���>I /0��!%3��~�۴%�2���߀Aɸ�p�W�&�E/�!�$�>�rǵ[ڇ��c�z��p�u� t�K�Ѣzv�"$��;+��T`2+��H�������
y��0������}�e���4݀s	��F�e���)�׬3�����L/2���Y�>MA�"�S%��!��K8��;6jI�
�%QY�y�{�͙�L4D2s!~6b4%f1��y6:�0��.E9�/6��T�J��P��)�ri�JHN!��]��P]Wf6n#K�D��!!��7L�>H	�V@�K��_2D�<���Ŵ���%Xt
�^^���O��vT��0��D�Ń�^�uTB��B���hx�/?�ˉ�F���r���A�F�I��[K0���S��{T��R�ӡAc՘���������e�$ZOqY���un[�	Oަݙ�@W.���?��O�`p��%�_6 �:�(�6#�L�K�&ec��F�����ǁd��ў9�2�*R�ݾq���|=cE��8c"S?�[agf��
_�N,)��h�q��>�V���fz��7�4�I\5��mg�NU��_������sl��d���dTH�t�{�χw&�aoS�8V�H���@'���u- ��8_i��Ε���s-Oq2O����� -}!���Z8��Z.���(��aZ^c�V����t�/�~W���21¨��f�1,�p�v�Bnk��G��M�t�X �E� -���d��ȼ�4z�+OWq��k�f^���"6!�RM�NO��_W{�˟v�d<�e��k&t|��d��)�,��##��VA0>'<�4�;��|hÿt��T]mV&�>�}��>���g}"}� �8:u<��|��.$ݠ`���xJ��v���,ѳ��_���3�����x�����Qa�R����j@�l�F!'�?��[$�R��e���F�JgV��HQ!��*ƿ<9w�n�	�M���3���N��������%��z�:�9L�r�8���^�֤|Q��ڮ�P��Q�آ��@b��r�R��1���ȸ��O	�P\���*+�l�c�vXQ���h��yV
<�W�W�ê4�?��FQ|C!m��Y���	�����(��4��k�>_m�h7+�FQ�⨱�$B�ڵX�nރ{�U&�P� If��x�.v�����~�p�aB�'�?>1Z���u ���]�I�Z��!�J���E^,Ņ�`�-y	Xr#�I��]w�$�&'��������~_l��7�1�j��Q�~�)|Fc�-�+UyT���}rT��_�m�&ޮ�a"�00���Jԝ���%��'�R*�~� ���ӦZLMиqB�_k;Ĺ�c�r�:	�������m�/h����v��-+��_��yk�|�&z���~��T�@� ��'Ř}Io�����;�� ���G�`�,/Xs.bˠO�n�����:�W�Z�[��oc���YfAldhC&��W#�C���U֯a�Ƴ���*A�v��HM8L�/���U\\6B͎��Z^LQ1sf��!	sM1�}ʟ�@g6�y�	Ӕ��A��2������3��7q�/_H��CZ'+AW�Ǧ�raA�N����(0{N��ٴ�����++�Y[��`��e\r��b����XO��a>�_�'���Ϟ�Nt�!��$�c2Lv���,�+ .f�B�1;�n�+?�����k�$�� 尉�D����$%����w�а�%�yK��ӰXj\�=&l�U1^���6�˂5���H�b'/����W
0��,�O����?�+��T�M��sh��f�@�N���œ/\�h#�&iZ-j�.��5�Z�S�2I�����Z�,�S;@�c���Ψw=���:��:��2b�k�RE�)+Ƅ�pb�SV��K�8M��2��3����(9�~U�d��)ۢ&XSyA%����4��?���x�7��AL��"h�O�m@�~�{�mb���֤r5����A�oN��0K!T#�Ne\;�b E`�����L#c�k�����	?B��i~��#���"���Y�0܁�	wp�!�wac�R�d%d0U5��xr�yőd\� Q3z�t<6�m��(a	g�jqG*R� ������?�.�i<�P�c���MM�z�?�A���Ϊ�L��q�||X�a�p�Wĩ��}�n4Ɇ�=��bJ^�gK�:�)T�6���s�߂d3F�<u�	�,T�~-4s�y^.^�e�a�;�Y�o����r����V�	7����ޫ����;6����R��2� ���{�ЮC����5�K��r�#�[�M���Ex�	}'@���UC�n���F�IWA�kT��KR^��56�Kci7_L	;`2���`A?�Z�wS��9yQ�X)�En�� ��o<��/�ź�L9�i^j�g�4{%�a{{ �$$,�����X:��C%�'������橊��e�	���\ZUԭo�2����\+�:6�c�E����i*��\�v�S&L�d�9�;L�r(���i� c�G�$�K�{"iQ�F,�ܯ���YU�*M��+�o�b�Y@B�u�3B�<�(�	:>��S�4�QE��(��Jy� �C(7�Ka�:�翥�ٲ����]�<�Eְy������1��ٿ{|�e�;�@��X;'�"L9���[��l���4!\���)�"a��[3e���%�1� O8Â"
��llfД+7�Oj���Mq`�|���d��ND����ɖ�p����?23@0�J������p��7%��I��pa^���؏�������::�n\W�^.)��$��`��Z~(E4��@���y4����<pL-1<�K�Ǣ��J���g�mՁքMMn�]����)��DH��v�JB�.��Jv��V�pKO�5��?������p���뱗`XTj�`�����?a����z�W��ΐnc0K�R��C�w�5>��K��n��u��X�c$TS�=��0���,?F�+a�<����'\/Д�؏����i�j-"���q��3r���l[�GS�m�B�m80~�0;
�b[�9Qv�����d����ElIZ)����!��*P�o�K��V$[k){0��@t1�
��K���Q`�]l�jzd���E��f-dXM=��}����U~:�/��*=w��%��3H��.P�p1�W]���ּ��L8�[�����c�4���Fp�T)o�O**e���� vt�Y���)��N�j�Ѡ�LS�(��5ڷ���ppH�R]�4�����UK���ك�ͳof��umk� ��@E����f(- &�ټ�e�D���J��	�xx��c�JT�j��&G
\qz���*��=��.�Y�=�1��Ǉ�Ƶ��7�*|8�΁E�>�#�o�b@���^�����1��y}E�.�C�zWi)
��-���Z�@���x�%�̈0R�J�+�|
�e�Q��|bo���>�?�����Q/�̚GQH�����Y~�C�A7z֪~�A��K��ƅ��dY)0�=�E�M=�T'�;	9��|?l�ވHrך�y��}��i��5�ш`S���T��ޮ�_�'�p���%bfa��hPJp:��a1%�u�įO҇A���o,�uq��ji�3N��'1n�C���E��F�<N[FV�(%D�w9���I�Up�C)��(���W3�W��E?iP��R��4�d�q]��3+`r�`ޮE����쓊ֱiA��a�j6}2�ۜs#�?|r8�N&$���up�<��Aأ����(�Ҍ\�Z^j Ar��ĝ��bT�2H~!v��<�FiMu�%8T��Y/����X����'�$��1%���a%�����ԅ�9x��~|
��#֘���O��?�V";T?8���	5��q�s��nV|���,�i?�ψ���J*Oy�I����S��4�ۺ���o���atQiQ�Om�7k���-F��<A� �Q�+H1ځ �9��EC�qܕ�j ��
���v5Y,P2;�?G�����AZz��}EBX9 a
W����ٲ�Z^�k����KC5_��UF���3>�M��������:D&7H���8f��(�]W�Iھ���@��fxM��G�����������R��q�t/una ׺ 3���U�Ԅ����
���&�h%QB0�zn�ى��s�k-f�{��gӁpp��$��������tV�[����!��pzD�\$7dJ�Ƹ��N�!��g5oM�ӈ�Te�#G��;o��	���H�@a�S<qp5�� 0Ne��64��R2_�|���I�\o�a`P���&ݤ�˃W3r���X���Ȇ�!��jj��P���ٓ��j��9t��j�9�B��6<����y�hHߤª�'���Ҕ���r^EӃ`ɼ? �B �@M�u�����7�����,��ޙ�4�8;b݈s��d.³��ø��y!W��8�+�R�2�Г2�+d+�ұ� ��_#�V+�6p�����/���ĳ��8V��3��y5瀼�4{�2���+xYeʿr!��p=�l�?��1�U�Њ�sj�l$��&~��%������7�x���#�,<kW�T��5E����J%�8�c��N�ea�R�����_�����gs��)�%^G������|k�`�)�,�0N�I)����R^�m��oV�,�ػ#ڽ�l�qqD(�"�\�Q�o��q���l��V�<�;v?<�Hw���b�y#�.#7) �������.�lJQl��fұ��$��j�\A?)r��e�����'PV�(s9f��FYM~�|l��hX^����0��;���7�l(:�����kZ��B,У�)�J��C�)�3^\���2��;�r;�麓�bIC��p���:g�Sgs��>8�"�sS�^�#O�V*{�0��5�=߱zxy�-�W��e�T؎����'����?a��0�O2�dɅ�c��:���h����^�2D~��:/��)L��6]x{LN��[iU
.�'u�T�\�9���(�:��D ��s7M����A}�`�!5�&葻D�jg^�p��%Eoh?����tC����BqA����/C��T�m�@ݻ�+W �M����3�/П`���L\b�v�\]͜�i���ͷ_����� 5M�:D�{�5��ٷ�5�~��g��N�/Av#�H���u�ݛ׷�	v}2����*Un��X�=�
�CY
1�\g+�&��AynB�T��~l�4:�����o N���5� ������ ۶�$��}_cr������ebʼ�׌~� \�q���w��/�!�>�- �n#T5�f�Xo.���<@�H�>��ڱ܅�#f���Z	��M�wcsN�v�`ހ~�{A�+�j�[W����@��/G�����ͷ��|��c+���0�Uz/������M��@`��>�p����6U�����	��UG͜7l�DtU*8�&�
���M����.�:�!	�$���^i�f�P1��ŠG]�h�"��"EK *&�W�˛EfB�?xT�r��7�������ۤ'���G\�Gq��ҏ�[JP��}5�{ޱ��3��
'@z��t�{=��59xa��-��p��7[�~�/ע������Z�����c�Z$��C��r����7/�.�.c�C}?�Ѝ6�o�HGGB �++���W��Z2�L�5/�/.#���Yn̎���xL&H�Ȣ�r��&��g)d�n&Y ��9���aiT�M6˭O^q!��ѕAרө=�`z	Q����_ Y?^��w1�6��V��}�?��8���v[-P�jI��9�䷧�^�J��jdp4!q�%�b_'$�k��m&�b��m�in��՛�̳�_�e���K�t�
<�$�� [�U��~<d]���<�odՎ�����P�j�P��h�lA	]yʳ�L��-�u�+�~~L++?I��Z ,��M|^k�:u@�x����*�" �ʹ�F�{=9�x��ۑ
N�P�iص�G���M����.�=2	>2+쪕l{T��Ga�d�����p��I�7��N�y
�Mh��&j9�U��O���+�+�$�~��֭j)M�sJ��R����	n�p�g�����s\�\�{�_���_h��Aϟ#X��B���Y�%^O�#�f*�����T36y�A�X�S���o������+�>x�|8�ڣ���b(J�a~�e�Q����̺�l߀�Oj�Ѷe�@M�e�����B��ƌz�]���Yw����S�"5V �y�X�-�?5�������, �;)�<A�i�T����G���̪V�9Us�N<o�����k.:p���^2-�AD�x�Vh ��
B��G4��������5����x�����T�6"��6̴j�Ny=��1����I��z��I��E4�%�4K���j�+�9���I���LtO��ܙ���9��M���H/����?�Ƒ���!��u����s���b�e� 6�a��vh�B��� � Lf��r�;5�K���ĕ3���F�#�����7�Bۋ�L�LF[y����Q
)�01�d!�#�f��F{��/��4G��}�c�XǲB�Hf���'x�2I��<���5����d򡼲"�f�p}�X���)B�%��(u}��ϱ���}�	�����o_ŀo�1���4XTHD�&>s�B�1.�;�E���G#�e�x!?!J���ۭ*�Nqk����Ũ�L�>]�L�0��&b<���u�
��w�C'ع,`�	[���Q@
L%"��tCZc�[`w������O��oi�:�ɖS�h�e�x��	�g������xĵs�"�� ū#���X���$q�0aM���+�'��d�(%<�[N�@(2��8Gt-� +l�Ž`K����uex�BQ��dT�if��9��l�<��}q��p������ـ����.q��ZW���
��� �Jwн@ȣ~�e��ŽA����z��p[�gzğ>Ɔ���sj�ż���[���jY��]����n�9[& �	�0�"�v�b̜M߄�mU���t���_M�ᛆ���Ìz�7a�5�E>�S�#Yu�L�֦��{�Fi��[HM,t���l}�5���<��D�$�M��d+R���2/&��T�%�]PLr�&=�� L=D3k��YQC��z��Ծ\s&��|(��Z���޳K�Ӧ���z�
CC8�$ �Y.{d\Y��u��i&W�M�� z"��!܎�ɳK��������,D^\�#	�ͥČu\�L��5.�������0:R̯��R��(�5�	�Cr����e+�x������H�)�a�[َ�Y#�y�ABzM��.Hǧ����	UV�$���zB�W���*/�J��0;î(2����x����*|��hȡ�7y.N�;C�]Ǹ=�B���a��R����Llf�P����G���%�i�
�8�Q���ڑN��%��	�uա5�e�hΗ2������0 F�؉�X�B�c�7���8��"LS���C`��m��*��Jcb�J �����;�$F����lH��%�IM[�C�:��N���?��;��c����L�2`�" |�ŭ����/;|.��;��=����<�O;�S���O�"��-�i���j�1 0��Iә�o���CȻt?�?	��:��w�Rp�8Gt��tx-N*��Փ"4S,���}*&C�&�XfK�*���G0��9��)LG��\=%�
%�+|v�AZɘ��V���l���[8���w�h� `�3QL�y�]��2n|�����#Z
s��r��3�0�v>1��("�W�B�4ts���?�楽�gk�jfu���]�Di����B%dۚ�K�-쀱p�eˢ������'�o-f���d���FL���U�8�b�d���zڦNlI ᄙ�L�!��/�D����+d6e'��}8��J3�h7>��:�7 G�k��O���Ѓ_��@G���-�h��F�����-����~It�V�p��%�z̆����˿Չ����ʟ���,��(��̚0%��:ۄXq��l-U<���*�����2��]�%��r�#�W]�h�6V�h� 1�OQ���Mk��TQڥ�q�8YB��兯N��<$���18����/�hP�6�oO�8 �I'��eY���Le|�S�j/�C=�0�8���V�J�|B���tE^}#j�:���--�թ�6b���~fꄁ�ӷʻ�b����q�Oc	*=l1���z�e��$�ڹ�E�<-Vn���Z'���b�G;S���s�5���ϠٌT.tp�!rP�ArD`��3+{s3��=(�M�T%	L⣻ؤ�H�1�4���p�t��_����k���V��:�u_8iGnڴNkOS7���s��$)0T�Z�G+���g�s�>�E.1|E��C�^]�K0Cu{������u���8.?TU �S�C��k�ƥ],����6�'��v.{W�Υ��aǏ";uf8C�` Oa�P%"� �iC�7N'�1)5H(�AyP0�ˋ�.Ӗ��SRX&��x��uC0n�e�� LZ���]9�"ὧa��q�OB�w��dɷ�<ǽ�l">XDMgx����c��*����&bJ��(��Q��߫���ݪ����޽R�#��{w
Oj������m" t��Q�fI��$5ve�Û0{F���6��D\mYޫ�l͸U���fe�c��+J"qR�^as�;�VJ���l"tR���Ek�;������1��J-�l��>��vH}�#��f&R��L��K�눇�d�%���`g�Yq�[��د!�N�g�2��)Z��-��7�hLq�e��{0�a����.6:����T������+��:^�;]o�>�]vB�q�.�A�Z
�Yg>�Zv俬~�����U#٪x(@R�Q��Us��-%ybQ��~�WYt����>�"�p�ڢ"��vn�-b$v	�`�Yg��ٓQ�
ތ-2���-xn�H/�*�۳����!	IY-�^���Q��D�qp"��)�W*h�9�6�u����|gOk�l'��6|h�>���N��	7��I}�hn��+Q7Z��()�qxn�#��nW���\إ���"�ХF$B�BVe�^U�4:�&x�BB����1~u�۠�j��Û;�9�zrLt���z�c߁]5IV�d�?����'wLGY�.S����\�,`��� �і'IX�����S:N�&�И�p��ij�Y�ouM�K�{ ��I
�/�z���8�C�4̄�N�� e,L�����σ��X���(�)ő�(��?j�y�n� hcL�ԷK/��� {B�0���oD�h��<'�W T��w�_�S#�����&������p�Th4�Y��U���gy�']k�0�A���4�����Zr^m��N쎝;���ҧdNڙ�������:$���x��x�}�}� ���'��J��M,���
X��o�e�+'$@�yVqt���4u��)��5�扜��-(3Y����/��_� ݱ;=)�Jc�͗�T� ��*��7�q��l���<\?h{[�D�;�bqݛ��S��]>��W�S����{��(Y(͋p񪔡:&�I]/�P�5�u�CӰi;II�]���}H�;�#Wݗ��i�����G�Z��l��eى%c$eG`�#	~*����VԊMa�
�&[hW�'x4/� �J"��ئ�N����i��Ho��܁�Q�$���s�Y��	Y�+7'e��*�����@jK��O9�;��-�]|�"i�Ǫ�����⾠��f�� FHߊIǟ�R��vS%�'��yDN%�����܈�����DkCbz� ��4��MhŻ`�g7LW���;1�%�����w,p����܄�cw������iM���w��ATi��q�y�FXG�|��%9��~�������\�~ch�Ǐ��){:dN�ez������A�td���N�a�h:��C	%����iH)�A�7�K��|�=��=��Po/N�@|�ꇄ�ʰ�~��K��ll����BFj1�kI3�.��m[�,w�����@Jo'���^ζ�!��ɻ1��Z�H�P��b����:v��ՏX�X�~[>��+�/�Cx9�q$��w<��b�L����/_m����Qx������A{�Gg�l��K�Ȗ��~@��Z��O��Ծ��uГ���\�2v��BP1��<Pݟ*�ĺG�֊�qX�]t����i~�؍�+��r����iwJ�٨�$�2ٓ0�~�*@l�fP������D
];2_U�����[bIh1���|�3��T�Ol�(�:Y�Nhy�Z�!�T��s/
I�/�G0ձ�����ZK��I�FNv$!d��1C,ҥџ��0�#�����S� �C	�n�/`�4'yʖ��a0$�9���.�ك�~��F��\���C�����-%W�T��E�I>��0���.%S�a����EKx��Ό1zX9���uK5VO������S8y���|AT5�vF�_���/���0ɚ5P���&@��hƅlB�T#a�����~��לR&�㈁�R0�Ǖ��l��1\��g�+�d�?�gj3�m%0��ƃjx�T�+_����G!��/��t�G�ZAu��B_��\�Yw�!�y"�ٗzTA��C_;�e���k�<�]� ������S� �X�>ϝ'SMN��U�a�77?G������N<K�����`�`V�ש@`)�g�+���寱_<t��k�t+��LZ5��s<�а���da��娛���b����j�o��π�����|��^�Apwq��ϯ>Y��s�@͂�\�H�u_ �d��.O
K�]C�^����CIQ�@Yp1\�h4�&w]��>�J�ק��V��I������ /����O��pqN�Y���>�pE���Ԭ�p?�Bm��Ȧ���B͢�k%Åz���AzX���T�E�h�<C]�9A�a6I�C=�.XbƜ��5 m �� ;����Р��*3�������Q�~�_��+�qŁx[5LI%�y~0]�}�Pۦԣk��q~6$>\�E�x��Z�ݫ0nܼ8u�b�Ma���Y���IW� �:���=ܭ1A�tihI�b�+����ӯ64��X���
D��f%%���^6h�峨���s-��c�B&pZG&RE��tw� ]�i	��Z[���f�@�I�PP�/�m�!�!�8�N�=T�n��>��C��=����9�0gs�q�g�N:p�� G�>_n����%b*���D!q�BN�
nx�����.��.۵6B�ߙGP���
#r��*�����d(�0;o2�+�#�r��G"1TT���,5-K����rl�nY��j4 F�M�:���E#��PjeJ�u���{��V]7+K#$	 �$K��c^J|��P��%@o��C>Y�;%býB��M�m�����ê�So��k��'���D@��p
��	?����8ꈮn@<�ޫpaj_��Ra8�ŬTNs)��D_ �x?jF!�jg jE�SU`�j�P&id�'�[�{�D�<�葪'a��9	��ڬ@�V&C�>=���G�1� {��K�K窳�,@�bޠw$��a�"�P�[�g�/,�c���G��q��0*�/�����b
KyC 䘼���p�E2�V�b�c���5��q��_Y�%KM��*kLm�S���}�D��*�O�|}�:%����,�gL�Q+t�F�E��g�!����`�x[	<Q�SF�����t1�xw�M<2muO]
�G�:M�=g+��7Jے����($@`�����������`��a*���X��4!��҅�R�Z��t�/)�jy[zV8Å�q���퉳*~��)���rs0OK�Ҡ ;�*�02�?q-��ak%��ng;V%d�@sr,��J��!9BEU�6&��(EdPeE�^/|Ԩ�*K���,�g[�����$�Ч����B+m�.L��4} �e�8gH�1�YK�Ula�������%�ֶ�1��ǌz ě(A=�t� -+5{6�g�7q_b�"�#�IAG4~��ZxA�	����O7 :<�7l6L�ɫ�T����h��zU�A�s��T(�P����mه��bQM�$m�������:u����E1$���B���<4�SG��x�q��_�(�'F�O�I���)�6�c�7x�^z�
�m�J�X�n�y�;N��2��M8`?�(ş���\�P�b���㤅�,Sv���?+۽(���zr������^*f���JMo��)F٦�t�z�+ϡ{���1�<�H�h�S���S�����1Ĕ��Q9��YWA��iM��K�#�0;�|�yO���c��<�@����;ۯa�֚D���,��hMI����"NZ7��˻yޟ[\����o0q'��Ŝ�,���茱~��2où�W��JB#�����ظ�u������k��u��� �||��N�I� #-Qz�l�}�n�?���J�~0���p�F�=a���&�kp�����sGZ?(�0�,Ɔg���C> *��S~◯ߣ�ƪE�^߲���O�.P��#g~��H#�G(;�JtN�C%�>�!�2����@5�#%6}�{�Q��*�b�k���Osn#�=1(��Bh�Z��T� �(Y�ݑ���{��;�\.��
> ~�(ۻME��{C������P��Mq���i"B��[*!���ߍ������>�����ZA=��	�^ȶ���Ǥ�nx����~�
�$Rp�X���XBi�d;n����ArQ�h]+��34�~���ه��HU�j�������g�؄j���b�OT��"��B�X{�����m
iY�.�A�f-�f��u�( P꛳��
z��\oѾ��37��R���A�9Y@j��z!F�ƶ �����D�,+�Ќ��+��ſ��\$�T���~x�3r3ς�.��͚�p��I�V�үBUH+GY`���0%�v�]yc����<Zu#Oy�����L��-	�G�=��ަ��j�����
�Ƽ�b�����H�1����� �lǔ�dg�^�텊0K�K`��nv#ʭ7�1�(B�g*����U$)�Z_���c׭�ו8�7&׈P�'(�xGL����-v����@L_%�l���n���/��fQ����B.�>�z\��	�N�Yϳ�6L ���o�}�&�q��bǾ�O�Gj%��Dd����Oe@�cv]�J!�����qww�mGG �I��u{�2�ƈ�89Hf\�K��4a�jaV�(H'�+�����&�Փ�v��
�&\�'�+4GNeEb�*
$}��쬾D���Y)�ͫLKjY�E��hW�E��_�%�����;'�o �FO$�sȲ�GK?�9}}lDC4wƪ# ���"��W{� +f���m^| #��G��;��3r����i������b���:yM�D"m��6!ΗT�&��i:1��o�?J�,1�Hr>(@[�?��pV�S/ٿl�vPXY�~kT����dv�o�8֧s��RJ�(��!(��k�~�ǃ����%��P��z�|�Ycf�o��s͔iET���8���L8ٙy�7���%ڇ��f��A?�����u/�*�)ZŚ���g��[L��8z"LB4]�������+�GE���&�e�ϔ��)�J�����������Π�!i�l]�!�� {�epU�f����� ��
���H�۔y�-�;��Q5��~��~������wad�I"b���0e�*�~Q��q�y�"x!�Ӌ%d��2Y��k��8+L��5��+�|�;�"����;�t�����G�K�Ar�5�a��&g���m�+w5�G恺�3���}۽�����Ɔ���נH�Z��4 W��Y���Xl��������eT�PQ>�uԛ�ā@5[�^�����EM^qp��cV�H�D���.�����u&K'[� q�ߢ�rdi	:R��£��\J�X4 ���;���&WW�ؿ��\���xk��(����B��&c����f�2���\�x,���f���m�9�O����z!��S�N\���
�/`n�Y>=��t�!��	o���l�Z�P����a���(O~���O��G)�^S�=�` ���)xHjG���Ѧ� ��U�X>��ozP�iN��u��/�c��)�|�iXw�[Q���Jэ������r$�S2��>��<��<��OU,ն��U�I%[Me�A�Á!Ē��
h���12x&@���t�!n��
Ԧ����o���.�.(P|��r���坂��1x���y�6��?�;��R����u����~~���ṕIFrBF�9LZ��%P����j��ӯie�hJYΝ�2mڒ$���9�bH'X	�"QȺj�3�l�PH��?w�0w�G��x@n��0�j�Q]0F�Aܯ���]d���Ɣ�s�R앩�}��'3<��89!@Tv��ֈ���r�oc_p!,
��۔����ER�Z������V����l��̃�	X:�v��V*���#����>��iܨ���е'T���*B�ٖ�� �[�~�3�*���Le�뼾�v��2���y\
Cu��3Q���,�W�x�S{�f�{��<V/�`�j��ԥTg�2���
]+��S�9�sſԿ`3%����L�IصM	Y�7����ZTY�4TΠ%/�U�e{"N�����M�f�d�_��^�3F1�[�t��y�{��o(�8ڌ8�-;�Tf� ,�AOL�$�f���E��R�*@B\!�}��x%�bΥ��A�rr�5���<���.�р�_��V������5����`u%+�&���}Cw����$���C����S*����&[wV�����W�k�<a��˘AN�2sF�+g�`�@��R��?"�ZIv���Lg�􆇃"塡����\�[�_SfQ��m������xOߟR��NK�L˂�:X��2�C���T]>5"!��V0:�*&�|�=ڴ����Y��t�ڳ� U�4��a���څ��!	��.�n��d��g֣�q�"W�ՅdÞfFݵ{��5��	�È��U�T�/M\ }Z;�Q�S?�����*O�O{
ʰ].ކ6{�$�^�t߉n�֝�0�%9PPlzW
D���N�0a��Bl�ecc��S�~>��~	�R�&^Ւn9'>b��#zE��m��"yw7�?Ѽ�  �^|�J�c.��U,#v�_o�D1����3��H�:��*o�tQ�1Ln�1�"�ZQyY
���Cu@�^�#��˖��֯8�u?�f<b�
��Y�v�ۆZG}z��ޟ`��F!�����ZM��~W;>	��N�1y�<K��I�.��r���KW�흫��K���!]Uj�=��cЉɔ��XO�9/�k��(��ݰ��~�WW�4fM �O��t:5M�.��5�I,�0��_O�mL��N�׶����jiG��X�+g� [�OXO��Q�caV�Xu�̘�Q
��)�����T��������x�#q���ԥ�g������s%A}�`f�D˧����׿����O(񚑙'$c��N��A�B��J+,�$X���	���D�ex����N��}j�*�?0n�ںK}�z�4^��u�B�w�?��Z!�T�y�ɉ�NOs�/�x�p��n��b3u� G	������NG�ds�-J�N�d��p��3��<'S�i���{M\�ýƞI{>��h��܊zf� ��xg��t�豀�R!�!�b�:��r��bˬ�i�V�Y�-�m
���>��if���)�mfyG k�Y��.���6jg�EGTp�˿�aX��^"OvN�����ȽAԡ���oCv3����y��4���y^P�>%"���$[϶���F+r�S�bL�.� �;q�R�T3�O��Hg��.+#"����s�������� �)��J4�ho�<j�gVOUx���u�Pc�L������������O['���e��^)�<<��M�Sh�|��nĂ�-X���^3�3f]^�CY��0Wu��|�qฯW�Ģ(��u&{ I�3x&��Q6OY�3_!'[�ě�B��fÈ���I���cm.��3�[�$1!'Ơq�O�B��fe���x�d�M~n������n9���w!B�7�Z��/6^S`��Ibj�)Θ(+C ��+�cQ�c�Q5�1�u���o�Sqͬ�b=􄳼����e�$Q�k�&���d����Eп�P���5nO����C�Y�j�� �`]�K
���V�u!�i�;h���XM0,���M��M� T=^�cd)h�ڥN]Wd�kBR��m����f@������x�3�>��O��X09\���i�B��n%(D��he��'~a	0O+��5AT�.4�e�wunU�F^)z�G(m~ �̈́�O�\�z.!���i�5>g���q�Q��I����V�!�^����%�n�.�J

{�N.(�u5a�0۹��B�MB��=MYL��P��\S��$�ŰL��3�	��u��m(���LWE�X>���f��J?��W�f�`w�'�U��{��jh����[v_#�
�ɛڀ�}�r	���q��6R�7/m�?=d�C�u(kJf�cN�q��!�	�����	���tRˤVwh�Rx�e�N3�2�8v����*�J�b=��%�,�N�_QCߙ����_T�J1u��z��xO�-�-�QN�5�r��6�x��դ����yAP2��{h�Zx	s^b���8:S�%���  <�WN�_�B����U۠M��Hם��~Z���;?�0� f�k�g�+�~C'��QH���r�#|�*������rH���s��[�����"mڞms�y���,u��zϻP2&-9_��o��d��R	+�h`8�?nc[�"�u7&��;~����s��\��&�Gt�ԇ}���"����aXVN���D�⠫����!5�/�9)�ރl����'�&�z-v���ޑ��'*��H�F�Y,|�-͑݁���G���"i�yh�E����j�M�K9��c���w0�Tx�,8z�=��]�6�ܢ���wg'�Y�B `�oh�$=�L��3�P2�n,�wcM�g�i����l�����2+����v�1�O*za�uA����y�[M@�'�N�]���-pc���n�R��R�*��$�wIw�dq/5du��=W߃�����Ȝk{/��Sj�$��3������O�]���ɾ��H����u�.��O�Ж���p��������f�;iXI} t�N�:��&�gL����%���l�u��İ%q
C���FTQd���� D����my��ˆ�����	�3a�������Ҏ�~�6��i9��8lH,?��M4�b��
SS�\|��� �#��h2ĨGL�6�L������0�Ç�3�>���� ��������c�K"��p�<�N��t�8%�-eÀ��٤>]!;���Y��?��?t�8����VR8q�������N��ټOX�Z�]�ꚸ���bV"�j㽝z!�S^�IZ��$�y����ܙS�+�y�G�]p���
��K��4v�&=/8��O1X<͕I�0:̞Ř&0{�����O��x���S]��B�Q�k���O|�Q���H0 f� |�TKtbi��;�yd��$VA�03$������:�|%*ߡ��ok[^T_2�h_�.�6<����Y��v�&Q6��M���vػ���z8�LF�1���VP���[��͟�Ml�1�o%�s�
�"+F��&���0���Rb�N�̼\��.� �BA\��#�*��Հ�	�����\�;���Exs�{Ln����Ka})�3VԂz7���׆v�5��a��:�]�ԓ�1n����&e;�qw8����N���0''T����t�/V��GC��ODC��(����]4�W��zi�VI����%�cm:�׮��?x�}	M�>A�rxCA�'���Qu�����W^�y�X���BT&��d��Sdy����}]G_���&{��LXxG�r��Y�h<!ڄ�B�UZd�r�S�b�4|Y��֕ѓMz�&�3�jV��Ƭ^U�2IS�mG�
���{�ef��u�h��N�im�	
�LJזo��J�)<�ѓn[,57:��� �ވ"�̠22�U#��</�1rG�Gx�E3W�tISe#��%M&�����tJ�܇�z����|8[����т�bP��|N����H�H�Y���;)�S��Y�	0)\w!(��,W^Lf1�����������%哖�[�wh����*�w�R�q&+I��}\Dr1&�? 	 4��FB�NE�һ��1(��5i�	�����%VM�5�$���p��S.-=�߬�A㦐5�,F�b�� Q�ЪWݎw��7ˎ�q4��aB�t��5`2�l���:��&�)�p�T;��g w�mY]�gԊ�m�8��.x��wt�8�n
��F�Cla�iW�J��
�-Ui�Y7�Y@����t�~���j2��p�[���w&d��i��>��=�Zu:!��q�=���+KQv(�㤃�8�1O�	0L��->�om̟����������c��M�)��ֲ�n
6��+��
@�QOsʦ����b�I���@���ag�[��i��-b��:�	E�S�Y�KKs�ʏ�oዧ/f&�aw1��� G6���J�L�6�❤�o�L.��l��G�x�z<j���J�a$K�=��Ye!�>S%~��%�7m�xCJ$Kb�FX�j0��'���h���C6 ��/s���l��9�c�	������n=�w��	�r1�;�B����6���a5ٶY��N��,:��W�IS˒�-��a��~�W(�8Y�Y�E!{V��@�5�́�c���%kk~���d�1���p��p����6L)�x��RRBݘ���i�(|1:v�4o���HUF+�� �~��*�f[xmoU�����01�Cy�~�	er��N)�����}�]��<zbJ�rv�u���a�3��\������emµ$��P#t!�U �k7N��M���v�Zr&��"�7p�
����:�z��	�P;��\.nu{���Jm�|�|�s(�A���sn�8���l5M�+T��Y7�l�Q�t�i���� ��{�������{�<B��ck^(w��4��/�]�z�e�w@�Y�Wcۑ�J����9=T�{_�eõ.��
�(o���	|�P��d��Wl4}��(ATɆ6vp�<���-��O�
�g�'4�S�q�ه��\�.L/�Vδ2�-WQYG�!��I���S��*,~&�%�v}ة�t���B�Ok ��/G8��)�%���\I��p��8��FWRvW
��8����|(��-CdlwYK�;-�n����ΤBp~��-պߡ�-��M��,�,@��I��CCF����)��7�6��D�C%L���ŧBUx��Z*�rn��ݜ��V��3���8�N��c&m<1�O�k�hM���ԝ�i�b3~�N�y򟟔����P��/J?~%�~�v/��k��q!C�7}�$/�:�/�4ݥ`p��6-T���t3�8Yش/�z)�� 2�>�
~�q駅~^A�s	�W~59 �8^��9ꆦ���-1ywh�ɟ�:���uqa���ɚ5puٙ{�Df
ľ��t]�����HE��7���b�_=����?�&h�	�&���2�1�\���sIȳ�=�u��r@����ƶ����z�(iOp�e�z^���0CI��U9����<V{ǰ���{Ն�.yQ��Vq��L0va��]D<�`>ڭ��x��)�{\��%��t�W��L����5r�kƫ�7�ʯ M�0"bn�ؽ����:/JM����U3�����_����Ԟ֣�`7�2���T�������J@����#�����:D�tp���lb�^�Wi�H�H%L�5���`���U�����z�jհ0�ZVtS�|e|�g�y0y�X�C�i�P3� ��۝�m�A���	��]�_-|Ͱ.����
��s�]o|�
�Pw*徭�R�1�NW�(�۸&����	dN�kJ@c���Z2���˧_`{e���7���Kq,Es���gKs�J�;uHАs���(?����u�6�bIL%M�Q�h[�V�.��)�/oJ�B�#q���X�P�:'���>�snT����3�0�`tUq.�B�y�!ם�,�kE~kX %���&�L���cA����}�=�Cb�[f�bh��k�<i���"c�־6�6�M������B�,�����np��[���浿��'&����c?�Br��7 ��������F3�>�j�9�8�g��0R���
\wxbR2�|����b��j��ץ�5�5T�/9]��G&�C�����DB��ȳzd4��%w&��i雎1$�Q�,����>�������-��	v���GMke�x�eh4���[ZbS>�
��4d^)�=�%�p�
L1�g����>��?�������L�4^M�C�U�Q�E�Kd�	�p�3n��UQ���iY��3�]�2��!A�=�)o�tJmt���_��
���³���z��EO��6�lp�� �t�0o����BCUl>������Wݡt*��;�ʀ��Z�L|`bp��_<w�(r�x�k�&��֦^�?km-Wuy�RD�:4;���!УII�H6����S�|k5=���l�ȋ?0�PAl�?�֠+�Ib�uc�E���8��0�2��gev�`'\CT�������S��GM��"0[֟ں�3�o����[���1�j�ބj�6��GT�x��fGn��lr"���F�?|�f�B5�0=�.B�6.�S���?ϖ�N���"�_|+�o�u��b��2M���u����=�lh��L��䗇@��3�w�c�<�F]k��$��X��9�S2���cweC�7pX�iÚ��_	C�hW�����͊�í����9�����[�R�,V�ϯ�kT�L��a@�Ԟ�Fte6t��A-�D�Eh�U.܄�>����Ej�Xr�M)���C��r�!'R�m��ˢ�0���fkœ[D�v&$6q���ث��C� M�� >���چ"���e�·+��<o���n�(G�����W�<���/���hd��v����5Z�'C�ex��	�"�������r�"F�xۯ��:Ă���x{ٙ8�y�{��9B�Lu���������n<6�i�"�j����Y}<_�ۋo���2ר��cX���|z2�<�`���W��(b���yGi�*dV(�փK��f��a����v��89A�3 1F^����Z�~q��Yk�ڐ�G_�'��P�8����s����+�^�����W�EE��~�N���!� ��]&���[� �b1Ia�#S�����J��r�
�XM`�_�o�~��4�p���� (����[��~�=_�d�h���{�����!�X�A=��7��5LV��� 12G����!�[�Ef��Q��"(rf�'�}���U�)�B�����T"A��_ă������a�����K�U}��2�x)@�߯{�$u����Vl,��Th��h����}���iE� ��y9��4�����VFY _ar��R�xbATNzoK%8�~�"x֨'9���Z{(c���-�U��F��dN�ޡ8˔��iK1���ȠD��̬�z��g�8�O�8o���0~R3��~� HTvB���/���꘎ۅda���cŀ����!��n�&�f�vŘ<�Ҍ3��y��D���3��'+T�Ӱ��G�e��`k.._i���UuL����<d=M�j�����kr{Ē��Y�K*kM]C�@���<��a�zn @]�X�Eo�d�QZ���B��l!���!7�Yu*��x���IC����bIi���lbf<��M���}�6t�A�3"���N΄+V�:��ei��z��L�D�m6�P��T����nB�!Ն)��V�v�T1a;8�u6�P�<f��b.��O���a
Bi?� Y?Q���k�9ט_|��l�x(u(V���h�4-}t�*��F����'j����e�-�q1uj7ǳ��rd�c>SX5Xv�/�f��/���o�ƈ�u�d(�Lj�DD;�31r]�|�cu�\���C�8�$��.%M��Tn{�Sߌ��:o�����^�CqI��`��6�$B�-�E�f�>u�^#
c�mV�K귽گ�"��0�]_���D�����d��Ó\FܫJJ}�!g"NH�Za���F-N|�]U�(�$$�؜�n�oO�׵�P}�@��ϫ��[�4j)�H�^�����{_��P��1J�(�Y��W�(�j�q%����me�
6*�|J�Z�1�������e��ޜ7�1�4�����+P�|�RpC��W�bu�#I�6����C�itU��h��[�v<3�暸���ZĘ�)䉴X;?@m�����f�l�9Fc���P�����{8Ybf��3���]"?�z4�Ȯ�#q������~���ۋ���Y�E
�r�e�;����|_�Z=j���>�D���>����.'0~c���Lnt�K;Ε����P�2 Z�E1����9$�k}�'��6�! zߢ��G�]�˟�3�=�/%�����,a����&�j�q����ZFNP���D��^��ZC�,��2>�j��=�IO.��`�p,^2��fB�]��'����Q��,z��L��iTiK�s���m8��K�A��08��ҝ���P��xm��II�\1u�а����p���Z1��,��N�ۈ�՚Z�?�g�# �Y��o�����"��X�-A�ܡ�g*a�s��J�T%X;+�yK �����c�	�x4�i5�.qv�O��1:\�1@u-J�2�b���KC�~�n<��;�f�G�o;T^)�euf��(ʇ&2Du�n%|�V7�T�4�S�g�ިl$��R���]'0�0�� �?\�N?R��/�S�����GE$�W�dԨ��<�,�~�;������� uk���ۚ����5 S�3�ʕi-���jj����c���?��m�����)q.����r}5��њP�$��J��1�1�"�T�	i0���	��0b���s7 _Β������/#p6�� T��
U��M\^y���xt��_/o���z�� �H+����~��!�;u6LƄB�H��*���EI[��b܉ͻ(s�55c4ȭ6�u�_��ց�V�B�`��a�ZYY�9�mƸ/��<�͊V8�=XVJt/���Rr�o�K5�#pa:ƨ�r%х~���ԗF�	�����ݜ�߄"C�#t`��|�V�.��0���)��0==�BV�����b}U�)�H<��gB�0������� �;������hO��w�[�^*�	9%��HhG����~�9��%��������%��be��֝��B���L�Z�F�eP!`Q�Z��r�Up�Lq j�'����iѶaJ
c��Ư�N��֬��Kt<%����=)M�aD�h�J��� J�AI 4���\\)f5�uȁ=0�o���dX���v�;[7��~�E�����?�0��ܨ���Ʈ��:oO�CD�l#��}e�z��˷�b2?�W���74r�z�[���mXDSJ ��R�J�a��26� X}l< zU��o�����`g�73�����L���Ie�@� �>�m�P�9�͜S�+׭B�w b�CL�eg-����͢ŧ'yy�uv�^8"�j{3+�wu�h9�R�R�0�L
�,��1�����T!Q)4M���O��#D����`�X��g��ZI��>�c"G��&rO��� Y]J�I��{v͹>�hMq`l�1$O$�P�%��_y�Ag��PU�#�6Ϫ����d�$(.�<�mnwKŚ�®�E#�w�q;d���<���<^ �b���!pm.#_�1Q6Q�h'�h��<��%	�u_%���k�%|j�[@�%�"R�Z%����� XR����*�{!M��@�-0�A~o!�56�|;������KAּ��TwVgה$�?�t��γC�*Cǝ�o��*���7 ��"�Ǹiqc�tF����� B������g�O�f���n�W��N��櫙+F�5�6 ��3$C�G:r�8S��Y��A��7����>��Һfnq�~Tډ3����Jޞ������U��C6?x�T��UE<A�bH�`�@�������̵�Apk�sh�OG���D^��]�GՊW
D}9�pC��=��fƚ8{�n\�柒1�DE�I����Њ5%~e�\2�A8(~���-t|Ϙ �Y�"c�0�Цʏ���I�Yi�;�	ɚd��S|�;�[�\���C귬�&FX�;ճFG��u�ԍ��"��aX�ꠂO<k��&����_���);�,�'�e��yr���4����V�!ۮ��"O[G�i������$qJ�/L�F�bh����"D�,1��?M=!���,�U>��#Q�����걿a@u,&�L���}���M7�.q8�wA$C+U>�s@��Yc)��zR��$�]]��h
D��FT��F`9Ѷ��&�jL���.}�L��T�x��R�r0������Iۡ�X(�k Hǌ��,.5����` �w����Rmڦ_�%X[�J&���B��N���)��)uі4mxh�8��"*,�������Z�O#�p�N���r��f�L���g���(	P�O�w��F~2��lP�O���|�� Z�Ǽ�'1͎�a*�(p�Ӎe5�꦳v/�	����8T��6=����j�V?��7�����U��K�t�I%)Ŵ�X�>c�����c�/����a����x�������9�G7������*�D�y!�p+>�wy���ua��@��|��*E=�s������a�ޣ�.�+�������%i��o���ЖVU���C���4GW��XW���sY�J�G�3�3Jp����xg>��χ���j�}cQ�w)O�v3���s��� ��LF)^6/'�|�BC/���Ly�y�7���e�/S@�����\�"�xO]X��=���;q#/0Gʶ���@Bn��J��H��0u�S�s��L�z�3��{��dh���O�������AX��R�.���5���L����L\7�J,vl�Xf�T��.��e�7���Z�� [���[�	�D�$K�.����g��������1��\ � q�0��㊼z��g�+,�ڠ���Jq8������ݒ�_2�7�ٮ	q		� �*���1�����:#������O9��!� A#T���q�%�
�����z���c���Hk����ˤa�#��(����x��B։M��"��0�
�7�"/��5���8B�3�cLhD�Љ���U�Ӕ�Ȳ&���/�c�چN��@�$0�!A2&������>�_��+k�>�u8c���Q�6��,�x�eU�}���!��DT1���Ջu�̪^]���؞����6N��)�@V�.�8���qZ���6��_4<Ǒ��ce����s�%8���E	�P>�&JY|8���,�`��%)���*> �L���QE�����'�D%�;N�Ŭ�5��K���������5�N��F�ʈ������6��J���S%�r�Y�՝��g(�
��46Zc��~gu���ȉ�����c�W�������5�-"�Ԗ�"��s�K�����N��1��֗��4Y)����]�4���Tu.��q�����!{��"��! ��"[����!kq�dDy|{]�e����hɍr8�;d��!ߚ7�L�p�s'|\�0����j
~�DN�h&�aZ��Zv�o�Ѷ-�G{�n^əOD����-P�$��(s��Qjf�]����Ev2E�.H-|�a���m��6.�D��C�S������֧�2-3'��K�˺5�bHF$E�}t[";�Ep�����M��Uqf�\�����i�{	ĵ��d~�ͯIE@�&��X�u�
�[��&�6��Ev:���j�����NI3E�j������e�X7�A��>�(;:zD�5<�wS.�/w( ��2Ò{v*Q.��Ҕ�rhL;�H�ʯ��I�_YS<�И�lN�t �l��q�|�h��"�gr�Ŧ̊:z��k3��?��ł�P����)׆�d�[(��>xyԩ��ĸ�����6�� Ӛ��zR�#ٓ�f'�,�0�|3���(1�S�����w���\����5��9�\��nK��������Z�!�p\FR�_ú�B@>=ȏ������ZJY����>���y+"�b�i��U}E3?�J/��o�����hA]}�B�����}qZ�oi#Aй�6������|q�RVxct@�!S,Lw`3�	o��k��ڼw(�R�ă�c6��PI'gI��w��B�[)Y�N���� U�b۪�I��RO�	��t�x���B���˲A>���8:M�!>���G�@�[����<���a����=֙Ռ��(0���/��HX�a[�[(�*��]���|nf�K��k�9kW��8�/����𒤫'�,�R�E��L�����|�(�Ǻ]��OE&�d^�(".��`�]�LMI��bv�X�F>^;��A#��Eb#g���l2����Y[�/�8��e�n�1I0�G	��_�|�9�ڏ
+_���L��~�N��Q��X#�Ѓ�ǥ��mm�Y�[�8��X���s��7��(GOp�B� P��Y�\�(�@5xwW�0��mzP47� pX�d"���]��ϛ�gM.�g4����T�x*������6��4����.)en��m���x�?�W;$�H[�L^a�β�	��/u���!��e�)zC0,�M�������B��YgK�5�zS͸�v)wmK�C�h���u���<o��v2�����:G�8ӣ�/Ki��Qm$!o^��"܁���6&�?��|KX�j���TAZ����)ڛJ%Yt�}v��%�X�[�nNxR4P�n�Eg+�;��d���)�_��3u�E�zo���[����99t�v*�#�Q���z�3�����_���Lc��e�Om�}�O�p	��Jw&]H���� ��S�>��&k�?�u�=.�P�}��� Z���[���Xc"!?$3�E�̊�lѼ���4�Y�Y�oa�m�����S�y��� ���:��aX��3R�e�1
S�!๞Y}�6����"NQk� ����*�J���_2���Ԡ�����xm�����/�Y���"[�l)�GN񲢤���p��Ʌ�����oZ�5Mʠ�w���D�l����&XӠ��=���l�N�����$	���M�l�#���"�W�e���or�a�vs*�۪�2�����%X9܀�/�w��t��$�=Ɗ�^�����dɳ�^�׭�<��&9!�o��ݛ�b�x��t�8��7}ި�e}�_�`�3>��?^�W��gn$��(���(`ncE��h�3v���v�6�V��d�Zj��Z��i��R�#��G%�����n�~�HI�qz��A&	 �,�RZ�A���&���it�Ķ5?�:ۗ�9��t&�tID��¨�Z�-l��h�KZ�[��:��q��ߧ}�������f�y��Z��b�������ׂ�6>(]t�wVv<<�U B���s�U+���8��l�}�lJj�~O����AB��׏��}_`�f�W@�����: �Q��I�jP�'�Z4�U�u�����o��z#����-���w?�.�x�-O���~���S�y�a*a5B��A̋ԥ(�7s��ұ�/4���#-�����l�X�@����!>AeJ�%
vH�4���
�5�b=<2��3Ȗ �3:�r:�jF@4�����99bQ3���/Ђ���GR��GD��#�)����
amR����l��Ea����5Z���V:h+U��Ǡ<^H�;�d(�Zi-A�[ ho�d�4M�� Z���j����8��V�)3|<U����z���%>�t��N-t@�\�$mO1��x�rJ�?W��\��j�:�c6���Z=��>�"���~K7Uq�d�	�$�9�|wҒ�B�D�R�lzD�st:/���?�|�i�_[Ҙ�#(���N֣!�̇�e�a̎���a�å���_�_�N��X�[�]a�����"5�3�bU�j���yW@���jb��<��~�`�J.��έ�3�ho��t��3<��v���E���-��]7��UɧЈ@`$@2�e���7Guw?�O�[�xQ�Q�Z��wJ�,cr�K�*����f8��*#S��O9ʼ�Yp�j���0Ek�Չ��S���>��_���)nY�ȡ	"���yLG��q�.�aX!U�Ԭi��nV�o��WA�����!q���-b���G�H�����MiPܙ�xE�����lX5�&����f�
j��H[�
�Ȗ[Tۿ&�$��'�	����wK�e�/)���7g�4�¼�h�{�"�S�@��F��[ }��)�fL�"+5�ផ�$���ٽ��p�~^����_�Ũu���(����{ZԠ��oE%+����@2�����h�hʯ�.�v.8��놸�\�}�ɡ�ϛ?�j�u����vȹ��"�R�I6�w�%n����a���oR���К�^e����7~�U��2�`�/5�l�I=�1�H��"���v�͙�"�ъ˴��K�Yқ�c�_XzwZ�uҺ�
�8cb|���Z��v���C��Ÿ'���=ǰ5~���{my��Ɔ����ju��Yf��A.���� �;�B�0�0��1Sm�:��,WO���xۣ�j&V���T'���~�_�h�q���5_KK��%ˁ��g���P$[���d��Js��98�n1�
r;���4'��D�-=Y�FV��"ym��hh�5{p^x)$`h_�1�(����]M!i���9�&�ᨡܛ&�u�S����,��6�R�%(�L>�q㚱�����-�]_}��8;��{7Iz��:����]b�!3��s����Z-�re]�Tٿ����[������
��`$����jhT/d�c�j+�vſ��P\r%)Fg�m�HO���&7���]]w�.�����Y�����
.K��T��{�͉T^�m��%9��d~C��#"�訾j�"�V~�Cb8�s���O¨[��G�J�]���?���mǣG31[���b|�l��Ń�ßb9{��k�!��ڹ���=O�<��B���dL�s�L�Fؼm2���:�6�]���-R9O��gW�D@�q!�>V�`(�����F�85�ܼ村A��OG��+�Br�U����%l�ǠlO�y����W����DT������g�LYj�F;u����eivD;p����_�����sӮD��u˜~2�� �Ud�� ȺU*E6�3HMLjxFv�l:���r?=���oP9���ħ(�φ���A��L�,K?�e�,��&�ARL��.�:S�N-�����h�z��	����/�V�32(s٦�\VYƧ_��C/ ��t�]qܻ�u�P����b��0M���*��ҔA�.c����M�j(�����T�ZpL��hq�d�1.(�`�]�#�]�@v��Qڊ@�i"K�Ԯڍ�Z�+����`ƴiS��w�h&�H�6�:�����u[]�Y�˱��F�K���Λ�sa�1�����ͱ��u��Zb��P�('E��y��7	���4��'b:S�cD@n�>t�B�V{�������+� '<�. ���_��u{N����;�S��W�/������R;~���*òȣ�h0�T���Ӛ�P��B�O�]Ҏ����!_5����I&�X���R`�J�Ch��t��Ͷ�����-�'y.#?�����2�_��)u���n��.�@������y����`.̙c��!��V�\�����D��7����d�?�Z��� �[�fV��<����^�e�;l,wBi�����P�%�Z�P�!$�[���>�(���)x%F��zP�	�}�2�`s+g��;-D�~��Y
��2(�p�&�[}�:؝փ�����R��?7E����^�V9[xC�$���ə�>�ʔ9Am�nh������1�u�����(��f�F���t��z1��Z��K��iѻ�=��dE���#�h��J�&۠#�S���(�d	����5����uG(ڸ�7P���:�n8#�uѩ�5��N�CS�xU��U�h�m5٣��j8yo���f�ɖϹn�������F��ʧ���<A��	ԡ�VJ}V�[���^^���}����ꉠJ��9k�~�L�����l+NL�>&$��E�Hw�:Ae�!5>Q/���$����O�K��������d�!���%£{���K	N=���ؤra�̪E�{Mj�;#�)��=*"�9I�!|w���_C��g*`�8]��&<ښ)e=30�%]%�qi0�:�A��待�#r-�D]��2'�jK8Ə���� �<�Ʌ���[:�7d�?+�y���|ps8u���t�5���A|dz��v���h�@ʩ
�at��N�~�N(��RL��R^w@}
�UR2Jvh��T�Mٍ������u͛dO>�ߌ��!�������D�q�%~�@\�����;�<���Y�R���ר nó&q'��}��Ibҹ%v����y)V3�ݻ�
���2Ug��O����[�R^�č-���}H�oܐ��+m�Q��T\#��)%�*P�f�����)#^p�<z�����|���p�`�#��x�����BC9#�Pe��]�.Y�Ʈx����yLY�F��2�p�)$BkZ�=V���iM�0V�69hί1b��?Ŏ{�����R7�<�_u�K��6L!r��v���@L�}��
��N}�V��=mQ�n������r�V�)[��F�.z��@��JI���­�O�Y�!��d���֝��e���<+8��'g�!~%�oJ�{�wͮ�{7���U[\����%Y�$U�~d1��K>
�
�ُ;���9�:�<vQ�U��� �T�u'�|l�	{B�a3-�<�&6��kXU
Ā!
�[�}5�,<�,�ٱ
3�Y�dar*�`�/nWbG/J8�"��2����Ϳ#��~� ����-t&�LL*�A��_��@��qV0�w�Ce�RX%=�l�����$��)yB؄C�� ��B"�@1t�3����%ҦN`"}YĻ��NceO�����i������}�K��ݻç�4����q#os�Y�هh�TH'��Z��}/ڻ|��]޺�bݠ{��O4/�C�J������Df��P*U4�>6�e#k�e�+�A��ӣR�gъm��0�"��t#���������}��Q^�Jc�e~{�����9�Rx%=T)�v�ap�N�`�7�䕆���b�:��� �����i���ί��Ȱ�eJs��d�%�Oܠ{iL���,:ʢ_�kz� �z�۩���G�2�Q��AY�\���L-	6�Jz�o�I��<^�&��|6_9���a�`���"�s�9�3R��{!��{��sY�]�͖y�*��M�C�����o|��73�g���G�I[� �N���=�X��
K�KT�SB��"��5Z��68d�3�l�B��Y��s���;�r���iNǽ��ȫ���g<;��#�����Y���EZ7`���9Ԍ���Vݔ����^{Яhɱ�,��7)nն�����f%��}8�dte؉�Q�)�������zE�^�ޢM=:wkCP��d���^U��j/�O�Sf�W򧘩�XR�W"�@-)�Sh݉�/��o�]�z�a�f��x�"��V	ވ�s���o��:�8.R5hJn<K43AF�Z|[����?5�8ύ�F�mz���ԍ!*a	*�d=���0H �AY�D��X�ᑁhw����ٟi��[F"�(�u'dF��jC�s!�I��ٌ�|'$m�"ú|�!*P�4җ�(�IG�H�qA����~d��e��E+ X�}��3D��$�2��;�&>o��)+�o�g���} ��T݌���[��ۂ��G���[���r��O	�&n�d�r:��!m5��G�K��c�( �G~*�~�o���H����N�.}�(���_�J3Q���=IS
��J�:������w���F�}Ϊ�<y���@QJ �zLnډ^���+-��L���p��8U������w��+g���Y�S�M!��P�ޛ�����H'��򲼀j���m@�į�. E~���CRC|شOqh ���Lf��ҠL7�L�}Sc��-�c��-i��b��Ƌ�B����9�#��Iͨ��%��<%V���������\����%�"A���00�DXܪw�}���S�M��������o��&���M�˴���{��L���`H��� ~�y��G�yg���T�K+��W��t��xƈTcp��ME[Ed���4lk�+F�H�U��Qg��:,�;�l0Ǔh#7e��w��?�^��4BGG�Mk3d���w����&�q�UM!J����e�v�u
/]��2/��w5�?�M��@�SO�C��\.@�>�r�&��B-"�G�G)U+�|u��k�h���{������_�n�eq�|�I�E�Ń�8q�6LZ/�4�z��Om�������r�9o���'Z���CaD|G���}C<+��Ë�-�+RF>���Jы4�����d�d��D���!ac�|i�`��s�{��ĕ��S>��b�inE�M,��7.b䝱�=��x�E@��n��=Ksv�^��Vd��Չ#:�u!��ࠣq�L�S(
7'δ���a�Gs@3ۻ�jlY��H���31���J���)��$�}X�S���vQ*�e���u��Kp�l�ft\�!��iԄ�
�z�j����u��Bd�w�&�8�<o�aP���Z�	��$g������0�;����O�.u���͒7��/K��ٯ�d7��{��rTs����ͽa1�dp�X���b?�ƿ�GD���]$������ڣ-9f��c�wzR?2f�1mMdJ/�#�j�VC�T�ʹ��Bӑ�C���I��U�{}�����@f0a����C���9���ƢX>�U�	�� ��#��:�4[E��"?�9���8�{��H�?��(�x9�x���t�aYdش\2Lv%�x�wR�?�wͽ]�	*g*��^�zE��K�Tr�������D�!մ�xr��IHȯ��J�����PJ�4�,�B-<��A�=��>\�d���h�]P����r��st2���aY�I_��:�%���g@�z&S֋�C�~�J<�&.J�%J��ӊ$j;g��N��+0��X�����w��$�B�qR���������q����lY)��^n�[J��ٓC�(L�ӕ[���5$S|d�b3�WӦ���li�+p|�^�C��ЄH�u!{Uj�kXX���H�������h4��˃�j���4?P�W�d��o~)��٭�1��6���ի���ަ�%ogzU��T'�6\�W?���I�-*���5��� a�OԒ$����s���L'z�O
�6Ts�\Ӥ�QY�)��f�0���V) ��A��/�+`й����9d(o�?k�o�k�
�C7:�3����@6�����w��Q&�B�;����2dp<�aq�G���btA(K��N�t��z[�]�Plp�+�AO�A�S8O2Uֿ�x�����$�%�k�r��yd�sЭ;ŗr�\����ѡ�����,la�dsL�r`����.d����Mx�<�~U	��������A��y	zb
����)1
����T��K���<I��Ƅ�H�!Tf� `픅rmg�=J�z2���(�ʥ�}C���<��� )�?_��r��H�����}���uď10Y��͟�.��x�����������	S���^����ލEF>h�w U���?β�ƭ��)<�	�ѱ\nG�w3'y�X6'���	>ǩ�7p4C���-qK#V�I#͋��pȁ�B��s�^�w͌&�S�G�7�8�?�����k��|�ӹ+%z�Y�PO/�	� ���2�nA�6���ʚ�R�u6��p�h��>Q��.��)o<[��.����8���L�e��r�g;�d)r�R_'��\�ۻ�b�6��!�Ī��ר�6�z9��L�Hщ�]�Y\���e�ԝ񽊦��"3�zez�[���&����������MxP�7(�����%\V����X��~�(�&Wݲ�4�@[����G�T˜4�?�S�B�Y��Q�Kl���`�|dt���}�(�]�{�A	@��|��J�qBP�5��G}
�[9�ɡ2���;Y|G���rt��������2�xS��*��A��[@mSk�w�C�"x!�$�wo��g�0�s�>�7��KL����.�1|{;����+�[�������~�E	)E���;3o�"Y^�~Quu�����H��c ��O�t�s�I���TC�
�^I�1z��cCa5���[n��.B�5h�����N,�;T���Ry.�a)հ�k������#s�C�]/k�%10 %a�l$�Vq�^W<��Ý�A�gw16	,����Jȧ�y_��d�6<���^k
���I��H�0�������.��s?h%׽X�LTTb��FC�Yp���V$pf\7�aN�y�<�ɥv|H��<:�����=dS<�P�cG���7��IـC��VM?���rf&���)�P'�MAc��=�{ao�d���Zc��a�1.q@��� ���7s�w �ZYf_�����e�;^ILb��n��+u�t�̈B�L*�"�)�xH_�	O��U�F�#�L�)Nq�Փ;P�+c��`��۰ ����z���6��r[�]�;ݧO����9�3�ou�$�b�@��B~�!
�U6��P��MۯߗBc@����[)p��=���&��#K�1��?�� n�P���e��>#�R��S���!4�Ҍ��#���ip*EZٷkkP�]
��J�<�¹�O�[.M�ɌJ١�=\� |g�8y��0�X�Ҹtxc�ӹ4�<Iɀ�t&���<V^~���C�R���\��W�����(��qgѺ�q�^`#�i��RW�7b{s)����ӟ7���7|�:E�U�[q��M"{}N˵�����C��ϙ(O��POr��`����>eo-(�# `U�C�.���`�?#U!���<{�4�;йx������wFNF���R�I s�^�y��T�� k&�1���|}�'Z�~ǉ+�Vp"gU�.�/�a��5�W�Sǀ0�!��g�}���G�A�79�52�B�������\c���e�|��\E��_��8�P����84��z���r���C1��4;��^6Oi�fV��PV������!4�QE�`^�Ս^����65,�B�� ��\��NxBf@�$�j������4²��䬚��poI�.l��t�@0�&Nu?\C����=�j'G��~')H����&�H\3���2�T��Jc�p��-=���TU�?���E_%��ZV����0�Vɦ���6�}j�
�� ܳ�>Y�7y6t���HJǬϊ��5~z��dX5w�te��QRe٫�܌!���6��G�����A�X�v�;�������z���u+�Z��i� 5a�L�����KWէ�[�!AÞʉ-����p�i��]yL��'_**V���ځk��-*�P������>f�nr�{8�A�*���jw�N(�
�w"���?�}�.ގdY=g|�92���wJpbb���6o��_(�ioH~�D��@XX]���m����j&��)�q��5�qY�v�-}����L���!Ո���s���54���Z�1�8�s(c��\�ؘ�	1Fs�[t���&O�.�A�[W�.OY�0����;y��7h3;��S��&�����kxH�b�\p�bvDVܛ_��b�8;�6�m`�O�J��P�&D��tL���kŏ/�8��k�ߛ�����Y ��M���8�*��_"A=f�� y�}mR�x�V�"0C<:�e�Iz�``&8�T$�aH{?.�dA�r��R�$�зt��E�t�	&"��ٚ������J<��|��*��56RG:��U���tP���{]�7�J5^}|<�Av���h���0?*0�T2��*Y��w��!��	�X�������N���%�^��YA����ұ�DT�c
�~z2�Y���Y9��!�#Fk�Ek����!�~�{nh��jt|N��E�%m���X��*j�U��n��sv�V:���,�'��>��)k�ܽz~
ݞ�P=�;�U,��A��8bw��D�����ߧrH��xO�=	|����eE�Z|o��]�:u��Be��:��V(t�#���{�>��#2GS��z�X���[ ��s7���$d����D�����ү�&9�9ҖӳJDv7Bg��3�����1*\=���xy�a�%���D���"�/�.�j7�� ��$�9G.�ϥ��<C`S �����O��P�N�+��5N�_�� oc��=JE����ޕa\��ݽsmY�y>�~���umP�x��w���e�ؙ��c�n��(I�����{K!�f��ۋ���a�����p�s��_y	T��t+:"k<���.��ָF��� �����bρs��NH��z�_4hm�k�m�xܖ̍r9�;rUg�5�`'�d�m��-}Bw�7�
�*�]��#㔙��+��з�!��fg�a���*M����ٔ��3��HR�� 28w���G� ���Z ��ؓ|!��»����R�&�.�JKS4�<�#����������P"�
%��U2��}�
�kg޿���I���Y��	���Չ/�����\�hoiˆG;�|��I0D��J>q��
�$X<dp�D���7|����,��]���so�#�̻�U2��:|������o�3��m�a��g�(��>p`�4��X���,�w�Kx��}w@���Œ�sB�/�#i+}�[��|��Ǒ�$��Ȏ>���k����z��)���[�d-�H���y�Co:��[T.�L0�\֖n��t����wD]?=+{��Ee�YCb�Ͱ�&p��?5
��q'��.:J���@��kܧ*�	��8 1>��Hi��#�����~���u㿊�U(�M�b�څ�w��b�1�@���3"�BX|w����ioL��I�]^b��xd�0hdueI�ٌ��N�ѩ�D�}����S��=S�z�=׳����*�N���g����=�	����� ��ב���k�)D����7��U��y5aۧ���I�����Ակ�u���S��T���~�b�槥U�?%|�c�z�t:�1�qMC������~���b�?�pD{�j�r�C��io꓿IzIo����$:?XG�й=�V�����|���������l���&ӹӯ��ʁn�Π'3d�z���|�B)���R��Pad:8�~x���-Bq�|����
�*x�DݠLw�����&>����
�c����woy�=i�t��f���jU�1m��F�&A�������>BM�`�����O��Uz�|�Km��r��Q�<�����������7��%.
�{�ܹ*�P�KE����'?��:���Rp����O=��K;� _�� �a¡�&\B#=�3^r�2̛�nS➼i�.]��-0� E�И7�����@�aL*K�\W �C��7�!6�k�7���1AT��>���H<��/o�H�7-_C���1퓩�2��ʖ�s�{�b��j1Vno�M�'�֣����
��8aY��qP IO���O��S46�;���Dx��A�S*['j�{@f!+r�P�}9��ڕ����f ��]SCث���G�Y�ڭ>���T?ҝ��cX\
�;O"���PZ`ꖷ�ՊVDy���O�,�,=��<����@	�X�X���@2�F<|1
$D�eH��b�a5,�Q+���E�sdZe����4Ʉ����1�Q����<(�7a��yx+�`�P�K�Ҥ��{a���t�`�Q*�+�O#Sŉ�샭�R�n7a+��f���DGmd 
)�!v,�#d�Y���պV�䛾죎�,J���V��܌}&�m��U��U�Q��㲴��ws���H��?Rq,��3\���,yZ�g4�_�'��A3!�`�f��%f[\��ɓ����2�t&��1��U��m��2�������&��v�@C����tG"D�/-��(W S�M���!N�(�˖t|�S�)����E���k�A�\(�k�;
_u5^�z��B=��;�ݐ�ܱ�SJ���Q0�m��Nvw~��̳};�j�/*�� B��#�Sw]��[d󴌇�({}Mi�1X{Yث���|x�K���l���BI��lO�mZ��b���tS\���F{ssJ�]��X�G��(��cqgޯ��P8�|�7%F��u�66���n�Kj:T�ח����[�_��pp��d��:{�>.P,�Yg�]��LsرOA��k�bo5���V�K�I����%\]�te��;U���C�f�a�Qd���Qy[���r7��N}{J� ��"�´�0�k[)Ҡ%�?���������&K� �V�VH�W�8�@\f=KG�4>\Z��ֆ���c�zDMwt$�]ڈ%�Rۭ������8�D�������ħZ�J��np�����B�L��Ta�wAIOnc(=͖�(�I��h��:���z���u�`M2�� ��6�Ə��~��d29����5>�V�*�4����K���#{JtQBƷ�\�R�,a �����.蒇�4���\�������}�wx����*�zR�:Z�Μ�Rǋgɡ�{�j|�H�����$�ɔiJ�����;��p@ 3�~��OQB��ǲq{(��X:i�UK���7;�@�F_+!��%#�:~G���~[C�;��`�D*y2ѳ��.��԰"S�9�0p�	N�]���zb�]��N#j�fGdA��t	��${	ƕ���bU�F�� P8�?a=PTҍӵ7�X�"�/=�/��j��-'�N�
��~��nJQ���N��/Eh�L���r�[r�$�
��"cK,rG���A��߸KAk0�Bptm޳��«aa����u�2�5L��!�\߱c��^�$Q)XDm�2�8�2�l��:Yf���<��o��GN�vBަ}q毠��t�`�6��$���$�m���Z �ZoM j���'�3�6�?$�����f��<ꮢ愂Fd{���!|P���E�Ψ1q�Ӿ���Rj��y�vn�aN�e!(y�-	��U�l:���%f���=٠<�v�'��PNn�W��A��%%D���@����p�8�כg1��趃�"MH�߰�	\��j2Ԗ�@�k���Ŗ�՛F
Bm�o�0��c�����O1�	�W�}E�^w�j�S�d�5:ݦT*�^���u��Y�0�<bJK���i�F��l��$�2$�h��A���a�A�mH�f��ՌZuO?}7��h�0,�Z0J�,��+'=�*p<���1|�f�ѕe��!�����	4z�0:v�w\A|����X�{x��X�*>lo�ė��Pe9��;l�Ռ�� 
PF=����es��Gľ�6�U�0���S�bp`7Dncq�����/=Ct�M�&1�}O�s:��֤:&<�8�lhZL�<��/�L�MJ�Kܪ�T�}�a�� �<�`k35k+��+�(����-]?YA��	�X.��2�+Ƃ�T���� �T�!�<�=�sjy� ����(�<�;�"'���v���N���?�r�e.~j�f�n6ϥ�����ʙ�f��Zlɒ�H��8a\*�&-F'{���obThK�=���}�����X����FpD=����0w�jBȳ
��ώg%
�Ka�g�ā���I�9��[b�o>�~�+=w���謠$2�씟N*���J�uth�H\���k�9�{�XC���&����q�K*���5����]�q��^ :����|����3��#R�FfY��=�}S�R�q!ϑ/����:v�_(�X��G�4k֨L".����\���W�:�b0�����h���X�T���l�i�IM�;F���+e�c\��ZYR=Ɯ|8"���$�MT�"!y�ʉ���R|A-o� Kǟe�H򪑔�wd��kU�qĵP��o��[`�4�K��l8�ܳ�5�&��̌��J����l[�:�*�"W>��d&��oZ��s7m�J� svNX�1��Í��EV
u��RV:��&��\��a>x�ʖcx���1�k!肈}����m���Wtip�lj����c;#�b�������Y������3,���<F��}���4N/B�Pݠw�e����*_W;����ѽ��8���'�4��2ǐb���7s����9�2��i�R��R�D&�<l1s4��c�Mli	Mf*�!��J?��S�`1����� ��We���!��C��Se��=(M-W�g��V����F ����sx���ϳ(<5�{~t����<�%�����g�[�=
��/�� �Q>�(�����7�������&e�z�BS"RdcP������������5^ƕ'÷�m�j����׭y�2�.Ǆl����[X��̐���Q�f�,I��>�a�������I��|��s;�ur�sό�-󭲆�%�1?���n���)O#�>��Y:p6�I�r�e�л�{�NFq܉N��$Ӭ<J�Q��/��޳a�Z��T�"�m�qk���o�\}
�aK䓐�g^�����Ҥ��$�����È���	U�`�nC�'h�3-D�a�-#�A�ޑ@�����c�Ӱ�4V2ulU�eB�����.��!G��<�{B.�>re���ݣ�p�� �ŮcV�{���\Pd匕	s�&��tT�����t����Ǵ̦���A�LHV����ϴ4,4�g>J;?�b��5��6O,[˝�RYM�g2g<�U��T|�q�ϊk{=�X38^�x��L��lw�)..O����b���U�*�we�D*Ǉ��U�ތ�>~���O�|���S��F5Ʌ�}���huo�,1q/��%.�q se.t�`/F���J�l�v^���:_:>D�N�O,���N�q�ń8�GC�_�?�Nd���O�NK6/��?�ss�&e�Sj;��qi�Vk!�+[# �h� �@O#m:���X�&4�3ڳ��(Yd��=���G�zT��/�I=����d�A^��Y*2��	TO�|�蟹-A����v}�yT����&O]qlO�^�g�G�O�����B���9&����\�ގН,��JR���
4rR��B<WQ+�5�]�G���T/J�
3\�.k����P�-La1`Оs�1�vAX��v��[h�;:��o�)��3����X;ƾ�Z~E��Dcd�I��z��� A�n�Oy/�;�N\�x7Z�I�g�A��Q���a>SZA]���{�E!�?�e��3��C*;��8sk�$ҭ�U��������F�����L�s��[E܍�MJ�W��S1�:mw��F��8��y�rص7���%��m��4rJ��9t�K��Q���H�x��j(QJ�o4y�����g�?�,��0�8�DD|�NM A+�V-�t�	Z��m<� [o�"��]�-�����,�pɦ����E�~�H�S��ӻ�CwX$����\%/�CAU�u(�H��`��r,�5>�9`��۲�,�-ӛu4�>Ж*�~��x��yX�"km���<�`�es�������,KR�h�˅Wm�
ܱ�T,�x�����	��<W	��N���o�e��xb���j"�TR*�98�+�1��Xu�<O�J�(.�hel,J�G�%6�:Sk6}1����C�&�X*f���oY?����g�� �L[ge��bʍ����9��#>��é���{N���)���<��E"=��Gݷ��6T������:��@&��8sY�(SȆ��$�~�L|� yRh�[�0+�-q�(��ɮA������_j���/���z�T��.�|���:���?�N�!��i����Ma ^��n�t(l��o彳�G�+7W#s��:�d����L�`M�e�~�T�r�m�'����6}�\��H���+��!o��w�Q����2��}��{��C����Cq�V2J��>z	;��	�	�� ��k�V~�h�;\����!
C�`nL��xՓ�IF'�?�_�")u�)�bL��f�Щ6N>Lul%�Xϸ��x� 
����A҆��}���~|݂���/?^8�m_�d11i4g��X�c����*�=�fu���~���s�ũ%Z�*-F-#vR� �:K�z.�ρ8����\Sq�H��q���~�og5t���<��'� ���C�z��UR���ep�-��>b&3W���e�է���|�3��7��Z�����sGs�(����[ד�[ �aE�������T�O����6i�pyLFa�%6Ñ!BL�+[���M��z���Z�r�X�\��̘����rUG�N~�#_kb#���||�d��۷�S��E���k/�����Kt98J��?�2b\p�����P�Ù�L�� �Dh�Mz��}#GQ�����
��]�������s?��_�V� OT-V>�����c-���ӹ������%hs��0v-�ƹl����Hr��7��4W^/��HU�RɧLI!s' &� !�1I�}Yk�"`ȳI��_��MܾG�����%�H��O#S@�^Q��M~�ۑ�X��b,r+e~���b����6����j�S� �2B%�XB��5��^�#�(6���b^�\x^=�R{	�1��5yS4y�\�Lbmy���]"��}��<&Z��<�{K��*�v'N����h#W, �B�Ԉ,�G��j�T�����z�yC �SZ��'�g������G�-<|	�)���qM�uԠ,�`٩�ŢT]��u�:�Y9X$���7ڭS���&���U��D�UX���^J<C���4W�ce�h��K�ģmf-q׸��&��!F�C
��,����k���]�!�d�XK=�%o?FQ+5�g�Ѩ�a�D�B}H�V�V�7�'eV���AP�}1�7�X�#�	B�E4z��Ӂ����OD��3FqQ�4�CL�3����͊�K�d8�#��.��*����Z��p����Ũ))7���\knm\AȜ|�v��O�r��T�����帲A B�rk,<���DWh?�ܻ�\�/Fp��z�^!�x��l��d��]�0j_\�X�lP�W-q��見)��+*٥�ЌI�40�t�ErtP��(F�N�b 2~�������Z�v��f;T���_;V���#�C�����Qϖ&ˑ#�c�#�Jf@9�����Yy�k�/j����:΃���uwk�n��N �y���(��B�G�UJ�f������z�e{�s�kr�r{>Dȹ�?;5|`|Ķ���yR�w>���P�P�gUT�%�R-�S�{�M��=�n��KDi1�"5��8�V����u��	�$����o�d�$G� �@\)���(��4�b��ɞ4���y���Z#t*�����찬�wius��ĉo	0�"���vθ�I��1%Hk�����oј��rD�ӣH�h�ٙV��1f:s̰�/�}����;���P#j1�����-�`�_]@�E�@��;��:Z&�'�XV�ɢarqE﫩�MoKS6�$�@�,\q�ʲQ�;��_�#L?����t�V/7�=��(5�va"J3ŵ@��՜*�u<�~��Ir	X�(���Is��%� w�OQ��M@x���>�7��5�"��՟:��' $L�i��?(�`c��B�r����2�s�֚��cF��V�_I�Y'���ُ%�o���3��Z��GG�����͞[<�3�8K?;h}�!&�Z�w������e�R\wi��6��~I3'x��8�:���,�K�I6�/�apR_��Ե��z��ǥ��U/<��i���IOĖ*$�t��:�
1�v�	& ����B9�w�)�U'�/�<�p^���[�ާ�2Ω�L��f��۳�e����F�Vr�ker��$�~S���������$s��	�~Ǵ*��fq!�B��v��a-�AfG�j��O?��C/�%6��ps�EH�j�.X+C��4W|��D
�%Daݷ�}�k�w�r�W������B	MA�}�7�Kk��o�5t�6���`�=+��)����ׯu#MyPrTcADO�F{�,�Yݮ+P��2n��͞�a���VrP&�5�|�'Й�i�l�*�Qv���F�O�L�wc�T?��C��H�x���F������Gɡm�_��|~� ��lq9 +Ih�E=�ӣ��:����=�1*�]~�S����џ	�����DÙ�8����σ��TV��&�_�Q�!�>���V����F�4 
�0LnӎW�/�k�z�n�~�]&�}����h-K*nM�e��=������6!~�07�� S���xNt�lz*JLC&���xʩ��z�k>u�g�mM(��e�a�
��|����@��Z�%������&8%"������W����J�*���ժs?��o��MY�g�~��rw�D����:��fg;+�@�Qɴ��וoU�o���o��7���\�lXSX[e�7�H�HU��D�a��v-
�FX��+�����Km[πC�vZb�M�$	�nd�`�����0�>p�Dԯ�4M����a�m.16"��f�}�X#:��ɗҶ��)->)�"N9�SA=D2���$��v��b���>8�3��w>K@+��H�����������"�7L��K�櫎�����W6�P-WA�..6��P�P@6b��*�fm���;PIvƂ��˄��=R�<W0d����_�6Yzo�v �~���R��*E��h�(����೺�H{�_}d�\�����֩��*�S�,%�gnG7UɲFM�Q��,U4�����B�Ԑ#imj�E�\"K��sP��W�m�@I��5���t>�<9�m:�����:
b� �]f�������)��&c���*����`r"���pd#CGt'�ŭ[����2����M��
0A�,K�)y?��ԉ,��#��H��`�G�{_�Ɉ���ꔁ!QaU2jۚ�(���ա�B��L�qT<��D����my>~�,�����V��ȼK��ʝ���m0�෿������D�M`���#����T��܍T����6���|!������T"Quy.Ŋ(��
X�'��#�ʍZ���T6�~:��:xCZ��s� �x����_ &p=�� �ҞkޝFh�(;�,���|������n;�t�Q�y�����-�~U����˥��28�e��ft->��`e��$V<��ǰ�d�԰`oS.�K���9C7�-�Y`�vo�������mc�`a�����xC�d}�����ٲ��܂�E	va(=��v���К�)���
6���/�����d�],؜�����C��텽���Q� Y�C�Z���T>�
��OIc��_��<�I*��;{��ނ��i��DN�F*���8\_��R�{s���?�9+�8����eʾ��O��ʗ��Y�(Nf?�zՂk����#��s�ئ����s*����"	h���|E�����Sf#̨�3�V��+g�2�đ�|@Y��*�ƙ]��TsKZM2.��	-=Z�1�O���L� Nӫ��mSG@k2���w^���
��ն�O�0م�PG)�oOЎ �Y���#�T�+h[18s�����AIH**�����5���m���.�ّ b�6:y`ֵ�	� v<���+�0�u-� 5qK(���$�t ���.��!��t�bF~��V�r>ǧ��I��	?���pg ��!�x;��ϑ?@�g�-���h��?@�0�Կ$y�l���]v!Y�&SJ������[�g2��u,P�EZ¦����CP�ӡf�o.&"LS2PI�-z���"�#v�(剻*���� �6�����i�Z[�(nWԓ9�v�G�+��mp=�Œo��� (�d����!�!V��N8U���ʁ���;ʭ{
7D��𣜴x�u�CIhǉ8h?�me�IU|�X���z�v�z���Z˩ �p�/�񁮃D���,�/XI�	��lpv��,!1�h?��R5�f1N7�	�s	�2� J}��J�M�ΙÊO����(��