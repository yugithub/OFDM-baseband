��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛdp�����/P?�RX�)�.�X�+�SZ�ð���өNl�7�Θ�v#����;0�pP��	,~�E��C���Ol:T�!� �mX�v$��nq���^*�	~	��܎�K��(���w5���Ƶ��D�ſ��9�AV�c����h,B�!�rW�.����y��὚���d����	�@o|�#e���ڶ����-��b�vzv$Y5����	�|��d��8j����6@4f�t�U��EC8{ڣl��/�pU���3�EZr	M�؈�����ҵ.��O�T�ZI�L�O)?����$ O���v�K�z�<z��~��F)~i���$�������s&ŕ�'�mX/?��Z��i۴
�����ۊX� ��h"����ܷ���AZ?�@�	OK)V��b[�W@�圭��E�-�ed*}-��f��������sm���'���$�J!*0���O	�㻷خ9%��DM#ʒ���-�Tl��[]V3�ҁ�q^�5�@�Z�+9�1�B��>����!���M,�r�Y�^���)g��V��q�+�P��.-WN�1(��Qx�ۋbU�D�J��b����+� ��uh[���d�7ς�b+6աs�z,u��^���o��^Oej �"IL���82��&�4q�}�1��Fp�9$�Qdmv�-���v7�ܾ\>�iܞm�)����	��-Kh��NO���_��/�Ǎ�"k;�V��,������K���l�@#�0���Ԋ�݊��\ACEk�/w�أcrn뉓�Q2M^��À�Z]n�M��:?�
!i����X�w ��w�!�!s��ư=O�K����]�*:��:�٪w�F�6�v�Ћ��ܥ��f������Ŭ�t�Ѯ�n�]�{h�v5����eo�l��ۡ��5l�<߽B� �iK6�{�Y� "���>�����~1������s|�-e��?i���d���Z���l�Q��ӎ����X�΍�ȣɄp!p���=ۋa���:UxrV��FsI�1.��	�8���٪�ț2oif��$N�K���'��k�K��죗z����XƔ7��MC>�[8\U*D�Mgq7D��s�u�u��ِ۪{�A�Ի;�5
��D[���c[U�z��ю[�ʪ��]���]a�-�+�3�½�_���[7W���P�,9�f�R��%56�k#�����C�uu��^H�S&��]-�L���T8@ZM��W���k�[u`62w+��B~�ܔ^P�5O�d�'1y�I���2k�Z�-�Z�C�fp֧� ���H.Ǔ1f�_���x�����z�H��ɻS&mʏ5�S�_�]��  1+Mi"����g����&i�������o�ю���7��=��{�ТS1pg��%�}��j��T D��d�����V�_à/���[	�2O��ѓk�R�(���o��]y�Az���ݗ��&���[|_`��(Fo�4W����֎\q�B�G"l�4�5�=9Ѽs�Z��<�Q�����A��UѦ��$�ڛB�L�_�8A�	��"�� �L�Q^ 1��!�6ǋ8;� V΍�{n�����L�<!�"�*Q������.�L�2F/ELe¶�� w�'�s��e�y�M���m�O3����"`~<FR܉����6n>R;�W$���zRz6�1� ��e��c�qB��Ҟ�!�km��7�u�Ѧm]!Z@	b�r��6��>r`8���by�G!�M\�v�ʗe��6�7re�]�k����}����+#N��+xx���s�)���O�y���u.Z.����dg��/��9R�i}i�뼁���?���<H�P0r0��o��j^P,N���(����=\�� ����΍D +���6�M,`aB�Ǝ��T���z�@Qs�T��f�"��"nn��KJ�
YM�$
��^+�bo�'��������Ռ�m4�dN푟�3P�>���]<���NZ��^�����W�#m?�+��� ʠb��x:K<rK°�.�ÿ�Bti[��]���˼#�bYb�y����F-7 &2$�{MЇ~�	��̥_bY���Ś|����i"0�y|��)K3Y�:�L$xk�|��ت�a�:��"-�	�C�����U�����on՛5K��B������4�J�~�H
�X,�L��ӂ�	�Y�h�Er�@���O�L!��a�:�A}��܌-8,f����[�ȱE����d���5��݋ѧܒ9��:�%�w�P�,��Sr|�]�Z\!d�^|`0pYYa��y�9a�¸���4;�`��ӫ��f�0'[?UCq�( ����*٬o�EYC"*���]�:����>�G{��;�Bm��װ}^N�݁ñ�G�u��ol���}__���;۰2*@w$�{v�Q�q��SLg�� ����� G֓eЎ2n7�'�.�9yE�t��?���]�b#`�r��{�e���t�rl�3���w7Q$���O�9���Us��w�H�FܫgR�?_��L�I��7�+c��[�B�~����ջh�O����v�܎ۺT	�(�Տ�Հ[-Ʒ�Nݟ�C�ےr�q�rsK���Z��	�3/f������T ~ ���L�`�X Ϩ0F��� )�;:Z�ֵj��E�E*��$�/D�3Yt��6A�5b&����_)�p�o{�әF��l��'��c�ɇ��V,�۾�S��x�>W����y�c���E�Ox'i��~d�#���<�eT�hp���NP�E��s|�i/�պ�zM�"gl�d��ou�WM%�0�wo�P�TZ�3��K!�q��V�:�*j�b���M[�G�9L� �ᦦHa��o��H[��y$f�p����p�.S�yZ�	��� ����v���P\/]�>ĕ��O����٫���;M����%}�jD\!�ri����?;Fm٧���Ta�,�4�b�B�I�W���뤙�@�x'��������\��e+��W��������0���jp�R��}��5��`[�1�2�r.��n�9pF���;�_Ak���! Ӵ~��Jp܆�`-&�.�:����
g�̴�t��<k�^��t� ��e� ����C���L\n�?�sI�C���������9"���~0�����p�	�Y_��P�	(�7�C�M�g֍E��M�Z�!��.(��?|#��	l��z  n�쐧�O[�ߩU}����xv���r���<ܾ����K�gԣ=b9�������pr����Z>�o{�'R��y�f�8Ju>�$�k�����fvwv��'s�ɜI~�n4�[~�$���*S�L�D��w6���p�$�4�ѱ�[:K�G,S*��i*�jd�@|�I���֛�P�ل�2W1������ r+�%d&������`o�%�I2�w=�[�!�ڥ.� _��L�؏���@��.�Pb�\\�i�ά�������E�E�מ3�D�b�{�Dڍ=�����(6C����B2|�%�<��Z@�k���b�!#2� wR_G�{�W�ݹ�?4o����rb�Z+�IK]���o�㉊>�\������hL��U��h�՘���ܸ�'��1�#��f�)��&�e܈��e�U�4�����z�eX�K��j��v!߅��g�B�Ś��/uw}�'g����E.r�*z��p<��C9�}�eMÃ)<m�͊�W���uLI�8��a:d�-���2!�ҙ,$E��#����^�����B�K�:ve�����Bl��U��xI���#��& x��z���G�6@e��\�Eƹt�S�:+_�q��cCL���&�;����a��6��G��TMOc�C��$���+�q����v{�t):�J��B�����e�?%ܘ����Y����V�ԍ���I�#/�Ud��"�f� ӂ��AXrz��ô�p����t�lQm���"�r�*���tS�W�?��y����=���h�.���'����Y�ACF��MJ��@�)�$���A#[-s�e�t�%�X#�g��iw�vU����c/���.��T�w�����R�_����H���7�OC�s	�=�����{=�]tn�d��,s�O����lb�E=�ڿ��Kv�*HIGh�c�M���9�B�Jգ�u��a��N4���	��	|�:��˯���Sk��Ss�<�N�~�>��K>4�3+7<�ݷ."�3���A���ċ�L/~Ԝ�Bd�D��/P{�G�$Wcͤ�t��Z��Z�[�
=J��{�}�1�#����!��]h����%қ'[�[r& `/��M���{���LW���KH�Lu���"h��N��~�>쨿�Kȟ������Q����5�(�
��#������*@�X$�NYw�5���R��b���U�c�K�2j� �#�j�%ϻs�ci��(������X�meCv��Qw�;y͵���p���u�ϊI�ی�S����G<>c�:.��BE�c���~t�"�-���v0�L�i���[��/��Vo�Ӥx��
��5g4������'�O�t�����H����r������BI�3ZT�5o�d�<a�|o�;��l�f��7��3s_uB�\ k�%�G�i����Xh�Uvx-��˷�9��:A�-���{����s�%�m�ͽ�5�%<��-o8yکm�yur�%� X\ZM+4�خ��P�)�G�������:�t&��y�<EO����W�_Iݕ(�6[lR��6����GU��ݽ��4ěa�ӌX�������P�~���<a���G��d��M/:����*� �����y�t��f��Y� k7�<Rƙa��|н���b&Ѕ��hX�3��Mv��������]��R�]U)���ѹM��5<_��7v.�s>��(���L��� ���	��!�P@	ٌ>�3Rq����-'4��ȍ�x5l7�.�DXoY��8��/�X7v�	��e���*k3��;.��<�7���3��,K
�nwP�����B)~��2X��r8v�j���osy��S1R���(ٽ�q:[�-����|e�Q9�2ټ�`�ȻkP�
q���T@�����۸�ڦc�J�b���$2HG�|U��7Ѝ"A(e�yC4�������_a���m��}d��g皂'w�P�,4�˭��"3/�5G�>�y�Xt%�6�|�[��O-T��g�o���IGS�oRU{J	(B"(�j���29��N��� q���k)t����A��COr԰wg4�8�2��=k��݈M���
.����3N^*3c����b��N�+�4-UgFhˏȰ��*��-��yA�286Q�*'o��O(8��E�T��RL����wG�R��a&~Ƴa^��j4�(29&��lĭ]��,z;�� w���zך�p�z�^݋m+�D��>23p��y���5S��^L��v��y�t�1��N�sX��./��oW��5�Q?�g��Q��s|��gO�.6�\	O��FA�aP�ū��\3<W��w�z��c����t�d#�i��I	����4�l�{ k���M{��.��g����V����2�K�q�|��j1���$vor<,;%�:�>�\��@M��C���_
r�a��l�G�d�b"䷩D�c�(8?��g�$..�V�i.��-)���_������p�Y"}������f~�k�����S"*D���HI�)�����L���\�%��L��W	�=H���Ҷ������k���P"���E{�b�c੕9�f��7o�I��>2��5c�>�B���)�Ⱥ! O�3ĊYJv�{�=j�i?����ۿ��o:+�w*��0kU�P�cs]
G`w�9�y#�U��nv
��}�JACzX%��v�L9S!�[��H�H�L?������vB7SI��h�/��:���9������0�0�%���g�sCqPH4�)qd�UZf��T�jẗ��\� �F�8YRxZ�z�p0����ҵ#c񱢉��(0+�ga?���Qf�݂���*��NY���9(U=u�"
?��Ͱ��	���
��з�=c��e�?S����Q��ۥj4:�D�Cc�h��OK����rݬ>�N南~d�Gҽ|��	�� �ѭ�46v�;Ơ�e?�4�����gf��?���>=��)��A�������7�1����4EG= o^�93�E��f^if�y&�dS�f���v^�5ҽ��(��V�/I r1��������q�P1���.[���$J��i>�eR�35��@Ȫ���4�C1����n"[�v�!�PU�2��UkJ�)H�����	l
޾Ҫ��L���iu��������,�{HQ��1^o$�9���;$;�U����^��%7 �Gq[���b:'������13G���&3�oEO�K 1q�u!����e��|V�ǆ�^<���\�Q�v�%��UvF�",���!��t��3��JШ��W����z;�[��ŀD���F̼$s{@6 /����d�>g'D��oш>+6�rPK�cY��:�����m���Pi(�|�FfV��H�F��M���|��r��Jln�ℎ�$!洞��� �<7�Y�Z����g�r���:e��AOs��+j%m�pY���ol흲��e4�Af��&W���f�����L�/Nk���t��@[�����>-�r���M�5yt�r�92~���c |Tf�kR+5T������}m-g��?�̮5�ĭE���W]�#���7`��I-�H�����4��hѲ��|���5������m��lB~=�&I�(�>�`8�d���i6c��!�<<�+�,p$�cύ��*�(#=-����|�Zz�*�����?�-�D.�ݻ{.��f/�\]68��~'G��	LM�	��[>�����F׻
��0@���
���G�Mz�$�Έ�μ��s�M2�8I`���N�~��a���X��-D�� w�b�F���㙀z�誳QOQ���Q���b_epM�µb/�I� gO�t�x �`����o0	Y���&v��L�����^iL�.?�SW`g��Z�I�ݞn�j�����s��n�x��K8��Y˪�ط�Iǚ�R�����6�zn�z{�n�:>��u�z����\^X2\JW���:�.�#�rD�в���28���ϧ,���z Q��ܘ^��5'�O�!_���p���W��k�����i<g�a�w��!W���E�&B��-h�l���Wpæ�8�I �4'�A|�N�����,�N��~�M���T��b�7D�gy�]OP������a��ܭ2Be��;fǞ_!����ɀ��'� ���Je��;��Ԭ\���0x{���r�����/��O����i��϶k��7vצg*�`CaΊ�姵Ŷ�T�LږN����	Ax��B�Yȅ���I�bN�;��"W�5����xEw��7T'@��,���o&#��F��/�݄����rw��TMoaSҪ�̙Js�:?���]aY�0%�F+����
2�u;z���#�^U��|�7R�e�Ht�Z��#��~b�̑�����LZ߶�e�x�13��ͷۀ�9_Q��O,��ZC��t�$Q[�"�\����q׀���������W������l�����z�oCˑ�5*A�b��u�iP�PR���[E( �Ml��m�.!��(Q�;)2a�G,� *��P~`���������A������˼��5�.���Ą7?UH�����tv�e�v"��/;�9O���u֎�B/����z�^��1�4Y<�2�����H�B��퇺7��.r