��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6�%�JbHZ�y�!�\�q�n��TB�}���M6��E�9��(�;L8�|^'ō���h���J���%��!b���Y ��p!ĸ�UmS�U�uf������A$�Ӵ&�{,�Eek痽&Ě5�4���e�"��J�sk��9�78A}��<��Z������'��{��!inHzVnҁ/	0��2a�f��w�3�����{�x)�zր�_��hP��z��@��5�GY�Ǎ8��ґ�����?�qL�7t(�k�ʛ֧L~�#s��Q��Dl�ÿ,��l?���IP�i����C�IqFD�R��9��=�p-?*��	P��j\�Ȳ��{�t�0��:����>r-x�:��m	�xw	��an��+ǲ�Vs�Qٯ�KH�~��em�1��C��oS�(��?�Ґf�U�L:s]1Bގ�|�!ZyF<.�`o��~�c9�p�Q�P#drNKq#�@Z�Hq�l�̑�d��c�n�͊&�V���G����9��8R7GAGj�^VrIv(p�J%��"m����:�>����s�3�-N�x���V�	�*�Z	�\�/��i��2�����'u@�r��靟Ng^�9�c�l�+���눿G]���}gnQ���t����"��|�'��'o���z���I�^�@�`2���i��|Γו��?%�X"0a
�(��/&h��[a,�*�Y!@3��Fj��
 Nj�|)�D)��?��H��^*nu�$�"��ZN�`>Is��<��*u�S3��U�xb0(�*�>�q��.��W�L�摒��2U��R��>�Q���i�
���I@��^���N�KN)�|��g]m��٨��R_zmr�uszMX�ظIK��d$�hG�2�<�ܺ0@�U����-O���*\�YJ�����F���>�|l�v&���;gZ�*�1��>	<`|}u\�S���!��u}��J� ��K	�+��!$/�����b�P��9uS��y�8?���jQ�fl�0��-I�j�� ���2����?��SJ-(��M�� �%�7o�$�N�ݤ�䒠
��bi?5<��svG���'W�ih�q?4��U:��%(�Ȁ�����z���ԙ���w�#$��&@��j���V�B.�=��E���<�:�{�l:�X�uz�R>8j(ß-(l�ٌ��פ�. �آ�������Q�v�����6��+ڡ&p�m���Q�<��s��1R	�nu�Οza�.ˎ�.��wtD���X'n\<�<�8U"�LF��c"z���x���N=�%�7�l����mS��K��Tq�x�2�X���.$�N�_֟�11��Ģ�v��	��1�6<>_���!����0�!�;~��rO�h��t�p�S�Z�����멓0C����#���"o\�)���o��Ϳz���cP�l,$��5�&��!7����M�#��q7�~�@io]#��S�-kug\����#� gMdM틔	ǥ�j�V{`�˶�f�>97���J���N�(&ln� �u��Ƭ]����h�C�L��1�� �^7U9XBk*f�!��n��>��g!�r��f�ĴpV�_���w��u=�\DP[�n���5Y
��N]�P�r2^R��� Fw3z� {�\o,jEo���z"��g8m["��
�t#�C�O����=��S] H5�a�`��X����S�|�J���.�T�ѓ��Ɇ�6�i�
 �P�&�s�0]���zv�ir��;X�4�d}�O.�� �""h���?Xnz�[79�Ot��)�~20X�ՌH�����¯e��Be��1�"����'p�Fe�)Ѹ��Z�US��f�f�Z����U�x��~��n�M��'05!9�Tn/Q�e�l�WV�Y�4����� ����;v8�8�ٿth�r���[\��AD��1'�2�[ﴗ��q<�Yr(,��u��:���Z���l�y���,�R/}�c)�o#�n-���<v�(�+�o��~�k9�M~ϲQ7�rU��Ko�#/;m��]��r��K��K'�)#9
̝�c�(1��X~���\=���H1(�w�"+��Z�����i���{ﺱ��ܫ\�!y���h?)[��©صģ{�T�fW��C�g�k'�w��R�I��ŭ�
���b��R�MP���i(Kv����,1�z9� =K=/ALʮ)Y� cS5M�����bL ,�҂������\"�ZNf�׍�{�Ս"f
�VK<�/+`������qޤ���0�����kռC�T!3(����3V�)�҃��g<�F3D8`Q;� �����[��9���]��zA��D�w�a)�X������=5���Z���-?<���:B��<Q����x����W�:~���H�n�W�rL.��Zq��W�����~�	�9r��GP�Uӹ���9���A�h� S.�B/��%n_ݏm(��WD��ۑv��8�;%�q���NAZ�d>^� ��H�}�L�'�2��Kd�����������FO���4iEL�?���o���_������_��c�Cd`�Yo2�����.X��mw۶�]ia��M�+����9M��i��T�h<=�Ye�k٘8��s���[~��2��¬������Ûy�aЦ��>*�?4�nzz3�`�g��O��P���2rzD���t{ϥ4��cfc����ʁS���hg7z��(N���ʤKC�����HG��<�-'��S�_#sg�I�V�}D&��W�]�%awr#���'w���v����ł�>��@@�86��$�e@��k����`�U�M�L�~S���H�%�a.��9���LV
IH=\?�rH��x/��hm�Յ�����K=���N���bG��'�l�'�e�I�:d	]���S��I����aE��uI-����7�?~�w�u����A噪G�,��A0���-��B��DFE��LuB��47$3P�R`�+՗,�"����=�<���X[t!�"��Q��h�12P3��;������+`��*wË0p��#���w�\d5��0��HtiB~��$��n��hw��L�R��/������bk{ED�r�ӗ�nmv��o1�c�{e��à\�������atϖNF��C�N�C�S��L���UEVc���JNt�G��y�����\�����$򐤾S!��B�q���j��&r1��� ȕ�G_���'�,C΀o�#w�u7���Ο1���g3q�I�%J�I�U���7���)�i9y1�22~����Q�s�E3,fM���(�֔	��Zi¦���6��}k��W��4b �1��Z�]e� 
��H}�O���s)ĶxY�����1��#�#p�]-,�k �ǘG
>�c>h�Ί�����0����'�������=�/+��ܙ�BY����{�M�BЖ*���_} �i���nyZxOPv��g�R����V!d9��<)R"tn�T�7�UMV�|��Ý��3v�w�v��S�D~Mw=kST:Z+,@�6j����,	�i��Y�ݎ%+��̏o_כ����?bId���	�!�B�=P&�7�E�f�٫���H�5�$�~�LϬ&i�����"�_-mZ�de�&���U��&z�U��'�$�1{AGx���ƨ[P�YX���	Tz@x	�+V>�F������zT�"�3�>(��MZ�+/e�0��eF�ܟ'�b�#�M���HF&��\
�)�B��K	l�{i�>ڴQ>��}󒳖UnA���e"�jO��l[�v�̕��[ݐ�eJ��rx����z�TH�Nè�_l,a� �k@�'�%-@p}ޖ��,����w�6|���3_��a�at!����ܩ@�_]U�bX��X8���BE��:�w( �6C`������6��v}���++� h9�Ձ�$S%H��AՐ�}o��_x�L�9��N�71X|-�w�w�o��S^"����?M�c��[�l	x�W}~���?V"�`��=I\�C�=�E�POdEξP�>�J�y����:�BT��u���d�\�J�JP}b	l"�C�,~���;��m�_2�%��wdFX�'�AV5�wvW��l(��.n+36nn�2�j�z���-ɶ�~A�"�f��U�����(�S�ҕwnB��f�6+�
����긒\3#c�=k�=��T ��ԧ���R/$�߷��3l�n�c�sP��N�����]nʯ�<:=�P�C�\�@�����W��b�qs�\:n���؝A#�߫�����xCMH��Ĉ�u��魣�z����zױ��$v���s�x�w�,���1穨!aGS��\�C6����ͻ�r���	@h퓛[�Ŕԩ������*�0���F��J�ܙ���fue��O�N�ۑ0�*��|�?����4�����oA2�Lwߩ�'$ �Vz��?�,�e�����#�8��N�B�Φ�����\�,N&2�ȵH{%~�b��`�di���x��jJ����t���-�[J|k�(����lT,�PD	������ ��o�{�|�Y]v���D%]n���%P��w�ge3J ���5%ӷ,~��c%���}��p������آ�� ��>T1^CP���gN�]P��z2s%RvP��d�n���"mfY����[�r�DE�Ϛ��K�U���ፃ��oߎ����x2�)f1�����Z��,ӯ
��Z<`(U��_�~�D1���dUj�PAM��垿����~��Y��_�>��O �1����F��ԣ�x���b��W���&�o�����|��/�r���>�N�:���S�y���'F>�@�J��-7{􊇕vp��҄��)��$�3b~�Sj�m�;3%��v+�J����ϥ*��I���0����<۹'G�)~��ʚ|m�'�pY������C>rDȊ�T��kX��|���d��
�6Ȱ1L����_vS�1"��F����פH�?��橷�������Am�ɨ�k�#ª�κ�(>���Z)����������v�F���rw�~�[.�L�	}��,����_�,���L�=����r[~h�}ʳ�^9w6�6$
�G�."42v��//���z��6Y�6�T�%Χ��"��������竚=��<�3k�e��43���X -�Sୗ�Ჸn@�.���gP�E�t�O%?"l�6�X����U�俷����������MǬ�;  �����g�'*���I<9o&�1H��~ #.��"4�Ϛ��b��W�iY�bKT��*���ГCO���b�SO~�`��.\�B�e�s�2D��J"�-�X[NuXY~������x�!�)v�N��Pf�D �/�:̳҇z�����t#���i��,ȝ����ĂT|�*�� ��P����1|lm�ɶ� KH�o��$�> �G>�]Y��k��R���@?k���J�*�^놯<e�+F�'>3,Fֆg���-��^d���@�v:S�"�Z�`V�8,�s�t��{tb�= V\s�;%�V*iuT-NF��B0�����z�}���mY��ķ*A�����v�0 W��w���nVc✾���� �ٴ��hi��I䮡m�3�sm��=��N�93 ���SO�*Aʚ*�����@��jta�W�P%3��(Ƶ�z"�G�^��4�k��A��*m�Ұ�!�C2[]�Gn�Vz<��Ima/�����$}���齄Bm��}�|�pN�����&	����T�>D#y}f��YghW��p~1H&�꼆�ˎC^|�ۼ��
c-`$��&���_���4�$���|a�x��Z����h<er{8:!����]������)�g�1}�3�3/E:ی�=��>��4Θ�\���@\5�����:��� (������!�YF��0r��H�]
`*`�����+��j{�F�/�L�B3����C{�R�.�ly!Z��½ښ��_8E��MШ�����~�LT�w~��v���9vY���E����:1�w�	s��k�����Ɨ��&iNA����9`	�GP͗���{���d�����ed=�|���PK�g�I����]u<�MZ���.���I4���g��H;��r�#q�S\/�v��'�Ng.ဖ�wv� Q�a�ī���r�R:N|j��e� �����5�l|�����"��T��_4�.�.5>z,�do'p�w��Y�6wX���H�mxQU��ѱ�7�>����Av� ܭC��=��j����?_My?���"� ͘���(1���(w	�j��1�3�"¦7�a��2-!n�TN��Ǿ� �бfY����7����w��'�4���K|�v��n���!��ؠWT��MŦ�`o�I�H��Z�<��M��(��B5_�xU���2�e��/-=���{F��>pY�T�l��o�<�1leJ�,u�P�o���Ţ_��<���']�˶9������Kf~��m������A�DG�-?�Wh�Kt
��a��U���]l�u��Oq� ,�bԖa(���|kXuT�{~���M��*��ec�5�S��h!���e��{�i����@Z;	$�+b�d�`qt.q0�-�P�� ����c�������ߛb���<НƧ�uǫ��-V���1���+j���$E�����M�{���`�k�3���B���#����?�k����J�`r����9��� W�yz`���2�Js��(\������k�	�+g�.o�,���(�no�n�o��0e[D�@r(�V��#��m���`��[�HLR�Ҭh�-�;�#��E��ׯ������/�\B��93�u0�u:���(�I�Bƺ*�MF�y�NU�<��Ǹ�1ERK�n��al���Zh�nؕAOl���}-�'�@1�VU�����`��f���^ފ�a�*g��{Y �q���5���}G��،�$z��>a�k*�_P}�3:s��x�X��s��Z�@��V?ɓ�S
fo�����wZ�c)>��v��Z�1s�DE�!�8���x}0N
��g-(/U��fS !���3C C�����ܞ�akTN�A"�pgq�ѫ}O|<�yn��%7:R��x��!������-����t��`���ID���g��R������}�p�O�ТxɌ�2��`�����v%�sN+���ANz����8=�Rv�^���X�q�e2��� S'��6J��r߇h�w9E���e6�?�9�\�*���ϡ%�@�4m�P��y��q�:��W>�A����8�Y�d�����/��/���r�$�f�� P�P�"�mզ^pu�J����58�%J��M�}�2�_�|o��u�D��`ZGC�'2��x�%�A�_�ᅱ��v�#Ө�Jv���3���HF��¯�Oa����J��5�DEGa4�`�?��O��jhѐ*Uv��;��f��}��ǌ�ש���ܝ�*|kBz/]2I�z7�5z
砐"�md���}���~�3s��N�BI��ꘓ"��@�?��\P��:���z�b��6d�:�_i�j?��}=h�������>�l@�a�}"8z���mݐ�oq�⡝�#bA�X/h�n�=��/�_~?�x��,���&l����*����$`�08V�|M���h�GS�A�e3�+�A5-�7���ST��B�M��搊nC����!{~%��Uh�MW8ʁ������rF�㐌�7�й2�����us�F�~yYY=�
c�����5*b��UhΌ�[�L�D�&�;�D-)hY��� 4�-ŔHW-��:{Y#�k�*��0��up�(*yD�Yհ����ӥ+ >�#����g��~?Sgh<Ę�p�9a�(�i��6���ӓ� Y�^6��۪J37=���abZ|�<��ʣ����r�.Cg*4jiZ��I�h>o������5��f�G6��d��k�u�?�	�~�X��*�B���h�wK���Abva�t��L�31NI��e$�k�b��#G9y�K�c�JYeð�����1_��C�eK�;��]��Fʷ�u��-��b��"�a5p5�D�x���:0��h(�NF���ߛE;����.�6�q��;��e�tB�7��s�dB�;��av�n�-8K� D�V[�^ͻ �����%�M �i�OХ%�G�2d��m
��O�
�F7�{�6�9%�����%��f��	�{�g@�yBAދ������;��,T�[Zg9/nv�xnX�ٹ*�b��=�.q�^1��ת��.���; ��<r�j�	ZW}
i�����t@�3N0A�!��w@�7�	$�VzhW�|Q�D�n���{��� &�*�4�l��t��5�G�&��W?��4H�`�|���������M�SQ�(|0W񍱋��!�8 ޸������V"ā��h�S�EY�B� r�Ê�Tka	fI�~�OIu	l�W����M�p���"4��
t]a���,�	Qk��U$
ma�:�G�Ul��u�P���Z�e��q��yha5�
����DY��%���<w=�zh�&�k�˥ɥ�'09�x�K�«���q�oX�OE7^��󰨖�@��~��� ��oc��X�����X���N�o���>\����e�R�����"c��+��,��0>]��<��yk��C�7�"1t6e���S�h�ʆ����8�����7�R�u�N-�K^�����;O>�����pb=��g��Z�{�CL?z9j��c8)8�f�Hg]Z� ��4.3m�c��xRJ6�βy�g�~����g��;^��Y ����׀�nf�HH����6�LR�)k0c�_��W����+|m�������n��Y�:���<�5�Y|��+	��^�Vb�4�l�L�u/��E>��V>�ch�/8�U�e?��Iq����C���0.p�8�![��pۜ���!�jOp4Q��/��nD��ɉ�4"e���sb��G�ɋ�M���49�b�Xg�`��'�~�p�$`�u5�}Z�>㝏�k
[=˂�g<��Z����#��ԡ.�EǞV�?8�vL�/����~{1�L��IR�����c�+����+!�s�R�@�ތ�|�/�?x�i���#�t>�������E���ԝ��cu��?�D�z��c8�>�[,�s%��PN�Eo��?�<9��z\�b���=��m��Y�Ɖ����A5Ʈ.{g'�D�A����f�@�պ���W[~}ٌ^��%a.ze�^~/2D���;���� y\��p.(ytS���9-(
ٴ@��ų��okD[��T��w�~gݗq�Fw`�I9��5�i��:�ӁQa�Sܙ�Y9�ʒ�+8B�h�G�a�>� �|�,���'�u�
T�;�� ��MW�D������d�h"c�3���+��o���v噎1�X��'7�(�L���{	O���V�t�}FJy\�1k
!{��}cp}�7vU��1�C^��V��]K�E'��X�I�����X�|K�1�����N3ٛ�J����YA��v'�@��^��W�)�vs��6*���� F��q����u>�U�[���(s�� ���J��d���r�����_������\�um��3�e7�4�A�p��wdݮ��;�\Љa�1\V/^��0��;�䰳���E����0n����CPa��
�^�Ef	�u�K�Rs9��9X�=Z��zx$���E�񷗗c�<�?��%�:������v��:�
i%�	�W+y��/�̝�EQ���W�c?�{����m'�ߧ<NA"3)�
!qn���{��0��¼��f��J����lǰ+O4#M��i�4��r�¹_��õ�+HLJ:}�lO�/��^�F�͖<Ra;B���*��K��ь
_�L�6s��:�%�`瓻�ث�״�[�ϋJ �.C��y��_����"����q�'�<wėY�/=7)�1�P<��Z�:{��{��(��,=���ho��A�� �r��~V���7�n����H�j4DҔ#�\�[a��k����R��;�j�#�26��_e:�#�T�_���M[���[rv�s�_��! d�o��>�R6b�3ߕ����1��� Nr"�Ǥ��M��4��)���?�(U����%�CoO�`k[�绕��m�G�����И�׬(q���~g$C�5��cၽB�Z�!q/Q����|э�Ze������O�$IB�}�'I�5GEzmx�K#��J<Gb��d'����1J��$�	⯏U�9�3f;����)$-����uD�U���h^�����	��;{��N�K�݄x�7a�a���`?'�T�:Q
�l��� $�P-�A�P^o����Oa� Bn����ۖ���,��E��X��(��C�Ǐ�-Q<m�F���:�F[AΌy�λԄ-��Rjw�r@���}V�!�b,��vP�p8��e�-Ο�e���\�Hă��w[�(���>?!�48d���6C1��������Sg��r��GvC8#�����R����f�4�� �=�o�x��hՏd�k��H�)b�PN�`l����H���e��D�swݢ�-!{�M�#H�My6$��?#Q[��%ϵ��I�r|Q՚�:@��L7��.�%�c�*���+"_p��m犦G��T>����
�r�k[�^��j˾��`���#���&26�Q�B���s�Nj�J3Y:��I)�ޯ��P�w��嗋�{�l��$p�.�`��R�s��̃���O*jY�p����W\�_ �����ОC�[�wg�(6lDʩ�1*�<?�$� �c�݀���R�@r�Ee����!� �I؃�\�S�a��zu��@��kP)���Kv���T
�����x�Hx��7��%���=%qv:{Q���;�-�c�Y�b���������m���'���*!8sLΛ/#w'/ �)��b��5���n������Sv��dXw{�����	q[�2LE,p�h렝fgU���W�A��,h���mMH5-9cs�,[���W��oD����<�ˀ�gIQ#	,}�U��O�IN��1wo'�h�"���׽�ql�H�Kl�YKѷ� ����$�|�!m�!��J��C/ճ�cc0�"��J�$T:��_����L<
��?F���K-q=��
炊�F�9�*?N|�oy,� �LPuާUޑÜǯ�Tw�Z������u�N��)�g�%�S[$˳��t����%���Ч���IN@H�ߟ�2f�0��b5��=�ọS�4#M�[#�9�hS����Bơ*t�]��[�~�J2�Zt��
4�J߹FY��Y�=0\t���\��-��_�=���}�Z �6}8�>�^?\�
��{��N�?�T��S=�nZ�5G�t���}�"�}��f��X^� \�E-� &H�y��1eP���熓��������6E|,�\�p:�Z��}|�I���JF�N�c��A�����\@9���m#ؘv5ێs��Ĉ�Y�C%FUq	�nW�,n�UpD�s�"�c� ���;*����r2���d��E�Z���K� ����<I�Y�h���2�o��"����
1@�Ou��i�2�Z��>��!���D2YF��� @O�Ż9� �2�6wu����4'fF��%��k\:���||�r�J<��!�J�������D�u?�q�0A��Z�
�k���U��)ԥ�]�����}����?���~z�}O��uc��4?=)�"+�#�GR�O`x0&r��1�<�o��k���|�4j���o�
t,����oH����0GW������냂h��s����Su,���K���.�f>0��g*��vkR@���g�6�g��w��߭�e���>,�_1/՞. �q�3�_(� ,&O��	���Ju6��7ӣ���NI�O��LA�>�D�TD���Ų!��n>4���������,���ʥl2�W͸W������?y\�W�W���E����kY�c�*I�,�g8ߘ\
k��G[� � ���W~g���j	��B��s`���-'2|�sN��VD�� /����t���54�r��<��8@a���{�Yު$��kڍT�J���n�W���`jo�p��Op�nng�����*���V��J�v	��o�z{s;�J�QK �Y@[��]��Bu��ԣ�8�w��U��jv�R��u��v=��-jI.�[�(V*N���M��?���F���)�1OI�lXVQ�$UᱴM*��Gw��jU@�����J��L�W�4��3���S/�	�yj1wI'׽�7vi����t��.�H��}>����֘�=�*�'d�j��,�Xȋ@=o����sO����� ��g����e(���#mJ����L�	�Ԗ&�� �J{�:�� ��[�Y&�h��޶������"�A3ŅQB����pJC�=��;��
3'����6��r��洔,���r�m� N�Ii"˗R�Ӯ�V�f�C(��Ν@�R�L�������ꜜ�����˙������R<%��c`}���1�9���Ju<�B��2�"]��GA���E�^gb�9k��AAUOv�ե�w	P�T^W��	W�P��w;��^TAN.�t��YO��