��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6�ݐ�௸U�@�ëA�L~�.{-�c{A�nC�<7F4t�R�cTd �]=t�I�C=1:�b�A{8�B!"�i�X��R���r������&�2�=���o���Ѣ��,I��:�D �������u��� �A��|��d[J�K�l_[���q0Y�A��O\��z�����y�dc	ٚP� C5((�Gx�}#?}↷?\;�C����t�P��	2,�I}J`mv��l2�@�D��!%��x."�s��U��8��A��T�m��ׁ���r����M��=���J���8G3QT6U�**�IM������1�~�����������< �����
�EC8�bX��53g{�� -�����%�XQ���w4-��Y�04a�C�.<{����4���F]C��IL��=�?�n��zQ�Z�@W�`�2eo����>�z)�	\+��\��0�������d4�R���������	��K滁��~�}�?�i�63��??�T�0SG�Ac�M7�"<|�H%'q���sI�}���Hd��Z���k��"����{��}4�z�776r8[�(�k���<����
|S��#��MOF�D碫d�t;�I���x�#,>��3����Z�#��$�b-W��n���ټ�MTf��[��rD�s�#�xz�����D	���%ׇ$G�`i�������\���qg�W�����GR%g�����8��������n���&��]L"n<�f������qݘ��E��fY�QL���8��X��ERex���;;�o�(��|��sU<ö�^�Ѻ�M+ �����k�ϥpm(��Щ����5j�I�+��'�'틄j<mw�M��w��k�҂��%fG�6`�W�WUr����*F{fڟ���;2Q8��x��Ǌՙ�(�q��Wq��Ü��$��UA�s�i��0=1zI�Џ{�|����3��Vy�jR�zC]��ER����{gf��4��Y��)��q1$E���Hxl�e�N;���'�M�J�8�F*�J��⋶~g�r��s��M�@���-��1��v��\M&�E3;���S��G�rm����ճ�e&��O���ڜ�U�NT��r3��vO��`q3�a������p�ef�m$�o�s�Y��t6�ԛ����B��֋*���%\���i0N8zBԑ��x>g��`�GFҪU��-�o�l<h���d"0�H{���	$�f�qGDa>8��b�"n!Db��dIv�똌��<j�\㫏������?s��6l$��(H����9�����E�'������ ӑ�v��l'��͂�c�u�V	����F��:u�i2�E�Ya�\�t	e��\��A
ކ�*�����̿p��mI�90)�鲩���w?iǣl�f�o�*7p�z�c�:]�U�h���Vڃ�w������TU-)O��>,�Q_)�jO/Vׇb�z�.��Ѯ޴����^_081n���k�nn�0f�;Q�����7Nq0S0(U��!2u��uS��:~hPÈO��t��'R��
}�5����n�Y2!�k��q:0cg�C;�5Qۀ�n���H��ܐ�C���Kr��TI��iOL8{�����o�\�$�Ǿ��>6R)+�T����r���Iv�p�-���
��.̉f�R�#�h�~X�?[�X�}��ԡ\�HA��U�l5Q� � �K�vc_�.^���1��π��<�����Q��'�nB���k�MX���Q��f���W���n9��8|��Nd(mȈMf��a*p��g�����'����2W���m	����F�{M�%+d}�͍4�[���PVk�0*�fI��Q4��|�f�S <}���6
��QפI��b���q�&z(���:9D�4yš�j+�Sj��Y��]t��]ԗ*U�4x��������ܺ�r�gt|�#�WY�%�N]nWY�`���(#L�-x�����mFR��u(y�-���u���|��]N����ڝ� ^�(��A�E'"a�&�d��)đzSsTM�`��ژ'�� ���ɜ}��r<��e��_��(p��X��Fa2�d�Ò����b�EY̖_LW5g+��%\�E��h��>4�A=B,�]k9�aV���ءqՂ�$O~Q��PfT��
�>��@ �Q�ۢk=���ƾ��#��L�@��;"�i(@�6��G&��ؑ�$w*eE�{t]�p_�I��/���e��>õ��f32��ڱ��B�cL�g��x|@Ь���o��3�G�Ǉ���v�@1�',�8�/�m}�$�P�k��?1l��,\3���6��Ъ�whK[A,�-��I�����`��	�t�I���H���CFbK^le�a�B飩f%�d��Q���`s��YD)��sY߆���/�wn� ���Z��Z�I�W0X�Ŗ���:�������6���D�Dg�����ON�!����� ���1����Vc�2$��,��{���S�mGּ��ٝC��8tw=b�D_]�|�)X�. �|_�O�~)�t;�5�y8����{�"d��}�ܪ2Auw4�ޅ
_��C��TzDÔQV_:e�t]�q����!�.�`��"�?���� o�wU����������ʹ(�h�j�0���ս 㟭����S�и1��s���*�!K�U^)�=n��U<�udT�2�д��-�(z G�e��oO�]/$�f�QIk�o�%�q�F�A�KČ���a d�+k�ѣg8FY1�n�v[�}�)s�Zp�ư玏X�nv� �W �����;�r��Z���,���,�.����}]=v	��-��+�֓Jm,�/����f=:��T�x1{W�&=�W�4{���]g8P���k7՞�(�,ul�����
Q�-����y�&�S��B�9�J�+��3�v��<��&�(@���SF犾,��[`���E"�X!����\�I��y�����|?llL+�Ïnh�I��ŵ��|H)5��'�GX��@��PS��*�:�@��_��)�o�A����KS����z�z|/�_�'z��l��
k��wz��
���S �9�H;5�>6�ݯEOMC�K*ە	i�ZUr�����f�d	7�n�^�
��'b֤�����O�[�<�4l$�{bI�O����%���M�FO��Ň��V��t�L�ܥl�������3�t='�.g�I����8�Ut�l'�vF�&�Ŵ|pQBcx�.2RT�zI�/����	�6�����[ݸ�`�1�}�������j.�а�����IϹ-�@��B�<3�6��n�8�}����T���ګ7����w�����N����*� ��_Z�-?2��k�_ؠo�@%)PdQ�[���H��$�{{�̚��`�����32<�B6P��e�v����Qz�NN}h� �˔$ b���U軣���(�qy�>);���D�5������&�r�����ƌ7�:�C�(���J�OҖ|!�@�$�[�!=�R`�d��_̷�g��#�m��v�X�%J1���p��I�&��m���٫c�( �%nn[\��  �x��HF8
��������^�#�d�1�>�m�.��bM��Hl[�פ �:�b#�E�$�m�cs�R�^j�5+R�\��e*���a�v��T��ۊ��K�+t��`bL#81��	�7�ҳ����8=k��[z�R�c��!fbP�zXL[���^�"%�	�ub���!t�e�]��=j-�4���MW*�M��b���U��Y?�ԡ�1|�T���[���7׽�c��%�P���n��1�T��,��52 �u1�AV��[�����d����jH*U�\��U3Y�����@���[�ZA/c}�~�3���d�8�l*���\Վ'"�P}�)B�{�#a�G�����3Q�B/�.�����1u����	w�d���߃��>�.���3��xA�6ԶSxx�F%�C���V�Z�Mfz�)���R��ua��[U8.U5#�^u=坑1�}��� ��Q�T������X�k	�DG0T�K��ؒ�	(O�R�W�#���,�t��d�b�{Ȅ"N�$��(�>�����U>H��E�0&7h����VI��Ի���^�d������|�~+o���:RF��Z��9Z"r��& Wx)�����u��/�Yd�t�؀�!:�iH������_��7]+&�vl����]�R��:��@��/2���L�á�+o��ǩ뾱��,���U5��v^�.�s}�Ý���Gl��НO��>{�ўa���"�2C��ʌ�̏{�VI]U6���� G����e+z�inO�i�^����}�v������VH܏뎻���$�ڔʶ�׾�(J+i������?^��7��&@R�~t�H�ج�V$�_�wXM��.L�HRpLh5��S'p�Δ �in��j�rpD �K���6���.y����jt��`���d�T p�n�J��3��\�R�������(?��\L��P5��ϣ�Z�~K�¾��5�BlzO��P�`����'�K'��M�	R�V0�����@3�I� 3o��� S.k���#D��G/��x4h6^����0J����p���Zg��C�Uӿӳnkן��[LM��i/�eB���h�Uf�����	����)�I���w�����X�^^�v�׃���7��-�:���F�K��p$�Z��~d�VZ�M%#&?��gD����`��zم�l����C�^̡߸ɭ���8_'q:���Ń��SQzJ�ƶG�I=�ęX�IF2����B��ZΈJ~{Y8U��%��u�38��-(���=*�ⓘ��|vn�A�8@�i`X^�r=
�OIt"���9�LF�?i��'�%|��F�*.�#F)4�����eyL3;²���lPݚ9OQ�\�F1s��E�A��*rw�D~T.ק \$��
��x����<Y�g$\#;�E���V�l�'���.�y�L�5�ե�{�DM��n�ΐTz����N�D+j$�*����-m��8�=�"���$���ମ��>����"	��\Xkdۘ�kT�FJ1��\�ľ�O��yYy_���L��]?+�)rٖ��Svf�K$�#Tu���À��!f�aU�g�>��Q�uQ�h,V��ٍ��AT��eB�{&�w?��)@7؄ʯ�٧�����խ���i��ϝK��♹�SV��hԴ��U��g?�9��K�&��Er��%�da�Pv��0Sy����#��L�c��#���W�m�������$�T8�X�a�5%������e�8J��~x6m��r���;�,{o̡���*@N� h����}�5�ځ9
Hn�*�_P87��;"������P�s D��ø��4��W�T���c�7X�f�.# ɏ������}~."��E �m4M lo�����'�s0)y'i �}Ɋ��L�V.�r���=�z-�/B'��a��G����~�pM�#��'�b3a���hD�~�����f����6��[�P��D+�,�$Hq�C~>bi�e)P���z)�} �uo�S:��)�����n�]1>������ e�j)��EP��*��v�l�E�Ð��0�,S����&^�o���-�I��Xh��N���S��ӻ/w�r./#qeДg�"�F��?��"�������GeӼ���K�z�N#6M%�Q��$+�5k��6�_����▫�f�_H7>26�X�6ZS�LT�YR\R���5���z{�C������ѩ�ed?X#����B!
�^�%]r.�ˑ��:o~�)¥?�p����� Q^2�_v�^�~��Bd(�Y��p����I�π��,h����+�Ě��(��A�_����J�ME���;�����q�� ��̤�)��˅Ŭl�l�f���ܼ��@pB��:��O�/烻y�F�ƽf��t �5��Ɉ�?Ee��o��6���0�̘��T���zb�E_�w�n�pר��Y%��X�ȓާp!]��R��F�=,�y����oD�~u����[o�$�1,J����c�B�T�	1��,Ѱ��[vLʵ<�&BV�7@�'$z2�L��|�	V˚���{$s
cng�#8%$�#���EJ�02�iZ�ǌ�,*��ov�i���+ޕc�ܚ�-@a�q�Q�T1��D��A)����1b�h�I(���נ�*C(��&�9��N��,����Z�E�=�6�ny��ʪ���7THb��y�o3+�Yㆰ��Z�4����X�O-?�3���a�L��É$�-��R�>�$�I\�h'�U���u"��C�S��NS��}��m���~98B��g��r��ڧg��4+����myC�Vq�-����>��{K�±T�]^nߛC4�����ug�f\�#�T��o>�2�j��;�ѣ�����{�]M"���.C,��)�ى��'���`⛙�D�oi~q�Ү'o�F�_��������ō>���Mv�x�!�W[�\
2:�F��9�/u���c>�y����,�3U>�E�~����g* �E�ϣ{�ь�B�9�����{3��j���ex-�O�=[���qz,��&I`����)��a�w�e��WM���W�+:k��F�!֘lI��a��W���'�����{ESG�;��w|}���3��.������P�|���$b��-�
NK3"�ۅ3�e1�ƶyĩ���+Z�vl �M��9��i�>�L�!�Y,�a�.��A�G KǼs�#b������&-�渶`�2�2�͹���k�9��g�C����!�F�j�[��<�C���&�r.VIn�z� M�
^[�"=ǌ��yT~�ز�6 �J���b(��c�28�2�Q�o����G�p�MOO�%.�X�'^����i����lԁ0�;I�.�b|1��K�=���tu셹sy�C��"�~ֱ�kzE�]Ē!������z),�"^�l ��{R�����F�r�� I�����rro�7��M������6����o�x�����ar<���I<f�)�y��M8b�H1�U�`�+�`�K��Y-�R9��:D�'��2�Ȕ{=/k;7l�I1!"*,0i���[�?`�/��9^A�0��̈́guޕ��pm�Ht.���M`���B�@N/wE�NvÌ92t*�,,��u8�ڔ8��N0��$��Ӕ����|e]	y@rO�tH����3]�]��&������t�a�9�8�j�a�"�H㐻�Q�&����Y}�~�o0�>d����b8/Z����N��Ӏ@ZhS���W��*�������!���i�����q6�B��-���0����eA\��66X:�!R'yL=����Nb���Ψ.Lʆ�cq����)ڡ��Z,�"X�ZP:D2S
"��F��G���H����I�=e?�heb�r�I{]�X�ЏtVyC�'����X�R���t�R!	iI��,֞��m(�MY�H�;=q[�e}�1���v���M鳹�4��݄Q�+��D#�L$���;�lz��߃1���N҇������$seQ��;�Y K���{�f���� xz�|d���t3���7�3���?Y{kC+H�j��!�`}�f��t6��(Ê����%2�KZ7*�h�C�;��{R*�>�eO�H��f�0��h���|�Y���@�K�zm_�Q��Uu8��%�� ������n�gi��;@�1�>�ԑ��E�N�IƂ�O�6�N�1q$&�UƔ��ũ���[��b��G�`��*��{I܃�c
�x��ܪ�'��칲ZT'?q��!����xhK�Η�ir9I�3mTo�RxG!��(O�lykݦ��p���N
��ї7�1��N#�!��4Ӱ. ��2T�)E1��ϻO�Pr�*p�|^d�.~i����d�i��7#ɐ�P��k����L��?Ӽ�1E	$*΅�%�\`�8Ӑ������v9�D�d~o�����<ڈ���2$��{U���3����p��
1SZ�
���{V��\����h�sr�Py�TezU�jH.�w�~YV�۵7n�Y
�x!��H�,춖0�vd|��E��&Mz�7hq�6Gd&��̬�o0L�����dJ�"R��}L�7�	ڼZ�w/H��,A�P�F�+�Ș�~�71��|�o4(���kg�u�s�8sN�q�_Mɾg��Ǉ��� ��ۅ��'�p���h{�z	��� u2H��l,zZ�O\�vH�������)��J��u��ZǊ����PIWQ����E��4bΥl�������ᷙZ��U]	���6Zw]���}J�(S��3w��~���!���z�*�ŝ��?h�0�u�p}��(t)���c9�q�!���K��GF�?M8˝>��+�X�f��?6eTd����M��e"��i�~�_i����ug�_�m����yD�>A�9�xr����7��(}=M���H;>h[}mM[?��h�� (��r�4��^3�<3<;���F]��u���$Z9�`�<�Q�E��kX?�U�!1	2΁�8+~
m_�H���������d�P~�/�s�ǆ[5ɔ���t`�\Ej-�y���/�jө�mת�͊�2�Xy-�-�L���K�St\�sMܜ(_�V�ʉ��y]�R��IO�
7�1�D��;��T������r�S2�m�8�*�?�5�ڣIߦ����fq����ύ�}e�.@˓��N�l鳪~1;I2�M}Z��o��J�Q8)r?���U�w?�c�a�r��v� h�{y8+5'�����"K
���Lt�z�m�LN
��g�e�X��u|԰@X٬!���ķ�H6N�k�����G%���9z�Drm8%�5����˃�|��dkT5p����E��k�8<IA b��&��X�<�g�܍�ث�x2u_	��5�CM�+�'�u^�2N���	(���l�_��Ʊ%g @�͈���Έ ��?�#���HTdW�&d�,p,�e�Z䲸8��f;S��#-���8A��8������c�M�sq��0 ��UU����}�rcGk���Ԡ�n�*�K	�P���� �N��	\1lK�i��#����Dz�P������i����yU3#�&;�7i਺Ci�b���)GE��{?^с7�eV���B$J�5/X��纪�U��&z�u�2��9��5M�ϒ�� ~�o ޅF���[p>&��wM���
 k;��i���^�IGͺa�0p�	Z�uZ��ڙ�W�61\�Iݼf�rW$EZZ�{�/W�����BeW��sX�!:�#k��
/I���.t I���p��=����Մ_H�!���=��蟒�s^�<��4�,�����P���%D\BaU��'�MO	]՝����ӽ��|�ƅ&|��.�焰ö����ч#�WYzZ��,��ۣ�w��ꅩ���1k�J�[�G�̚Â�W��J5�y7Z�����\�a�KQq�A�c@K`�vn<���jҜ��d���,�oV%�}�e�J����,�=I�ο��5&4�ݘ��F��r��:��I%�nuo�(6���/�Dد�q~�F��Q���Kr�nM�����],By?�64���ѳ>�Ȗv� �����,���=YƊ����Kўӧ���.+�CzX�Iü~݃犈�n�٬�Ѕ�D����%��y}����,�T#e%�z�G'�_�p�D�Wlk������q
�F`n�.Va�<���-�ϙ������9ʿP{I)�04k���	���bLX�S�`�b粺R����=��L<>��ʚ���^�Mr�Zl��<X���V`�`^�pK��u�ǌm�����>mv<���w�d����8V�,���"%\��ų��#�p�{Lwf?�<�%[1`m��6R^�?����f��^> )�h��TM��m�I��M�?��Ky_�LOPm����A )X�nh�J�.�y�|��*��>�����'�/��sc�Z�h\]8��rd-˸H)>2} ���A�R^H�9ꦌ�G���B<��w�Hk#�E��<��l��8�?����h��Uz���u����J�~�y�ݰ;H�ۑ#�]:abw�>�d���~l0�C ����o��81��[gA�̛i�+�\;�[�U�܄%�8ƴS���rJ�I./JZIb�>���S��`D�M#��Er�eΑK�]{/_R.q�q���&�nN�HPN\�q���ת����'�/n_�XB'��"�љ뜧�q`�8TWֶ�V"ҺI���a^���k&=�D�2��jLO�崕���k���6�����&�1Dj([�e��ͅ���)�t���A��F�N++M�pi%�����-"�iJ�5w��miw8�"_�)�st~��NO��c}�����Ys(~����K1��ϊ��Z�Y�]�6L��^�I�p���t��Q�qž���P��C�Wn;7�9�0�'E���B�xMPs���mW����L��cRi��RN5$Q��[�ir�嚛W����k�V�n��7ċ�-񭫫��Y�P@8�٢��ڕf?To���S���7�8���S���Q@����^��k�NZ���l�ĥ��O���T�hsyf�O�53G��ă���ʢ�/���gFvP<b��W�AZ���΅f_Q���@�Q�!�&�]79���®�#W�o��F�ŽPOZ	�E��j2Q;�$���8_j������T����V_�ד {��$�|B�"���)�5Ɋ����3������r>yMS�IZg��莅�Œ��茉���b���ͳ�����JU(A���>ih��N=�<�y�;��6gSf��Ȱ�
�y�\V��M�%�f��l�B�e}cse�H���W�ϰ�&ӆ�d�s�wF��u��)B%L>����kˉC�r)����"<Ty_��q-J���Q�w�9Ja7�(c���Y��+|
���_AQ`�t�����4�=?���8��Z:�M*��߂���RzT���)tዴ�9-���A�ؔ����SR�4�����&Ї� '�}V� �YhG����5A�J�����Y����p�g�� ֥���ؤS�8֟DE�%�!><\�`���qh����XP��?�2�3	��3W@��T��F��Y�&`E���*����̰�~��щ4��<{�迊m}��� 7�V�Ew$����Oh_�> .>����n�q��@�ʛ�$kk��k�ݽ0CMy���FZ0�He��R��p�ԏ��G�i�1`.b�2	��_�<�t����v�U֜@'㖬6V��
74�E�7�v!y\JŞHD��l�m
�'!Ν9)9�m��{�wA�<<^˅���c��;sU��=��*+|@���9jҽ�����3'�KJp �9����?�?���|�&Z��o=ä�.@�H��s)�|��	�rbZt��!�HI�����:)�jG�ƍ��V���S�繼)���$ڣW�{��@��NϐR���)ه��� }����ԾL��!�c�k�H�����@���ĕ�o�z�uN��� \b�,8�t���YY�`����ӻaKr��Oz��eh%k��h�8Z�b�>���
����^��P+�C��a��"/�����]���EQB�╌����?����d�����a,:狂d��a˩@!��������D0\����������;ܤ�x�i o�	���O���B�=�q�Ԉ2h#pRE#��n@�����8���z�� �͢'{�
������zb�˝�!�q-��&P�m�y/�`��~:�c�|Q��Q�B�iVzS������OA�5�Ӫg�>?B��q�|4�����M���//��-{S��6C���U��[���D��-��u���/�(��9`��GP�A�l�����`�Sҩ[��[5]�:'�E�� ����C��	�k8�Bٓ�	:|:��W��(�y������V.�7h9cQ����W��S���^l{�v��=�G�����4!fڽ��M>/�O�H���S�#dA/
r���`��p;�Ȏ����R�pvf[�����|�N=L��4��+<� O���1��ݭ��Hj� �S$?��18�������Ami��;�_G �;!��Q�-�Ӥa���3�����ݞ�M?r�-$�S��k;_����Z�}���/�(�S�5�'h�z��C>��XAr�L[�}���6;
�5����B���Z��G ,$��l��W�f��ɥ ^��8<�B�H�}Xw���W�Q���=�f%���|�%���Z�Ru��N�r��e��r�8��f��cTj�	�n��pDDM��T���!�_�_�3�a��`.6��Q�;�N|K���E�ݻ��R���z����ͫ��7����%;7��Hٟ+ɻOw(����T��zԖ�}\<�l3�X1����`�z����β*�y	|�̎����`�������E��,{�ַ�9����	��_���A���G�#<����Ui��nS���:(q�o-�|��gP�g
�/����������oj�cF���{J0.]�����xʐ)�Q�9�A+g�n�ke��3O�]��[�xĽ�Nk�C���G��0�%���>�H��bn!���X��T�C��=�?E_s��,R(��B$|�b��%�B���!��G��3V ��|�ט~��˕\p��j~�=a��Xp����Ѱʊ�,�)�7��"f:�9Z3���Ԣ�PSh�XP+C��p4�j���Q�LU�s'�-Oc���$�{��U���-��t�pEЊ���!W[2"oϡ��H	�PL5.��c�JC���"�{q4�,�{�w�	�p���hZp�	��6-E��?�zr��y5Sbz5k�YmU�:�����~�h0h������%�����މ΃���T�~����2j��Y��ü�V��u��P�M����!/K�UA5;��[x�<�v�C��7��ӆ����U�Ě��9�����-{���ܲ���Y��t70X����GA��;�ݡ�hk�	�؇N+�u_:�q�(�je7 I��ǫ.���H�
���ԗ��3��<�ru�O��ݦ���񒼒�7��0.����f%U+�Y�
V��y�[�-$3OqЀ���(��5O�XU*�~���&�v��~����a\1��+�Ğ�$BTC���u_rM(X�N6����=�9>e)��+����TKܠ�g!���'ɧA8O�6+^�U8O/!�"z&��f�4u��u<Ң�ӥ�G�N> ���.i�&����,��%�-'��u.�0��G
����c��5)���*�}���Ev&9{�p|��%�S��)<�L�ѝνՓa�Y�
��1�W��i��<+�?:=����du3GhI½�n�T�퉣�s.8�WB�h���0���nT����AI�$hTC1�5v�vnrR�/�|�iK���U��\ƒ�}�k6�9Jݧ���i7Nr\� ș	9r4*sB��$w�<�A-����(*PNQ'�v�~P�A�Y�{�l�Kv`ך8wY����|;6/``8a��zG���!���)w2����������:�CFX����{� ��ǟr%"o������і���a��j�������A���}�H��9�Z��t���X���`O�(Or�a-��?�
4�(�'È��'���#E5��Y��Q7P3]� ��� ��R+�Td�l���&���d#i�%���+I��U����(|7�������B����Y�Da�G�� ]�U�� r�Gw�K�X�1��0Du��u����R.������㸖�~L�C�*28GD>��۶��&�4��m՝���+�[�c��/T��<Wˑ*�p�=�4��3=���
�V�?��^ɘ�]'S�t�����[Z¢dI�� 1C��ob�G(�Zݳ��8��6�B-_ykl��C,�6�c%"�&�4:��J-Zg\Sʔ���Q�<��Fc������&��nA�趆[��WZg��� ��n�G�1�K��{΁��:=��]���Y!+�x�Ts�Z^_��!l|8���G	o>��G�Ȑx�?�����w.�YęH�Ϣ��}�\��S0R���t�����¸��J�N�_܃�F�"#V��zDX��~x��f��ҬK"r�[xM:X�U�9ub���Kw����v���VC/���Z#�W�uO����e����fT/��<�^Ţ�5�oi�����X`���Āb���/~`���=7fηI�r�1<I�Tԗw�h�j��q�Q�dXaxfJ�DF��e�2��5]��}V����8jNXak�֫�Q�(�˪��Z;��Z�2��E���0f��c�^�p�}����������2Dqt]
j�mԌ�
d����Ф�Q�7�!$��,u����5�3L����V� ?g��/�A~�F]�]쀌����-�����Ͼ5~؈C��|�����=���u���`J�ME����%�k^˸�:e���4 �K4/�)&B�aw����'��]��ʧ�,�E&���!������O���b/�'�_à�r�IY����lо4B���U�Ȥ#��m��x��d���K#�)�k;���T]�/�U
�~�]�t�s{7I��t��b�?�ړ�n.@�R8�jn�3®|+��y��:��#�]<�˫�)*�l/�u�>,Ƿ�t��=l}��� �!Ws�T��%pS�?��m��qE95�x�#��j���C��@b" Hp����^λ��u�?/��Qe�� ��?�®������8��K�9�P��8C+�g�6<�dӌ\1s辷�=�����vW�!,�u�l�p0.J���7�~�3�jc~ph=b�ԉ��K���Kۑ�4�e�ku��M��K�M0��<L�Z�kC#5ϱ���v����U�A|;�d�T򫰦�TBQ��͡&�qpCɣv�$�me��$�l�6U�F�Z��p��g�	���k�A/#�D�d�Z����/��`c�AQv
0��<�F.2�w�Lg�LAx�l��H�*�Uo*fqɀ��Nm`#��g7w,����E_ �0*��J0�|���\��d��$�sA�Rܠ��x���خ�����V8q��ڳ��Bz^���W�S!��䍖
����Ì��{�oPv5$�0i���ú���&���:��ب�]/!v�}$�}�?)���ډ���y�1��mv�%m�L��IF�k��L�Ts1�+n⠅�x�1�	����[ �����ś6&ԋA�����K:n��۶шGL��_�A�8�;X_���D������s��]!��oz�1��^qK�҂Áb���
71�n�I
�3֜E��t���*�jꅏ
;�֕nQ�@�w�@�<��	a�EԝW�NM��^��2l\��n�.����
K�\�@;�Q*���~Tse��xA�
�^"��I<�q㉩�����l[�А� 0ԟÏ�Y%��*%��N���_&�t�a��J�X1���rJ� W% zݸ[dЭ���n1��g��h,���p[���_�9��,ۚC̦� JKĜ����
�KR��_ ��`_ū��X�N.��%ɽnAӋ�P�ڶ0��:ꖣ�=�$f,q�0Vv��Eܞ�-��]�TZqG��|�֧�� "�O��A��J��g5��1+#��|�	=s�<��jC.���@�_���*�?z�\�
❂��F
�n\��� �PU��<�;���c{��7:U��Ћ��{�B	���]�]�ѯD�0��$�ԄR���	����V!�������>2ڤ��{�������������fr�L�:��F��qg���7Cƒ�N)3�*��X	\Y[s7����wJB���:�Q�~��ب�㠂�!>����������%c��~�4��6c�-����>٣�0
�9b�Ɲ�H"����s!�<��\?�f)�OeR��	�L����.5�����6H��YԞ���<�2W�fS��KN+�-8���[�Y��������g�$�.\Qs7g}/����&h�t��~S���Ϋ�N��b@�w_�DDS�4=��";��Tg���џ	R�FH86Bw�ӭ3�>�8�q��R)5�-]�#�1p�G��=�?j0���<���5ꝥGuW�{�@�7B�T�D��2�(y|%%)��}�]I���ɲ�a�h���Ð�*��Hc����g���������k�8�}��!�z���М�H��ŵ� 
7LAu�V�])K�8S�w�Wg�w^y�lƆ翪������*5'7�q��V�����e��Oz"��m͎þ- �(eX:MP.��� �ӧ�J������%�Պt��T�R�jz!ZPkSN�Ά��,\1� ���qwÇvG#��8��.��SJ�l*�&��$o�V&O�u�Z� �n\�cl�N�=<�4��;r��b>T�~e�&]
b�����3�&���д	��.�$�o3+1��ylX=ȭmÀ�����J47�	���n[3w�<." ��ɭ�Gx��q�׌�3���IS�����ĤW�K���4����U�^1뚡j�(ɭ(§�al��a�NKk�<אUź/����� BUM�P�Mᚼ���$\A�rU���q�[r0�y��_�ν/�/r]����O��j�F�zK���3�����.	v�}+w������x������ը��YgP��_]u�����>����4�i2�v����߫��1�ސ�)�[�ݔ�Y&�v����,��IK /�"��ys��.|������ٸ��3�X��io~�V6�%�ΐ����Q�=���#�C��j�x]�#d�1 �������V�A�a��)ȼ���pm�,Jm�>�����*�����<yH�-MWs��v�����KF���>���٭��5�&�┇a����&��$�qe(�����J,�0�zWf b�����u����漆$����P8mf�GK���`<�J�CO�1]k�Ӗ���j(�ϛZt)_���(avݓɾ�K�=g�Ey�)���U�s�3
^5�Q�0P��>wOC�(��#%8\���N�s�t*{��wz�������Ӎ�Ń���РnRqR�������Q'�����2lǈ�����{~S�Y���_�%{��;�ث>哯��r���I%h��<	X�)u	���*h(���&}�u�g~�M5�:��u&�ۉ�
u��8��b�����
�����M��nW4��9���,�h|�������\�?=
Z!��_�`oB�� �����",|O`z�XO����R��QA`4��YC̽Z�5�yð�Wt��H��/A�0^��������4g
�9�1'��rtF����cvpa� ���5WQ�ZK���k��Fc�n(u�U	%E{���#��{��e�W����"p2.��A^�s���al�-��	��P��8L���7��d�SKiL�����!�$Qර�A�=�Md����XE��g��װ�	g�DrY�C��_�ۿ��+D/�BZ�N�T}70�(e���G����x���˛	�.�P���*��4[����d%E`�+�M3��w�������V�!1��UhpHGM�kƭ�Lߞ4�r�&�������GpTuy������f3�/Ք��7����)i��¿��?�y�	��kya�U�H�1.��[��3���t�4��R=�����C�oQ�o,hO	':)���d������_T��lo�-�f��L+��,?�	@�T�K�Y�*pV'���TN���_K\�!m�v�8�zӊ"e��b�:�����)�Ej�׿���9m�&��a��*���%��]����53�&�
�hԤ
�� �ʔ���YC��K&��Aw�w� �9+�θ>\
 �V������o ���zMo4لȐ,��z��UWF\�Z�_^Լ��R/��װ�V�o	�J2�t�/~�Ų���p�`	�n���V��V��Z/'�^�[Ff�{`�eC���F��N���/L��v�%�k4ξ�ܽ�I�W`g[x/�if�C�Q)g7~�{�ep����o|���L��E��֭>��,٠��k6aݡA�4p��lx]�!,|ҭ#�����!�Y���؇as��)�������Un��kЮ�lC��S�m��
!WB����)��@m������9�қ.��_�g�9B�/�")hZ�n�2LgE�X�Q�Z��¹��>��<���O��n�I����~��;y�e}���:�� �)�+^��KaN�p� ��1�Hg�� ���(́<aE؋���!n���k
ܪ�1
@x撚N$;�1���^.F9 ��2�B���o7�����9s�?�%�I��<�����Y
l�H$��svhFy���E�TZ	���rv��5vTӆ�4D�K�m�.���;BY*6���Q!�0/Q#�j'����C�֮֘CV8{EB~ٜ�<�R�ss�Tk#S����b���񎯰���� x1�6��O�]!�.�ĵr��V���~. �E������)���'`�ӧ��F8�µ���Y~T��אE�D�g,��a%�\9���_�~�|��'*!W����al�e� ��d��@h�T �T2�%��!j���l��E�G}{����o+O����Aj�$}���/�D���P!|m�������D�-M?8=��`�E(�]C[(��:�>�AY�w��!>�y����'1u�=?�ӃB/=$��5��i(l{E>�Aജ�E$o���Fy�sp:#I����9�,=�⅂��D\1�7��~\�q�A��E8����!EG���4�yt[F�|sR��fSwh��Tf�Q~�& ��>��vjT��gZ�!"f�����1��V�Q�R�k�3�҆��}#�4�˴q���_���O;�"r�\�X{��2v��Yc�2A���^�k���|�I�hU��-��/�&�ό�Bt�j�B���֫�1���.�,��O0��E�I�G�����"7F�4H��zS��T8�\���,hZ'��Z`H{h%9���<���v0�	-�y�[#��0O�'�� �+i�SEs��6�F@ǰ��	(��B5eƝm誺.�g��e��6w�c^Ĕ�$�
��&79	N�x$ 5P�+9؂I���a����@{Y�&Iݯ���~�����օ��YX;O��?=�e������ 譵�����ҭy:$&�)���z9�-�c�;��q[����FN�	Mqf(@�I�
����\m�.��'QI?���{d����ol'�cH�B��Q^Q��<�;��JD?�m#�	�>-F%VjHr��*4�/U���d�Z0�l(aj. ��K��
�~߄��^�G!�9 ���(�<�1 �%����uJ�|`�Zd�9�Q]5l���)�-l�M]�S:u<q���:к1]#�*;���1㒡����^��x�x��6<�pȘO���Z�:^T��7_`�Wi[G��:]x���~Ɵ=��t��cP{Ɏ�?�#(�YdM��r�,���8,�^x��$p�
/��͡�\�:���n�|���c
�b�V<Ɔ<&CY��ۇ���:y��CQ�W�7^@'�,w�MJu1�Y�eA�5�lb�RY=,%"d2L��0�=��A��+�j��10��El	�D�?�R���܀x��3V'�qH�!n�&6�[.nQɓB�c�ƚ��!4q]X4S~o���@భ���x�M���^G^cI�N�W`��
	9�y���;闣{�o3z4�kj))��T�Tvf�n���w�>>�%�F6�Z)t&(��c�r�Z�8;����Ghm�s-��<u�{$H`R��_H[{[�y�N����~w�y�H��RZ2|o��En�u@�Z���P(�N�-��^�8��7�׻�2�����ު�z�dTf�wR�xb�y	c���� �z=2��ī�t�a�5=����m�M�_V�:�x/�z7Þ�����,�^GR��N۱��s�	f_h��P��Q'7�)�~�vq�0 �HzmN��w�@�3@hƪB%!�a�.�2k���(r���K��(#��Ǔ/:������W�XM����x�W�D�p�F_w���2�&�,�������iy_����z�%-�2I�{7�����>܆*x��x��� &GZ�Y�V�Ԯb����]>�x���&�$���}-��l��M��?�u�����e� =	�j�c�}_vG�|�=�@�A�IEp0�a9w�Ok�L� #�a��Zݡ�4�*!n����d�|�6�6j������=���4�:�*ɟg�*�5TLP���p�����a���о� ��y>�M"f�:�6�V��)���C��J�,�x<��)��Q�_�����y� x�ws傏)���c��B��;���>gf�n �w�8^E�&2x��uE&e�dAx>�TX%dM��Y��4�M ��5 >��e��u��=1&1�[�'��Fk�	�`�#3wvӀo=�:��&�c�[f�A�����yA*���b�������"D��b]Tn3�0���A�����6r���i��]�+��vN�6&�O\�Eܚ��3w��9�|4��P��Ĳ�j��EU$AH�X���6P��w�8�q�_. ���p
��I��go˳^!��7Z�ͭyd�TS��gJ<3�_�F�f۲l	E͐��a���:,5%�;Eč�������KEJw�َL��jI¼)�wY���x w�dj���e��-O�\W=��C�����ICڅ*	E��Cl�eh����B��ݽ}�.X�d���� m|�X�w�l���A6nKx�)�i���i :��pj/��״Fj AI�ﴯZ��D5B����A�L��r�7���w �I�C��\ID]W!���@f��.��vd�H�q_�m_���I��Au���jv_�T���P��� t�2��8�<Zz��h�׮����+7�in� 6����� x+o���|}E�Z��쵻���|}l�n���8�ɮ=W����W"�: ����?��¤JAJe����C����~{�G�y�����~�G}�&+U�k�i�wr�kn�P��˾'g����Ff!~�s�=_O������1.�8�ǃܥ��;O�G��^Aw��v��E9���;�1�Z�`���9W@���׮���k�uI�>s\C��<k��L a6
�ϋ����:����'-�|[|u�P����s#�:nw��H��fSW(������T#��%f]a�w�D�&ţ���i��꺍�����ҹ�/��6��V,AL�����np�����w�Q>���3J�� ���2�dwIH�s���H`PQ��~�[��8N�dX��k�e%F�ʤI 4�B�UR����2�K���5�W5��隈^�@F����`p/E�\���x��Z,�����@�㋌N�&1^O6�j�Y��R\[��"���
I�D�]x���?����� 6 �Z��!�tIs�>��̳��?)�VaI~���*��QK�k���' �^xt}&<�6qX�P�	��u/��xஔ�"��*ļ8�QD�̑�S�#��=�ODA�����j�\=�4l7���Xk����'Pi��`�"��r���m9Br��W�AsT�hH�$�v�`���~	���W�x��B����oޣ�dH�k f�����7����xaS4�tb������a8���k��
)��,�@�v"�n�gj���r���U}�x�~r���N��'hMH��s�H��:�š7� �#��J���S2�{'Q���=���0���s+H�吃��O� 뺐�c�rt%(	6ћ~�jR�c�#0�� �Ř����~c�7=D2�zʧQn�}�5jIm!l,!�����Yyq�y�&�_���l��҂�2N�z���0�&��5)��M-iU1�ʅ�s���&1�����@]{vN���`�}�� )G��.3tk�7��]1v�����'ĸ$27�Ԛ�o���RQ�(<�\9�u��ƳN���⁀z�v�c�#u�m�'�G'�8m�Hة_oG��%��K���Ү���`���Z�.Ч�ro��CKt�tYìȖ�8��I54�<H�Z
zYȭ�3� t��WqN��CլE�_���|�&o}夨
��r�����-��P�D�,Y�S���7���6s>��x筭(f��k��1:�O����-�P�!g,���>q�eZ��� �9g�	�Fb�6??qiXZ�3�/`$��ՙ����n�~݅�RF���p�z;0ߋ��}���=sz�l���.p{:��f�،�->��T>|��ղ�*Q���p+�8v
��8�`6�!וAY������v�I�j\�=~�γ����+����*�Vc�7ķ��Ӈܫ�Պ��Uh�ٟ(����T&l;�ZK/�2����O~�%Z
����C ��C`���s�6��B5tX�y�E����y���4_rK)g�r�)�s�X>p�k"g�JljY�Db ���Z���������[h.���V��Y�'P��&6�~�,��^�ɵu;?�=�BaT��hp�<w��^K��h���WX~	��̌�vK�A�t+�bُͭ��D㗓��ړ�ٛ{uh���#��0M�����S������P	�HMA��f��a5����{="OC�l����q��X��؅X?�a���=1`�ݢ\�F��d9���q�Q�1	�#hy��LP?7`ꝣ�Xn��"�ϴ卽?��K;��F,
�G]��k�Ez�?8T++�^iP&u����Z�)�$�����P��s�!0&�7R8�"���uvnC���>�a�Q�g\�h�p|��&v��E�;�����G^���4z���b���칎��`KA�嫘g�J�r���i���`	�3�����������i���V�'U�v[$3�&�ي� 	R�6V������Ҽ�Ң�*��Z���2f�d��������iYI�L���6ǘ� ��p��}P�@��.���g�u�9���4�}K�V��>�EX�7�Zb��3tJP��?�K���Fc3�jd|7�r�O>��W�VG�:�Q�Di3#�Ѐ��0t�]�q��w�I�6ig�X�uyܙ�|G���D�s��G�����ȃ��^e\�����hɄc�4~)��f��La *uzr^�ML�����ʰ}C��Է���:�;ȶFB���c�� =u;k�x��<g3����~�F�Ow,ɣyG0Z�FsY� �K1�~�/�x��������o�H�mL�sp�� �e���g��M�c�Kg��ßl��Vw5~��Zp�v�O����l�`�xK����e�ik�������oie����-�D���\.c�%:h�k	�W���:<����E��ҳ��Dѭ�7�4
F����1_�di:�.ƥVm9bV=0Dq3]��F�����T�,� X<}�`�Ny�;�u�����z�d�� �5���K)����.���Aeh�m��ÄQ��F�MHz�l�0���`P$�2DH-V`��|s�8ގ��m�I��嶨�cOB�e����mK�<q枊��2�ޥ&��J�-O]�:>�����463��d2���T��T5�~؂����/j<b�l;�,�����)ֲx���W�����5��)��������%�a�ªC�x���p�_Dn�)�8�gx���K'��(^���o��YZ�ȗI�n%�E��S���0K��Y#]b"n�G�YMz�T��W�3�8ׂm���q�b� ���-����R�7�W��fr��Q��mK��rd}:;�B�e{|\�5|�j�1ȑ�B��<��iZ�dt��-�9Ͽ���𹙚��7�Z\��p���{��5�24��� c�Ce��V�q�Y}�8�t�:��݋��}��S'��Q�k��^��8l�N�ay B�4�щ�0\]��?��d�L�w�˾p{��:�D_��|Ѕ�8����D;�5������!���i�#�WPU#!?7���L7A��<ƴ�G,
�4�r�aɢr��S��<��cH�M8�8k��^Jj;���-z�	���4����>�o������zK0<_,vK�9�_xF�x"�808�5�辇DR���N�~�N��|���$w�Y�R���va\؏�w��YN4�/^���<,���t��l^�!3U���iY���5u�	�*�ߤ�����"��|w3�n+�6Q]*��9t��2۝^�re�����.����dp�v�ˢb�O OW	�-���;�@WTz� �*��C6���֖�Ywk�N�1,�k?Wd���8�]m���4�v�d�R����}�db��E,Tmn]��ÉYQ �l�?O5%V�E����.���NJ]�����wE% 6)D�{�e�̟ϟW�TeN�	BO�@�g�Rq���G����a�����*���ؖ9/��Z�.���O]
!�w�W/=�	)��o'�u.gh��ah��fߟ{y�L<�R�� �#��_����T8�j�RW���df�T�n}��	9>�����ف���s�
 z�F��/69��ZC�i>��Qt{�
��`t,�x9b�-D#���*��㛪�`���0�ϱ�� �x�uB��<��w Zm��HuXqo�g�`���,;�P[&��������%��3j#B��	��f�&��kC�`�7":�-��һ@�ny���.U�p#�b{Oy��2S�|���Ry�7�2�ݟ�f�G�l����3��O�qCP�p%��%��Ⱥ�ӏ����o�.���7�xT'2|��?a�z�7u��a�/�#��6��y�[�{)����3־R�5�%�Cr�4)�SK{�����W�����A�͐`-����t���0B�~e�1u��-��s��OP���N�t����^o�]��5&����;}C�5��DKc�;�F��mQ�C���fӧX�S*g��7	�*�I�Z�=F!G@���I*��q�R�e�����������(�V��	03t�?B���[J@ߘ�?%�U��I>/2A yzr�U/���4�.�|,��c�f�09�)�2�p�ˈ��!�|� ڜ��N��΂���բ�[���ME;wP��p�'ڋ�ey<ٰ���ıDu��s�[��%��hc�N�����ƕ>��d���������3J������U�F��~�]c��^Us�/rh�&�R�X�&O� s)��J�=VS��#���QW3L<�ǩN��eB&':�1?����������;�)��o�BΓ�Qz?K�o��Xn�<������|m!��y,RO��ij͍����y�ܙ!�Hd<6t�J�#��ا"��"C�L�](Ge����¤?�w�W�!����f���kq7M'�NEHf������!4���)�2���N�m�>v��eA�� ��Ì�:��g�7ݘ�)�o�Fi�qt�V�iF/��=yv㕗�U�݈
o��c~��jb��u�Kd���u��C����Gi2��D��}HE"�t �� :	�d8\��mH#�W����{�P�9b�~��� �9�3A탠�!���x��1e��u��\���;},Ed��il}�S��¥Q�q���қ��7,����w�ʰrz�9E--~|<f�D�!MI#�m�2}��{7Iek�����'�W���x��a�@P ��Y`IƠ�Uئ�cr�h�(y�1d؎��=6�G�'?X��>���e�1�x���؉���p�]�|�.ԏ�L����,��}�3�m�),�ֲ�!��aROH���P�8��gGV�7R�@�B]	�O{:1���9Ǚ=k�C#K������AO��DN6d����[����?*&qL�P~��JM��25�}_�����ғ�$b��3��Q��YNn�C����fk�7ҹ�M���
|��H���)�4��as
uZ�gC��"mm����#��x�����SI��{�\'c�nue��;w	Q���n�k��%s��ӮQm��{��L��۱�����9�R�
7K(�V�����i���,�|�V��mnG!^<��p��\>)���a��@��9J�t�t+)�/�Z8<������t���/�EM���jEsԼoS��;^���`���'8�G���1IY���*�V���v�ޫ,���i^�ځWj9�'Tɧ���� X��\��S>���.Z��:�Y���K�	K�s���֢�R��2b+RE���*q��kU�{�ތM���(A|F�-�&an���.ϓd���
������Q�-%�r~�/MT�}ͧ8����+� #�P��
���q��<2Tq���O#&c�	���c�c�%\q0� �x�I��ĻA��/�R�]�f�����Gf�Y���,!3���DWm�O�C�r��DL�%����0�,l�C�,C�4Bj�CwAٗ|[A0Y�B��^�`3�31t�܀�`	�h�u X�2vo��v_�),���zv���*TT�М¿۲.�̥�j��̱�r�D%G�G��Y�B�s3I�0~�G%�	A�m(�N5[W'�]Oo�Z�C$8W�O�[��Cؗ2��/LRZ��)������uzZ69-y�2��
�Q�P��g�D]��D����y��R����9m,_N(����Y�z	���f[k���)�]���wx-l�&u����+[�H8$�&~c���0�F���#[<�-](Qw9��A��.��EӃ�]�1�����l�@­� +{�Z*�W��*Q{h��'�(�]�:�K�ڠf��;]�,�n���l~�jO�w$�t���f�q��٢?�	36��J���iͭ>"z}jE�-z$��T�B��a�>��G��BP�t�۠2�8+�����!��Ň�������!� f�2����w"����$,A9��ׁ���ˡ�p�F�E�ގ���ܲK������%�^�����o�F�L��@V� � P�x ��'�M4��mrN��c"�nՄFne����p1�A`�c~k�cu@�s��\Ś��!�֎n3oR�^�4������}S�=��|v^K#)��=��~o��XȪIK6L�'�[�>)�%*�s#�g�� ����)�7�/�
�xB�=�G�+����@�ћ�}9�Q�>��ǚj�|+s}�h{�+ �|��/���O����7d�@�ײ(^q�Օ���̇�=�A��&�K�vR�)�SLS���q����_����3���VC����K2�D7����~����ֽ�d`�#�|��0�a ��X<׌���6ʼ��ɗ�U�S�&�gb����C^����8@�&�����P���R\�T�qd�q;�* ���5�>�����y�y'i��#��ܶk�z�|��L��b#9��V�_�����=2]��>S�/d�Mz��L�����!gBI4��{[���,���4|�W0�7�`��hG��(���f�7�ͬ3��c\.`�L3X��Gئ?f�����Q��\��d�a�$��H��!1V�k�P>�1�5̶��8Q��(J����"5��'O�]ee��]bߌ�"Ȥ(3_��I�U�洺���h_�;m@_=�눻��Y⇥�p���fm+-"w����ib�g�O4:��4��s���%��6�v���7J9g�H��+�s��E��gq{�M��~����D8���3����n�V���-Ǽ��#|����U���tPٵڪB�]�a$�6,,%��z��Tե������ላ
R��8͖�2�O��D�x�PH�s�W�#7��� ��8B�*�##�9/$�͝��}.An��f�;=����hX��o){aE�lU
E	j����j�E��ћ�Tu�V�3p/��r[p )�
?�f�hR�Yޒs����){ֵ�
��A���_7rB�uF9��%ͮ��|t�pm$��3rMS�\�_BW{�$��)+Y�."'�:5ͨ|mC<|LB�WN����w;�W���Ő=��e.��?A�c�>b+����~�d�Ͷ�f��/_����՟!�E'�����'ҽ90�1��gD�V�G?4C���c`�q���W�;���z�#OA����c�k���˿l41Oy�D���Klc=��CN@�ʪK(H�شؾ�M���@v����[��c�h,>~�+��5`�΀YV������NPt�g!��$����{#��b-?؊����f[�g�F��@�� �ȃ�9hAc�-Iγo��M�ٗ�"C���ڥF�SL���  �#�1猰|4a̤ZУ\Z�%6�Ja'�rֶ-��.�w:������݃���v��plfB��^����&\Nց�jt}�iӄ >J���i9��I�}u�,@@8� �457�gs�uG��ᆭ�W'p
�4� RW��^��=�G7�WB�]�4�(�6�޼>�S��1rF&o�'�u�
ܿ��-�t�x����Z�o�-T�if��M:�ĩK��C��"*��B��`�{6;s��T4�sv��d��-�`�kxn�������!)Yx?b��@D��]ߏS���������̬	���o.��]
�<Q40l�յ�O�+yi����n"C��i��_���mfXZ�E�4�4��Z;�&
� Q���&^�����v��#��F��ş������|9�ls͆I��d5��=<��u�����!K���뙽�O�+�ɛ|8����z�.��ZN��)�G�W?!h��ﺦ���-pIc����՗�6�c�͐�t������p���_hM�@�@�P,�Q�*�դ>8�$_�J��SIf|��^զoansx�6Pf�v�g�l�Z��d��_��շ��8�u���fQg���vQ�^�2�Ui�\�=A-�K�O���Y�R��o��J^6.�ˏ��9���G��S"�/蝕+vײ��2
sah��Ea�����^� �ő��2������8�����s ��E�j���<IPP�D��)�hl��Ц�t�S�-c��5�}%���_%��=)V�it�È�*�ٰ�S���ǰ�vvp �Y|��c���!9'h��Q�i�P
^�X�S��-VL� �L�}��;3	��LO�s�B���=`��h1Q���u�X?2���[e@�m��$��墿c5�`|� �k�P	��<��1>�<3����O�Ky��3/�?X�?�V��!� 5�9��F@sti������V����i��]��hb��մ�<4���Z<Q?)C:r��댜�0��-j���Jjr�4Cs���۱��j\գ��}C��lS�	a��Q� ���Lb�-�Z��:�<s?�1"ΠmL���vc��0��&8K%@VX�X������2�ɩ�a��}�Oʑ���@mv����-IڕO��������r�dhE�}�N6�1@��~��� ��+��V	u�"i�N5h�@�d�����Z��zX��6���oo��SӇ�aLM��P���Ԡ�	��7	�_��Gw��+&ۣ�BϼJ����L`j�iU��9;$vdF�
��?�-1�3F��[9�ϙ4�fĈY��I���)o;�$1U�h�:��%yi��x��FE�Q&'Q+D��z�C���,�\�Z�]���}��*�^�3�ޑr�c��^	 )n��\@�K��=���&O��qe��x�+˥f�f�J㺩�s_z�q��K�{X���d��� �~'&x��.ViG�g��\%�=˅>W;փW���w	�n�@�+�8`L)E�[�c���;�}�ml6�9��7�ɠU���`OG���F��v����+��N���z)��\���*ȋ���ť�j�C�����k�.	�Qg.ϔ|Bʬ'.�;��޴_��O6����jHح�љ��蹞V<��$���3,e��D%7�G�(�BHK5.V��:?l�q������b�Cx��M'���9����~h4#TЦ�X�R�1bb��ȂeC���^I��
޸e>��}'�5�C�Na(�P���zl	$oM~����Ş��Zm��g}J0�@�e��D�ً<�����_I$��ƛ����pZ�O1 ��K�2?�MZ�;�oJRA���Q�����g�Y�,3lm�{�',B1��"nԲ����aLDfz��V�`��T���x�[x�9_��V�s��_�˃wԎ�����rAU�/FT���lB[���h�A�j��2R�Vd�dÄ#�Q*<���`�x040�|L���|_���Dmɖ���A�W�a��@d��� �A��h�d&#b�!�볦�8��ا�m�R�4-����p8��?�?�j=�F,4xVA�`��xC;�a�����$��> 7v�����n�Mk31a��lF���LNoR�YLl�Q���}�&�zxhF������w���b��Ur�?�Ԑ� [�Id\��0���C� ���#����n
��n�HG�n$�9��iI�,���dn�a'��(�uP�,�{(_�7c&���R�Gm�[�_�3�q
��+2?[��?�W_b��N[M�bu�V�ڒz�S�9�9��M�%x�5�܁�C%a��s��f
?7�j��Q�B&���e;�ɷ�H����7���+�i2�}���3�.L�f�H���_֨�������Wb�P�� �އ�V<�@�����&�^�%���w�U�3�h��k������Cc.j�na6�����Zb3��>K�d���w[^�[.��tVa�竉?�R�ߖ�u�+E
�a���d�<���|��?�^���@�ef�,��ֱ��h��ՐÛ�{��U*p+�B�T���(�g�dV� ��4]��0��r֟�:s˷JÇ\A�J�����+}�,�@y�[�e+���tqMݧ�2�Yp�*�^D��0�5�}�O�?5h�24Dx$K����"��l�G�D�����uʎ����B�@1�	��V�qX4d3�t��>A6��������o��3���a��/�0��uw۬/2�٬(|�-/9&�tks��N���(�5T���*ўDm[���H��8�g��P��.l"�k�}��	ZP����a�e�+@e�n�ޗʂr��(�x<����;���kY���.�����V`>zŁة�R��.mk;-2�N\�~�u6��+=��LK���l��g%+��E\�i)+0 ���$8Bn͘�'πyμ���WC���eY��^����~��+YYaw͠��i��������i2�����dl�z"/Ys��*te�A�Z�ݻ�������Gь
��D(��0�OAc�!U*�m���f��s�O���(_��k��g�#�����>�4�M�_y��0 Z�[!�H�K�W��:2�"{�t�N����I�'��\���&`��&z=A�p!�
,��{+�ȓ��>�|�r�~z̬*��ݸ˴O͈���]`�,[�>��P�~p#�)�ca;A⫇a 5�?��[��� �b{5{�Vb�l�R��٣�Ųj��~]0�� s5|�#��+W�*D� ��L$T�]ɮOY�cR��Usʒ�F�~^��ђ(�}Ppf0�w��w}������z6$�z|�e�{�=�{Ŀ�6)��"�� ���o�]Yc�|J ꎉ���l�`�!QB���&��ϟ7{������������R�<LHG�/�:��+gt�D	��@,ϴ4	1o�#��:> �D�q�E����&� �j�˄�qc�B��,���I7�?(tؒ�Ӯ�#.33���P=�B >�)Ĵ�H�}���v[�q�����]�{""3_-I�#(e&O�q�f��-����5חdi~���M4�`!�����BM���M5������!�m�e���+Y���a]Eoy 4;�nO4��Gi͒�kb� ���J0�El�N�1�;Cτ7, ��:��(\�{Qmz_q>?��|�ՃL���)C�p�,7�
R�o~Nt��ª������)EN}�gxu�Yr+ � ��
�S���}u��E�$�i��[�|�uW���q�9T)L� 347Hb�� 0�yZ�*���AO���F�
-�UW����<]������5^�G�\����Ɍ�ǀl�xeqJ�ef)Ѵ�P�W �X�F�َ��G�Ҳ߀^�=�T���L�Y����~Yh�u�W�����+��$)kT�<oK���_����OY�t��_[v�1��\{�v�i�����0���K�39��ʻt��G� ����׆HP�i����g���K<K�qGV�Zm+��VQ�WU����4�Ϩ��CW������F���T�"�2�Z�l���#�ڄ��F���QE�:�na�'�����%Iwׂ�����av."���Kz\�ŏ[���3j���f����a�����5�ό\�"�U�Ï�����g(�Ea���$���!0�T��YL�)qU�\GD΁�뤘��4u�@�"�:9�N��0��Ou����t��s�o0��Htw�����	u��b۰���?�j]�zA|?�>l��D���"Ũ'4�3����آ�]4��Q�����1��V0˖_6�p�i���� �v��&X9�f.Z΄��p�y<IZ%�l'L+^��L�P؝
ε�b��s �Վԡ�zcu�<ZH�H��m��1��7��QRM�,�˱+J��qH-?5�V��J�3^t��bn��J!��,��W����F
�S���xL�,l�T��[$�^_,����e����.��8K���{��39���Mc��"~�}wx�V�ZÆ���x�~��KZz�e!Բ#�~��0ň��cN��SܲGJz�R�d�,D��]��4�ƫ����&$e�E��đH��� ���!,��J�\��3ᐞA�ēl_]�W���
t*��SFXdg1�����Ns��L����;k�_�׼����� 7�sJST.� �rT�'^�@*�I�(n�=-�]K���N�H&&!;� 7b�J�|�r��4�+\���n�q%�K;�(1���o �;�z*����|�s�F�{�\��Ē��ؖ%�~���+^�� �kY�ײ&t��Ϥ���L�� �Kz�O�������\o{��
�E�b�牖�h6�ڶ/!�#�R��~P紏dIr_�ؐ-f�&{ۖ%3���yt���,l�d�5�v^��"�)�5]�
�r���>��;rY��*���#%�E��lψ��?����W!3H�d2��{�
����R�s����Y�?u˟Hn�f��q�@� "���R�[k�ӭ�r;�6@Wz(ۡE�#b��]`��~�M)������Z�}P��E�|H:�T1���5a �͸�Ro\ˉ� r�3���m�`�U4��:۩���i���*|{�h����Ǵc��>�\���k�V��;��ō�o��E��m�q0��������j
7�|]��6N{F�ќV�h���s�⑏=�7V���%�L�r=~!�~�h�ĵ6�j���v���T�<:���0�QL�(3,��uݒ��()�A�A��D)��:�zo��>�f��!�nw�5 a�1���H�e� �h������d�2++|�J�UQ�9l[����׺,M�v� �0�gga����\~�b�ͥ��-�+���u/�Ņ==���s߶�g�@_��Vg(�~W���{J�3�����e&�Ё8-'T���PT;J4�aL�o��8vL��e4�x�{ԛ�J�%�xw�rH(���G�,��V5�ʩl�c*>��u1�� 3M��`m��mv��m�k�_�	X4��^��ɞO;l�\�Gf;�z#7Tp _1J���ևz>���۞΋��(�r*l'���2�xϋw��vZ�ۮ��Ԝ1.��$h��#�\��/0	E�E3���#����g�������J�K�H.ƅ���H���oy@��|�sb֢��ߎ�Y|����I�k�7Z_�p������\�&f��V��l��4��"��7v)H���ǫa�=i�vW��$�k\w	���U�K�� PU"�ڵ����j�����G�B!���ṪU���*�Tӯ�Xy��	U�� �����n4�	?-�Y%� X�W=�Z���^�rDp���%��?9b��Irq�qDF�)P�k��%aH�ִ��<�� %R�kᨄ�T�Bw�y��/p('��0����ɯ��7E��K�(�)ю먳����2��i�Ͱ�?����m����dO�|}^��IQ'��qs�a7��F�ɖ����K��|�_�X�����[�З����z��j�J��ii�*�@�R��`mM�σ���Q�97;�g��fH����ߚ�)��+��޸���j��W]@︲z���>��������&a5$Z $���+ˢQS���fGs���+㩓�x���@sᏆ(?�t㊪Em����P<��47Y���Ҡ�W�kէ�7����@�(v�G�O����bM�4�3ʆW�.�\�5��J}'%�@�2ôI��!B�bFк�Ggǧ>�P CY��S�j
թ���S��,��/�{��5��aX�H�<�|Q���d
��a3;τ}�A̼Z�^�B���4��.�/���$g��T(�$.�3�GI˽�cn`�#�L��]�̒Pu
|nd��̵/b�w�i�����L�_`������A���Ē�6�l$PH]Ć5aH3ybl���^�]%
HO�&��z�P��ѐ�xV�*����R	h�2�7�@k
�ѬTsL7g�*z�F/����k������h��pk�O��t��y�U�p�i��x���d��%�_%W6�{ �ą��'��������F���?���n��{K�xm�e��U*�1%K�����b)PH%��!2���������M�r���ˮ�����x��WeK∥*�q��8"��~����*v�P#���m�����
39��$��r���uR�me.B{��$�%འ����'�܍�&�$�~R� ��mM}
0	T=ɮ��W�h�mN��%��T��J$��m��R�@Q��v�� D�4�:��̇.ePjJ�,�I��㵬U�9"d�$:uk)x6[8�m�07U�C]tby��	@B_H��=�Ŧ��Z!��*,k�J����A�D{B]�=`�e��M�9[�i
��D1C�?��m��>jU*����%������1���v&�ђ䧹��hz�uD(���6"��/�K#n��o7����L
��g�jW\��{#��!�/o��.�?�!Q�c׶�j{&�̼Yx�ֻ7̪O�ɑq��p�Y�"M/���bul+K˫�+'P��2{Sh��V��TOzN�Y}�:�P}#Ԛ���ٽ7L���Pd��o�Y�;	[�N�{64<@�%2�bPQy��Fm��S��5n1=@W��v%ou������#�c��J�k���#��~<�̮J���1tu�j���H����(�-�bN�jH�)L%�ʸ�����B��'��E�d�U���H���~���nt��:9���G���n��cD�l%���x�-9`P�HX����/�3[���̠����!�6a���v�zs�y�P�6����J�"s7�~��	�=��qp%�*Q]�Z�wǼ���ӆ�	�/TG�H�Ì
)���#�ҠN�H�Mƍ["�b�qC*>���i�^:�����i�����ڢ�IAFV�oM�����Ń;D��!0;A�$ĠA��np�Y+�<'���g��WPSտ��yF�~�}������~��'��9X
��N�%� �!b����M�U��zޅ!�?q����������3�u���Ej?$9{eXB��J�m4��,�$���
�pdX���=��o
AFJ�����f���{�g�EZHt��avk��7E?�y��I����p�vQj��3Jٻl��Q���=4vT���e����뭉�������x;��6_�M��΍
w��$�@�I~M�|1W�A�,�g�˧PV|��ގ5�F6�s�A�:�B&`�9��U�AM��+=�l�gʅ�ףڷ�Q�5<�?-�WCF��P&�7gH?�ܔ�_d��q^$.8A�6�BjH��B��háS�>��
��.��UfȂ�
�{�
*Ћ�,~��;Ͽ�@��~;��ޥ+�$7����i���ժXK�6��گ������)���4�����yOy3��T��KQ���ڰ�n�i (��ٱ�$}4�j����ӌ�}�Q1�X	4tʳ�%�P�X�vZV�騍[n��q1M��������-�UV���m~k`���gyR3V�8�Wx%���?q��N�uS�b� ��Ļ�<ڒ7�ﺟ�,�Ȋp�� �ORT8��� �l�,�T�{�(m���W��́��S�軣1.�-��@��׬kd=�J����|�����7=��|�qi�([��j@_�[%L{���lJ��W�d��B�l	���'`=��:�2F�X*җ�]�*�P�S��t{�A�Ln�`W���1�U7�x�Ie儔���P��OQ�ks�*��Z/��6[h lHfhPi���ߡe27���*��s��*	��[@]������= �|$K�_�p�+���na|��ʻ���1�@�i�PA�x� ��[Br�oE,u�s��%i~�Y�k�%!".��W�S��詄-f�]��c�۞'a��KY�R��_�Z��~���"j����k�0��n�@=�Gkꇐ�)[�)��=��t�(���j
�&*#�r.��R�t���JW�e�5׮o��� n��ǁ�<�r͆�	�g$�c؉ K��+��O\���y���.�'�X����?)|Dޓ�S�+ �~�3yM���d�a������X��ڗ�"�KS��/��d\a�;����~�S0�'Yp9ET��'3	��A#� �>�an/��c�`hhl��sا��wM�ʑ�Ց�g)����Lms�x?	�<�"�qK��}�-�7P�/J=�@S+"9���d�a���FP��u
�y��
�E�V�/�<�EAA�J�,�ׁ��4����00Hk�K�Y$��m��Q�/��i�L�z}.D���EI�T�o�H.��_�ً�!α��l�=�(��|E~d>����,肌S0��a��o�G7��t��۠C�OGIfuo��||���s�PԳٱ�Ho���%�Eh/��/�2gy>/�ya���u4ٳ#�=mŧ|�<��a+7u�����m^�5C�V{;��֛f�z7�m�X�e�9�de�T+�V�+�?B�h�:�pM�QقMD����_��q�)=$+P�We8�#M}g$H�1��S����-�_y|�@����ܠe�T{q��˒�e�c�w�8>8�ɒR�.�S8l`_��EU���������p�I�bk�~I��Ry�28٪'�G�^�ED��j ���5��N�_5M���Xc ]��8s(�-.� 懙Pk�<,�,�J�P�V<��������⏜��Z?D["�Ɲb������8�Ŝ��� ���\H���J�{�hpL|]��,�m�*����&��]���t�Ŗ��c�R����S��P^<�������lc��8mK�с�G�%���F���$b·���tP��K�h�kӘ�ؐ�>��n�mϔUlw��^�v:I>�lޝ(��Й �nn�,�޴�_�����F����Ԧf	���z�Ԩ)�"�0��6��(-�`�?�(m�K��4�)P�u%���;[}�R���u���D�u�z�J�'}���W`�T�pL��Aфd���w�a������.��D9�%�������vz)�kh�>��@XSL��>��V��n��������������� �-�x��/���l�W��Ǒ�?�YC�<��b,��q�^�L���M䴄�/	���#&��U�`�����E�f����T�#�n�j�A�5��Z�Wu8���.�^��
u}�?���҃"��3�z� ���:,�/����ҫ��W��2��N]��8%T� ��e��ƾ7-�
Z��[*㉢3Y)3_x��4�:ce7�V�k�S�}i�ͥ��T-j/��S7w�gÍ5�mZ���}�`�=�ӹ�r+2�R��n��r�J��CQ��uo��k����T���c�45$pЕ��l�ߢ�2�%i�k����9���ұ�L�FƉ�P����
����Eh����]�a�~�ђ h�kz�ӥAS8?m�Au`~A٘����C;�M�_E�؋��N�!�~�?�N����9��r�����t��zn*��K��:Xn*l�I8��;���ഊvZy��8��A~�8��Ĉc��[�͕t	tm����~���: ����ȣ��g�xX���cT�����ОQ���h�;��i*g���2�F	$�n�c�hf�2�O���gx)��G��ӂ�T���=uC��/�7�R���g۠�e�G
�AP�[�>�{Ta�	J]O>�Rl2�a@�Ye��Y:E�`P���ޅǠ����1�5����Lӈ��bgU��'�H��7�x�j�A�i�v���ݖO�5��qs�HRƈK��es8p!�`����T�����!K���)��6�*(- ���8]��YϐsR�Oė�Z�}�I8^��+�I?z�/�=��jIA��`���n=��0;�Ӳ}1L0��G7�U��2
}�D�x)R�� m�N�7��>_�l�F؄3�
�l�4͟�543�W�r����uQ�?���T�`�v����B�D�l��	}�9Mr����X����"ҵ�QVf�\i�H��n�?r\DX��D���DnD�m������}@2����� ˮ/C����pW

�q���1�R6}�Fjc�8�
Vg�f�Y����,����^������$M�VO�x�T��<�n��G��4oֽo5xRJL�q�$��?����Ϟ��9C8ta���`�ݠ�YC��*��?�9�a+ʻa T	oZc���	:�����`��h�R+���|���P%���aaBw��:z�����#�|�Z>�C�v��>A�>J��"���֙s��#��w˫Na�C����p�8*!��qU��S<������R1[�>h�(Y��F���oD0O��^I�����*kI����n�a� R�v��i��7毚���wX d�+1>�h���D��Q��r�7mO�G����ưF"���bH$��^m�[&=��#kڨ��j����g=B ������WE����&Ҹf[�aO��RvqN,�e�/���R�݁���#x ����W\�\���U'"ky5Iu/ë���O��mЊGy>�"��ϩ��,��2�=���A�d������(��SF�(&��^�V�G ��6P;��4~c)��NΊ�6�dy�j�c�{�W�P>;�X�zB_h�w� �@Ӿ�Y��r}��ϲ��a;Ip ܢ;��8��&|���x
�PH�M�Sg��6h�ۦ̢�>��.Í�QdF�����}��UgL����pѝ1�_Ь�˲;�2�D�s��S���~a�&�������(� �t�>6r���>�SucS�}�A9fm������ 
�G���6�� �va��[�OP�j�Էv�?Yu9�.)�yZ����O�SW�p�)(�d1-Z4�Aw�c��tj���<4��A���A�����=�!訊�.p�4�`mG�3����Z3���*)d�1�W�(�%��t8�6�٢O!
��O��K�������E� V����_�������>q>\��w�d���0���v�zz��bZ8��|���'�O8r�eB���d}����I���;..�S7�fY�b���& ˭+j�wH91��$��Hb��*TVc3�!d���5U���B��@���vé����l�ÞKd]�z�c��)�<~�I0�k_�=�䖴�+�6��쟓��uw�U����7�Ƨ>'�����=�	�ia���6��JD����[�}7TyM���v��j���ϫ�cDA�������0�w-�4{~��V��ӱ�	v6���5qS��sje��Zu��'10�\v��n��Es_o-�^N�P�;��b�-`�gB�î���g�qH���Cg�F5P�0��ئ�ftD�@\'�X�- ?@��Ф�լ�fZsNB��t�����{,}��$����_���q�N7���}m=�_쏷�x%'u��[KQ�L�
v�b����#�<��j^6ѓ��e�e�UI���	�`��zs�m��(Z�2Ϋf��RI7�b�M6��s��\���W��c�΢���IB��y&�R�u�� ����ֵ�Q� �{��;�q�(��<_�K���I�E�8;�q��,�O%��dЖ*�j�:�ٍ��[�64��k`XG�wF[�W` ��B��R�B�YN�w?�Rլ%�sU�1Wk#8��	�a�pX����(��z�M����s���P_J�o��j��j?LxPg$'�SW���4%��qfJL�J�� ���8�E���l��@�Y~ɂֳu��4a�ER'0����+K�]�q��^�{�J��o+��Yq�zg8�S��Y���� -J�1���j�|:f�ZP&]�H�68���M�`/Џ�������n�;}�� ��&A������1O��俀�vD@��%n���Z�ѕ�Jg_y��,pO�������\GbGg��@�4"D�j�a�U�|�=Z[�L����ZU� ]xp���[��j,NŞ���)�A5R�S��s�q+��s�����7b��I�c��6��nL�ğ���o�Cz���O��I@�u�>����~m��4�>�]ܴ�lW�N �5?�R�:^�[�,ۧAA��Z� x�x��� �_�Ң5��&�4�o��e���:�A�|��3� 	�͢���h�hQ2
�Y��A���S�i����eC��$�)0n�S-ƨA��$
ܑ���0o/�D/2��j!
���G�!�� �H���"&,��ęPTR���*!�@(�Q�e��1ƞGp��bn��83{h�J��u�;"r41 <��%t]z����x�geb��U���Ț=C��6a��;�O<[$�Y2��q������\��Le#]�4/�%��7�~��ݣ㧧5w�HԈ����Z��wY�Z�uܬ�K�J��-Z ��`:�>]��Ø֌�N���u�0Ӌ"�O�:� |~`����~6Uz��|��������j	�3@,3��M�b�'�)�ͭ&���A�s�$�)�y�I'JM�� ��<�P85�UUA�S��]���W����(Xp �g��o?h�Tl�U��"V�����c?!Խ�7Ϸ/*�B�E]�8Ҝ8�,Wmt�3{Ե�[��y}�zב�+�f�-5�e�z��Pg��	c�p��Z���E��S�~��g����a�O�3�����D�s�D��/�}>t��Z�@Ԙ��;X3_,-pUL���|���Er���Ѩix��]������04!ԧ��wϠ��Y������]�?�Qҝ�J���vFϓ��|�/��.Ȋ�Mi-Z7��no
�@�A��Y�Yo���4�kȺm���u�qjq����a���*{y����,���l�:�&��^s|�b����R1�͢K�/���9fE�\4��;?�M���b��#�ф��% �j�(^ڀ�R9�]�� ��sL�@�x�(���x C��!?�AX//�&�ē�$���~��
re>��uuB�#H�Ui:�� �橂g��Y?)�2��!�M�&�[�A�Iݓt�[���n��<�ד��^Ӛ���e:�g��J	���9�VJW�'�Pk>�G���p$��Ϫ���ؼ��M���DK�������qr��A���
�O�����:̮��l���	������mW���Tu��F����U��7� ��p)q�9���i������"���T	>"}��T\G�q�>����p,���8k���� �YK�w}֏ߴ-,|�w{�����b��7_aU�
b��:>C��J�C�ȥ��mq�Q�#�_�V��"�R�r��Y`O|/Y6�����hZ��m�w���T=	�ݪ�?@��j��TXk�Q��Ԑ�D�KSC��-%cϯW�2��Aۆ}9�t�K�2C��E���deT3����<��)�c�����]<G��'���p �c:�'R���A�9o�y�D��b��Z�h�/ː�[���b~�4`�k\5VqJΌ;&�k�:"�1�UU~�M�U���v;�M�[�I!���˿��H���`<2oG
�s?i�G�v��ƟϮbo���ޱO$�׮��-&5$�wmOx�o2��k�/�lqoO�	:G+7H!#ms������fOV������ݧU���F�;����$A���(R�s�A'6jJ��>�7Gf�)u%�m�۸5S�;�u_�X����3+i�1� ����.n���{��e;Lj�h_�}h�O-�Z5#�\l����z[h��,T����a�!�vx�_:V���]#��e�����?��7>b��\�i<J��	p�x�$YX��LvBk��ڌنH��5�k�_z����ɼa)J9��	����ԍ�PEL	����֠�����:9��D6�CZ�8�a�J���=��UtK�p��q<�$/�>���<Z���1:�t}ڝ��ϫL$��*�w��O��E��TJi���_. c�髫���l���8��'J��%wML���P$�--��"sjO$�!��8&�}M��Y���)�������5���b�@�XЏr�	�-��`<�-�qwgנ���s�gUd��n8/9���Z
�Q>`+g-��>'�F���m�Q3+��&z+��%�P��7\5�w����-��>UO��܍y<�̶l'k�_c�?��KT6/�s\q���/�ʜs���Ŀ��y&�,��em1W�q����ղ+'��/C�n'm���#vL��@FE�-����_���z���	�-~d�j�4��)ܱ���8 ����/s0al���:o��C[Wu,ਙ/�A�Uh�ӻ��q}S�/�~��<x�]�Y�m"c��j����c��Ħ����b
�zyj��I����`��U���n��j똯_���A2�n(�C�Q��M5t6ѫ��s��.B̈́��k�e�ՕU;���0Xp�ͷQ�	�V}��v���1����S��/��}�;p�0�6�n ^5��H���W�u?�C֋�<̹ߒX���G��D�_�d�ւч�`����E~4�?�cK� 	�r�W�pV}�WW<�+�n���å����0�j���+������ߘP3����gdE���|��w�0X~o=���˅�#��R�
A�f��T/}�O�vs�
rOry�6��	v�"=�+<���W�˴h+�a7G3$�TL�I�!��	\��Q&It� �~��=?r����FVf�ZD����.�t��B��`�HxЈ\�y�d�f�E���-O.��R�����o9���]yX���:Hi��4ƂZ|�`jv�)���-��'��t`#PD����=VgY�g$����-h	�ߤ�-H�&"��C�J�,c�9�
H�rdHG�Ӯ��ҤIS�:ߑO�dWp�����5H�j]��%�Q��1xp�޼t�j��4��\C!Qb�5�f1�ݴ���h�ք2悐��ľ�\���{¿gI��^�o���|��~}!1!�ڤ�������C�X��o�^�������%�	b͏��X��j�T�j����ÙS��� ��p�ߐ�-��~5�sS	c];໷9�1Yl�Y:�9x��Qy�#H�����L�F��c����z&����vU�$�^vT��7i�=�E�q�le�w�ڛ�Y;�o}BE#�um���L@	$}j�ۅ]���Q*۱��1����j�f�����}9L�Ԗvg�U�]jo4��3iG���S%Pr�5��`(��f/�[���YqS=����3�>�:�>@�F�,��0Fv�W�3k�-+�riPZ@�T��R�]����@<�̮r�N����j#ˆ{ϔχ��0h��6C���֝b��ev�G UQF�n���^D��ܩ��)^Y�-�_�Y@ZHHsR��4�S�7�f�!]���p6�+�ԣv��'�t-'A"q�F��1�n5��2p
�����d�N�wB�Z��?��Lg�9�w�֊
����ׯ�H�}0�z)N��d'�2�����<��n���u���I��3c,��@��e�݄�sTjR$$:)q��e���<�-���>�:�U�[WL|�#�t�T�EW_�jc�Ϛ�8����[w��5�jah�N���$�Zh6�q%��X�Q����Sg�,v�d���8Љ��-��ʩd���)("��o�K�T 3[����@���!k!�臚O�x��c�=���՗�Y|��}B�n�MF#b^X���m�`�����	��'������)��?�&��\d�kl�׋�_cPX/���bB�q�@Š�~���w�M�>����濸h��)24�O{�CPt,*0h0{��*�*����N�r~5"��9(A��N��xY}{��im?�D #Bj� ��-���Bٙ,�<\6v�E�jD��j02��Hl��!=p��]?��p�O���3�&�P�k���H; H� >���ڀ�������؆����5��CU��A�Y*p�&.b=�Zt3&~���<�䫸b4�k��N���ii��W�b��+��;���0�٦��ry/��:�/��M�h�ӕ����r���!�� �f�u�W�`X%Sg���9Hg��͡�@c��~�T��ͬ�S�O�Ng��r��2����:o�y�&�p[��o�{��P��A3�s��Khc��Eg�=c&ns���X���=��;�?c�t%�ˏ,)��Vl��D�c��ٶ�)�s�0��.	���?�J<l�D�<��$r��i�X�(�͗Xe�8��t1��lﯖS��v�91�I\L�m7'�����l��]���N���
�2{6;�(0vIF�S
�tf�nb�����A�zZ��}㦥�������Kj�����F
�;��d�y�BD�S_\��&�1�q�q���O��n)ξEɮ��!շ���/@�`��'Fs3�}��e�=~H>9?��o6���Ġ��M� D�+m�#���6�0�6p����#����G���܋v#򳤌~-�R=]*F>r�mV�p�;e%���l��2�uX�Gc4C�o 42e�4�W�ʹ�`��9%(�ƤC��am]Bmoq�����yid�-�����~��]t4�$[X3{�&p����� ��ުB���B�.Kask������4SU�Q�h�A�3�!��6��
5C��A/|��^=t��{���;�>:<�4.�B#�����uE啱�:<��ab��gu�j���ȦW�\\[�.�Iq�i/E�1�o��ji5{	qچ�P�@F�Y�:��ܝ�d���ҵ1�e3��$�ф"@�xş�zZ���%�<�9n�$Pe�d^3 �@��[��d�}�)���2"U���\��l�N�5)�A<U���p�IC���Vt���C��=��ޅ�-�bB�4���V�Wȉ��¿�܊�`��S7���_�F ��[�'`X��cq�Pw.�O����p��D|F2�!����Za=$���Inb Xx�k�a8+��>��^Y�B�D]u��pR]�-#���Yy�.e�4O�jP<mZ�M���:�@b�/����s7�s<����(���[���
���O��z�2�����)�܈���&#Lw�I�Û���B�_3����m;xEek��q��/��>@qZ��y� ���X�-���l��4)8�e��װh�|���wڏ2�Xd��|��v.�
�z����E[@ht�Q��x5��"�;2lcP��ᤥ�ܜ�q���3��f �p�� 8��_w��LCSGj�_�]���٪���PR����
�i�כC�q�؜�(�p)�_Эr�-��a�6)�hvƌG5t7f⹷�`v�#hZ�J��q _ ���lCh���.�D��
QG,j�P~PCҼIP~����,������n� ތ�t6 �&��(}��k ���xcp�^���M+��Bx�e��*�@��
�W��M�G���dH�"]��]�Td��	�&�يk�����;Ym�������U��@&�5�����mEL Jʳe�}�v�O�F˧sS^	�����|� ����`!w��cK#�ia���\�Wٱx4*&s��kЦ��ҭ �v�����=:-.֡eǔ�Y���^����\��·{P�Q���=妎첫��g�תɾ<�?.��|��z�<��i��n�Gz~���9r�ܚ�@���S�� 3�4�z�`��p�L[�֜j�?�+���O���w����k~ÏxK�X��vcU ��9�w�mq��[ZA �x�)��@(����k�����$����3h�n�����e��k��9�
��V�
T8��^�.������!�$��7�ʠp,�C���2L�+�Z��p��e$�o#���?C6Ɣ�O{�������ň[���gRsDە��V>_R[�i*<rF���Q�Չo���᥉�9D�4��cV�M�hV�8����܌�U�:��]N4��a�F.��%����֨0�ɝn_5��m|�L�aWF2�f�w}�I��1��1%?���`|O"�}Gn��UZHj�Ky���`r�E�po�xbY�4��>��[�9�g~ֲ�M5i*�sF�v(�Θ����;�V[�4���ˤO�sOV%_D
S�g�&\��01�Ȗ���j�����&����E�%;ɢy}< ������+J,GR4mC3�/�WR���˯z�m����	��gfӎ��y�A.�R�"5GFW����&�T��6�)�,�r�.BE8I��=K4>ʲ.��T�輈b�Bxz���ě��h"���OSXX��7�+�a�o��v��κ����'�M�T�O�0�5��L������#a!=��P��c<����vt�yAϽGQ����C�=��Z[d��e���&����6��L��ꡲ��	��x��g#f�I�A�l�i�N��?9Z�]���m�V������& $���tuoCx��dɲ���c����s`ߙ���T��Q^��y/�&�fb��g��k7���(�g����fF�3�����3(�(� 'ʷ�?���u�����G���-ژ�RV�/L�?%)n�'��ce_�I8�M�u~�Z��!��M"D9���[���C��q��BE��m�.�;�#��קW`Z!Yh���szCN㽩F~��� _�\���^"��.�BX ����'x��5�KiI������E�39�v����P ���w?�Һ�po�Fv���Sw�l+uی�I�����<�\��EUR�����ZM���]�