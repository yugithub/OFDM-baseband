��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6>�M56�M0x��L��?��W8�tEa��d-�X�V��,��̼�zjS��)��^H1CU@
�^	d_�&nJy<���lzs�%'T�����zhQ��_�.�oG|�Yg7YJ֡�oǘ�����Ѳ�o���$'\���+O2�I����ag9�5�`��'R��0�_�����vz~�;5��E��h��pS��%fA?����{	D�o�^j�r1�y��( �:�Aa�ފx�����Q����*3��sB{E�,����b�7)�c܋_g�İ:H�����4҆���$p���f�?d9tJQ����P�5W�B�yх2h��M->`�z�Ӵ}��L�b��M��7d]�O�N��
�|L�U	O�S��삓�*���L�,�?j�����������yr0�>�A�L�eb�J@�P�_���# g�cY��_��(t�m�5�K.���2�)��;��s��Vu/�e��9\�.^ٲ��k�T�!���<5S�`�ck���7��&~�qK�Mh[T`�W��q�7�|��������7�zM��B��V���'H��)�ȕ	��������M7�ACӐ�Ig�c���5���Vq�0�c�K��'4A3��⏙S5�g*�φ�8��v�0�f����ښP246�&m9��Ch1�*@!5�x������n�����Ni�ݠqkD���Z3u�5S��h��*smcۡ�K%,W���ڧ}y�(xI�f��>�h4��KV�|<+�'���M�Vb��v���6;.���p�m#��I1�&��E����gyu�٦*��sh	���}̰���� Y���Qͣ�]{*Џ�����i��a�������`�p�����������e�\K�o�v5��d��Ll<:�;l2M2l���`@j��L���@����ʆ��B�}gy[�ӆ�=���⧎�R���%{���.ǗwϮ��� ��yM�a>(g�:������@��\��R�žR.t���|��ag�n	����,�\�=�)��v��X�%`����nF���!��"U��f6����P�=�܋`�@H���N�#W�2d>���=���^��p��^̒���i�=��4à%�4%����=�M2��dP��B��屩��t��=��%�?�P���L�e��
_� !1O�͓�vqR�;�̑�
�z,eEJ�H��֟�LrP�����x���0�zu�*�@"�g�G�s�n,9)������Ǌ�_2����c]�8!"⭛��P������AA�;�2��1��iV�C&�)������e{!�C���8Ǡ.S���\Gu�p�_��t��yH���!T#=!p-�冸�b#�~6lG�5�z^�Z�����c��M��4�s(����G��o�х� �Q�h3�c�n	Z~���7~��˝K�0;�I@a02X)M�;6�� �K10�_T�3�ѻ��"#�C�'B���5zU��:do�,^�\j$��00.��*���L	�}�*7}��L���]~H1d)br�%ܗ�����\�h�ף,Uؗ��,��<Ә��[�w��b���bpf�#�Z��6��Q�i����B�C���b��z��3��s�	��B��8��~�����U�%k����9��6㉒��-�ab˾��)�߻�
>��GO�������[#��Z������=�w[ig�0�QM�3�"�]�eo�|hXԭȠ�Ix�����-���թ���&�j��>����U����x[H[��Z�����7����+r}M�|_�+>' �2�U��ӗ�����<��VU��|�|��mCW��m�0�.��?ʾz�3>8(�L߳�֯\��X#�<�:�s�e��'�٫z�7�f�Tm��n�4� j��/�b�n2�g��};@��&mˮh�!(�ȟB�j��\�3!.U�y���ZC��,��v�f7U�C)�^
u��~���Ur�c��3�T�q���X�K/^Ϲ7^|6�i�X��h�F����K�ɻ$��Ik~3�O/g����>W��I�6��.����~ �j����u���i�[Eb���K��Vkhպ�I8�=_3\�-��Ći�3h?��{��?ƹ1s����`�E�Ǿ���ތv�j9
��dC��Ơ���H���A����Af�C�L�$�\ؼ�2��Yɏa	X��7�;;���F�z���7��[C,�'�Z��Y.-d�&P�Hku,P7�&A�3%�9�|Ѣ�8� �-F_��_�����T^�{��B۪�cKT�.���ؔ��.��-�7>�1Ƭ�9���)+v����w����n���N#Ɛ\Yte�<{�w���>U��-���t`˦Ns�G�OXxt�V(�0yY���J���%���ΥH`Q�0�M��:.K/1f��O��Q�1�r�D���.,�'(�Y\��.!�;GG�/|�p%ZZ5J��Goz����+�y��Z2ͻl��1�]f�O�tT��pQ(g�����5۲&
꾨�R{�nY�t�-�aa��0���W���~�M8���hd����j\?x	�d��eB�]�O���C<SBbP��[�F��W��Zp7@cA|ʏ�|0y�������y����d��A]��8M%�P��o{q휓�����)��4�o�P�C��5�w��-���ǳ,��.�Eg)o84X� �~c�X�g �� q����&�P�-8�=)=D����qF%7/0�Jp(�{��L�0���ͥ�d�:"��v�a��o%��(F�|n2#�w2��lܞ�cdTHu�ٙf^ՅPզ�!��yA�K��r����7F2�E����a	�h���y�
��|�´,"@��Ϊ����hH�a,�S}�'���[�´�F�c��� $3~��ހ�r,���`�Gј]�_W�J�+xX�B�S8rZ�vk��¹�N�Ȭ8�8�9�bi�<��@@*� O��cy�����-�m((`D��p`�3����A'�n�8��W�9?����[ʖ=�p� ���%l�����?�>�KO0���D@UGkt�䅫t�+�4f�7��2(��X�:�}�슝�$�k�/��Λ�= 1�'~��oc��գb֨ �w���?"�h���b������A��?[&�^��~�g\�<Pd���̟��-���./}� �ah����q�P1�������gJ䡞, �1`�V�~�A�J���;-�aK�ar��0I��ltr�K��!w�5X��r��EDQ���-�E�I41��?4$ɿD&���b"��E<��P�w���1�j\$=2|9;�4;�.���&fiƒi�y'7]Q���	A�H�yT�E�;��rZQ��|͋~~jAم|ć�����E�2)�C��˦p�迓��@��$��^)������!羜+g!�!_��,'���^u�}�R��y�
Nhj��#�^;��3�r���G��i��y���-_dW��wB4�٠�=:���P������\�$筟�5t,�;�!W#�W��)��t��B��Tz�MT �����R!�j���?BJT7��������Z	k2�>�� �g����b'^e���&SV2�F��"*�2q�x��U�����֌�H]�l#�bg6�u~�7��M��♌��?[���-{V�T;��pFI }g�X��4�r�g�g�~����;a�m��yeq�7��WF.��z���{�[:f�ZZ��E_Ru���`Z�Qa�u�Ҁ�@��0���?yj��2�i���ʲ����~君=Y��3�M#���)��#�P�yZ0�Ė6��6��9!�	vɣɭ8�@�����$�Qi?��r������)co�����{����7���/Y�*�ǥ�����P� ��8}F�y�B�)A���T����:E�}�1��EH�[�>^�ŋ"ڨ�tz�h~s
�K�X��a:u/�:�@��e��F�5�혬�d�-5�|���u�Р�UK_9}L��vIz'���l���v��
Ǣ��n�j�8�7�ن.��*��cP9oD��?(��<�X�3�G�,O|��x�s �5�b�Z�5��ԯ��.�-Z5�q���
�د�w/g��g�aፔe0pUO��?���aC�Wlu��)���g���dC1�"���-��hg|��n�֐�aa�|R�yC汲z�2E���*�K+(� ��090��]�4���~����RH6�����:A�ҋ��bQ����$'1@��f�� �/&M$�p�6|�$߸���Ѩ��PB9#�4+�L�e���8�\���Pb$�8�XИ�u��A�5��~WL_��ߣbkb%�������߫���X1Tve ^��5�ț��x�����[d����odj����}��Y�L��BX�IGX8�����*�"�Syj��d�--�w�sg]�
)ḁ^��R�g�q�Lb'z�M:�}�/���-��(�*�-SR�-�yMz�&d׬� *��Id�6���	:R� (W2�a�E�`	��
[��E�3M9�D��0Hx����lkkָ�t�Q����V��EmF�s���߯_��|�qz �� O�t<�cl��l�L�g̠��M&U4(J5!�T�Ja�������9��Gr��M��������_���v��(N?���x��wӯ��|��O~Z�T�3s��I�}��X�����gw%'��G���Ͼ<�_�;?-j6ǅ}�+o7'� A� W-K��������
G��Z���g��:��>���<���!���(�#���Zڀ�!J�4���Ҽ�yX��ͩ�M�d�ܺ�2��F\�i�ٓ�\��~rS(�^Π�{��Es�\�ҿ
V䰏&�(��s}> ��+��Y���	��-��iz���t:a � ^Z�ҁ\���2�BB� ��p��^�� ��q��$�Y!2ޚI߱��\�ҕk�l�pr���L4sx�N��%wF�!s#�.F�k��~����t�j3b�d�J�G�pU89�	w�ǻ�>Z�W�N��y�C��[�P���6�����]mBT���r;`š�A�ñ�Nv����\�i>�
��c�������wEh�|^Σ������l��e��`�wTx��q�3uq��O�����Ca�u�d;�/����C�1E�1�V�u��XH�;Q9l�!y��?��7�cK#f֍Mr�}�Q��Qh�L38T��xJ���{f{� �����b���{��~�P��ӬH�m=�t���=�{E���l�X��(i�T�ӵ�~�9Q��^ܝ��fe��ko�j��Η�OF��� ��D���R�0�_ɿ�B�;8�(%ю
@(DJg{�#J��m�.��$��[s�E�V�lM�n�w���{���~����H?	
���r{�\Ab�q�TmsX�q�hD7sdE�/:]2n���v緇�O���шm�m��&�Ԝ�-ߺ��1]�p�05���s�;=G�ĥ����Z2�_�[U�=1�Uڞ!�L���!E��n�.�B��_r�zT�봧+8a���u:�L-%@��)��]�8 "�-�^k[(����XJ`ăQ�1ޕ��R;����*�$�.��oؙ�"
D��1�D(;�$��qO���pwy�E-o�`��&U�N��$�s1��#]
��oW~�y�ʒU��� ��w*���P�e�e,��_3�[V��2�vZ�a�8��� :n{x�-�`������p���NZ:2	ot'n�bFf�`������'�m�h��q��� ��Q��T�ş�b�,b���ƓV"��8�I����{�O�t 2���t�خ�Ɵ�P��j����k]��A���-Ez���dE�1Gk�<��>)G��齷m��M�a�|�3�N�#�Nԍ�-}"�W�2�}��*���R�*ڏ��qH�1C��
���]�Ę���Ё7�6@7*����f�����bS��T�W]�̰�A�U���+�ݐ X_�aL��_e��Ċ�]���S5�i����' 4��X�{L�&�Sl2��p�Ɵ]��̓�Cs�bZIЂѧB�ĺ� '1I��Ǝ��-�1s��B�q_�eZ辨��a���Z#w,7cxo�y̩�BO8
"
�KB���?1_����m!]\�r���Uq�Yľ�zQP�i_nLG�6���$z�WǾ0rh��[�J3�*'N�U	V6�xXq�����!`���'�|&S�O+:���&z<{A�i|ϫ��[5�J�d����$O2A+M����ה��-6wX �8��F��#�~~�[G+��W	�/ّI�)��q`�W=R˱L=�pPn����M~����v�FP����hR��R�e��$�{�!��x���9�Z	mQP�&tr�]V��܏g	^N��h��^��<h�boEX<�	 ���ry7���v�'J�ּԍ���dh�N*�(���S����r�R����ٿ���o���V�����.j�P��%�(�h�7����g"YT$K��.��8Q ��0����3�����X��J�BT�e}#����?�P��1�s�}���ni����#�Ga����V�0;�=F��q��ܞ
�|<<e�v=}��5��2���9R��~�b;�+���=u�����(�gQK���Շ��A�A�^������7/2��-*�>�i�s�4�X�j'�@�}�	\_�~�?z�{BU׮� �^�,���ê��@����E��#���^hԊ[�?��|ClMU�NxV�	P�!b�B#��Q;�蘜v�����W������aq0�f���,���X�!��f�萟�1r�iV'���V�����EW�R��f�9��2�u�-q�f�xJ���S*�8�ϛB$i��蚽(=Gl��5�F�sot^��kX�!�{�>zy	W|��l��}�W��?��eD��8�/ ���]��T�.�5�
R�.l��֌���N���6Q����+���S7#g�m�	K�`�]�; �_��^�L?��e=т�t
~:�ITV?*���؎�ݩ�Y��-%��b��p�D8�'��hi:�/k�I
�N�0�W�
g�T����7�6{���=��]�P�3~+�<tS�]O�[��,bG�Yb���� >�����i67���Ad\�鵓�w�܂EK14K&�=��}�K�=yE(��D��~�C筑a��	����ĬD�u�j�\��p*5��^�ո��$bK6M��(����3}~�+i�,Q`��%,��Nh\�I��Dw�nx�ʫK��zg˫^����X�����$���o��;(zq{h�(9T�\���N�_�id6B��~{�'�Z����#86�E�h�˝�@���]�y�]�-�.hE;����&v�7�k3c��qH��}La�HJ/�ܹ�3n��J�gq`���j���?�@@ȕ!�w��bȀ�{���r22Uc��#�wl�2ɥ\��U���QV��Gd`�aLg~����ƫ�z<�F�śt��8���M�)m��.�W
RP�2�Y�ũ�B���ij-�U��f\�6����7�NaI�B�G�aw�}8�񾜁*��%��!|�������H�5�#���#��9������s�.;E������x+ؖ�MQ1H��C��C�x;u������a/՛��y�
rȂ�3u"[1�4�}�{�����+h�?>SPXKL���.�P��J�ԟ���%�*ơ'#8�s��L�^�R��,�ʙu��_��׋;�ڥ�
�����t�Qٟ�$'����$H����o�a�q��tA���B�nX#�Nᘽ�ؾL	���>vz	!�Q��&RY��6�(:�
�)!�9O�=���R�9��Qo^���g{��GkH�(q�-˯�yIP�Ik�,c��4�N�������M�AH8�W��}�ڲ%�3��,_�:����82�'���������������B+��g���*~��������x��6��YV�	��}���KX($Hv��\��_�چ�����v��)6�ό/����/*�,J�w�@>���1��O�h�S3D�( �9l�2g�;N�CC3A���r�)�Bt�<�ɖ\CK�o,�9��K��o���w�4�"��YG�5E�k��w?�[�͞�:F�XEyA�������'�@)��.���� �9�%����_�!�K=z�n`��ık����� `\�o�֗j...�f�������A��Q>�ǩ�y;���h���oe�r4��QI��\z����3>ح 	��~�Éa����|Ơ���E�F��.���c�3�	�Jj���d<��܋�˚�M� A�>�F���z�-�e��P"J֬�f3(w<15.�K�����L�c�G����e��S��v���ZBv:;��q8T挥����<���D�15�ܪ�N~֪dVI���z�5̓z�~`�.��W@�