��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ��v�2T�(S�ư������K�_��K�qu�7�7*dg�3Qy��O���T��71�"�Kgo�!�av��C������o]��lRg�Iu��ߝ�[�%>��D����o�|6p�1S�5�[ �)LA���ː��>���-o�h�q��'^�7�O�Z������� �[l[@F���v+�u����M�;�Pܖܱ��C����9*#�ه���:rSŝhGRġv�L��\�^Kݺ.�Tu�C���#�I@ .�G�x�5C ���r^`���o�o
�^QP��.�����i=�������zi��K<S�S�,��.|�<%L�բ�+�@�T���-���h���@)&'�����4Ϲ_呮ˌ��eD�'�9�CO���D�g��C�%ՙ	��Cg���`%��q�F�J<S�?Qt�Ҝ�/G�f��?Ƈ�+Y��H|��Q#��!�v��_��������������@\9��4D�4g)��V�r�0u�Z�s}��يcIsI�����������[�[<�*���B���;~zhi㟚U<\�* K�.\�ſW<��b��Q<s<4y���D.�P`��o �*�~�%E2g�m�c���jS�'Y81��6Q��x1$��C�&Mw�ic+	%V��>LSM͚|c����A�M!��ƒ���,�0�D Z�0zzù��7��@�U ��'����� ��T輫ܮgS;�9v9�s8�X{:�Hϣ�{��ڠi<m�{�h�3S@���t��N���yj���.��ωzͼ͙eidw�1����u$RO9�Sj���0�<�.��m.�-��+I�n]]|��H �K��a�Ţ����=����_��}�¼�C��:|�a
��=��g��ٰ;HU��,�Ɂj͖|h���`h�:ȷwWP�3�����^-{+C�5����E�4��Pӄ��6%l1�����` ת��I������u4N��:D�׈Q��b �H� �Ϯq/�1����E"�C�����
htB�_v�pV�R�0��똞�$	�Lht1��L�5U��>mC����͙ �'ja� m��-6��T)�J*xj?�^��t��ݝ��Rk�gD�֋��>�Y+T��+�RiOl�`M�h�� X��WT	���W����<|>s��^R�2���� �~��F�%�A���H�������I�a"U�s˰Ja�����}��ifd��l�{T�<��՜�1@�ʙ�Xh��C�_X�-�k..�ڜ��g����>��,�
��9�8�AD�%UMM�f�m.c;0����>uN��3[Rp�(�V�2��t앲��R��.h�ɿ��]xK�+�ETL���Y�@��X�z�������ߟn+��`����3�S5��;"Ig��_�D��k.��rry���qq��E��!u�*���|G�P�Ʉ�m�0Yr	Wmo[�i�g?��S`d�A{O�,ҧ�~�B�[&�?m��3}oK�J�F�_�_�������ƥ3Ā!�]�}��@���D�鳳18Ypԑ�)eÈa	�?L��(��s{�ct��oOH��u7Z��zX�qܐ�Kq���7�e��� %�����'�.v�z׏�Yf��3WY��߅���|�'����GBs1�o�^W�J��&?�K{�-aB1�^2� ��)T#],/å�44r�{2�7թ�I$\s�>AXO��C9����K$�N�f������V���v��\��cP�N����MF��b~�r���R�F:���:�j"�pt�	��G;��#^4(��h���}�� }I�˕��tb+�O�#|���`BԬ9!V�Wv��Q�ޠ�õ�NB:iL���Xrp��EH;�v��C��J���'�a�s����R�F��1�H�)n�?5XN�2)q���j�ȝ�7���}�}��dk� �`X]%P��_t*e�G�*sG�����8&�,���6��(�H}�	��0�5�@���<�/W��;^��#Q`9���?�BV�=n
����?�4\ե���gk5�:K�"�쵉1��I�����|�U�8@d.p/i��M$�0MC�W�I|m�WG��W�]D���)�8\��=���z*� &���w��ǟ�J�d������iPG����}�G{��?��;W�N�Fz�'����RH)&�1�Xxg 	!Ϟ�4g��t�SSMr![��7�7��1�e+�'4�$�JŔnq(+}f�gm��ԍ��6w�X���4��щXt�����[i�[���~�pl.��/��e���{�����1�����?����vj	i�C�Է�YB5j�UHX9��W����SL�m��t��ا�{�=Dc1�*����ڴ�&�]���h�E"�ú �x�B�BS�&-f�\�UɥG�1��y�]C1��*�
�G(����#oD�1��y'CF�>�cK���Fx��/�a���)� :�dH!i��sa�l�+J/z(3�Bt�(w�s4"L�-Ye�-�����K1=�ϝ7�k9)G�Up�۽>��⍞��.m�%��x	�Č#��t�"���!�t��'`�#�c��n{�Ȑ��.Ft�*'�r�k����f��f����O�ߟF���ܬ���3�����O��7���KВk&�c�ꧠ�L�`�}����}P��-�?��,_�W��(��7j�/x[U�p�!�g3��Jt
�lh<�t�$����.� �h��_��5�u>�h�
�d�y�mG?K�P��'}�-�C	j�,�j�SO���ay�by����0w�xٳL�y����C���n�m1�2F�1o��k�#��K��o
��� 8� E�J����;|i@�8<���$�5+��64a�zH�$��)T>��Vφ�nFܥA�I�_^V;�mR;�ț��yz,kX��KLZR�����U^�x����|�-m�dݬ�o��z��0je�nm#��C5{�+�N���rJ���BR�Z��{^U��wk�q�&	=^������y'������8��SC�F.l���*�E'Z~!bPc�_UԜ�dB�0�H�֘9���v2V3d ���Es�X�������N��[j���b	�1��
����F�̦���I0㵄4Mů������-ގ�e�@���ip�@��J�b�H����A�4D�+pK�L"�W����>��@ս�ZB�6a�zĦG2�g�gK�v���gY%�o�s�	M�CD@��bz�]S�;Q =��yk-z.��Wm��G���l��2J�[����W^�WP7DPQX���6�P�-�)�U�h��x�Ƴ�Zc�`"o
�5W�	�&�=9Z�iߨ���t(-*��P�P�/Hl_�x� '�	���K�O-@��e�R��@PN�.x��w���Ʃ�qM?���幑_���ɍ0��B���L��(�4���x�!@V�X����*1~|�r5y��F�3�_�i�F�<;)��pN��H6u��W�$.}E��w��S�G5C8H�3�6�����\���0|,� �C�m��i�4�g4���^���!��P� H���!Ȓ>��>�|2�b1����B����*�O0�>0�¶�}�Q}�$���t^��>Z)��|��"�*~���C����6oMD�S���P���v&5�2@������eMr�G��G���ӿ��r�[k��{C�����-a-.g�U��&��#����+���*XI��f@M�;��sp� ,��VK����Ap�F6�u��-}����]4p�NΗ��M�n}��~����N��p��R���BIf�:�^��Г��0nѫ��}��P���:^�g��%�EN��l�乬|�[�p��|��ȕGt`��ؚj��Z��'-��I�i>4�����g��\���% H�/ƿ2�w�c����%�H#�����_���Ī���0C+f)�G�h�M�Rvu���/F�����h����0.D�译g�W�p�����\�b���s�UV�1��g}}c�\����c*��ۧ7�a��p.bJ$OP��	-�Fy�}���!B2�X_J�O�;��/i	�*dU#nr<�Y����[�eY4��
�Nf��,�����.�\���2 �u%;�\�@w���W{�C3�A�5�3^Px�o0	�~&�rI�T�j3�[��/���"6ڕ��x��m�0���^�.e3��~v�O�L)�uc������-����R�?s9>�L��N`�z���LO�������m���O� ��Ri��X��=�� sz3=ϗx�X��ʋX�mr�^
�&nݗj)��ߛ�p����<9�=B&L��p�Ғz<�1�1�ƴ炕c�Z�ƨ�x_O���)'Jգ���k� �fK;�e�]%M	JNq���а� �@�;D��S�w@�ŋX[}��k�wfv����G�OtV��~�ȿ�_�d|N.h*Z��Z!0L@!t�M8)�xGN����{�|�T��+���FJ�X�7��J;B,.R�[����Qm�^�kRqr#����D��QPm��9����Q.z�9�� Zt�Fa(�ht�(Bf���-�[���XM�B�j��+ ��9��Ly���T7ܕ��щ ��8a�$�ʈT����#���S�_)qnB��|%�зᇟ,�{OC	�����[zR5�ف";WcY��DlX�%t���B�EҡR� h��[ѽ�i�c�Ti5��d�on�X��?����dOd�Q�}��b�q~�bkPF�|������>T7z*vCe�"��%�>bы�T���ƺ�+,�?���J-��l.��¥���/W�ѧZj�_���Ώ52-�ŮA��~��1�Hg���_a�n�|�P�8���K�Fq���V�=R�����=0ޑ��h�~���Yu#�)�:�x�F��n�#�l�ײ�=�I���������B�vA&(�6__߷ćQ6�]�ʂ9Ը�:�hO��꼥tQ��J#��+�"�q�v��R��Ow_� 7�tk��d����)@�ss��ٙ���W�JM��~NC�C�₯Ъ��l�A�p~�/p}3�>��Û����a�G6�ײ���4>�dn�,�x�c�k�Ul@�"Z�t�y��Ȱ��s1�`/�������I\w���)�p��fӚ;<��s�7�*�j����z��몮r��^&�7�F�v�B8yB@�_c��Lh�x��-�����$x�u
]z��)��V3lί_2Y�~��dkA��[&l�i�j2/�!Bc�������`-70<b���'M����H��i��|�AY<j�?��g�@8U��ɒOl={0�ڛE�B:j�|{�M��p[s�:)��'>��$�NO;��>�@n9�I��v��ݠ�fV�4l�s`�5I�
�i7y�~_)ݷh峛E��m�|6�$��;`.�����6�/ޚTἾs�n;{	�"ia0rp��V�m��p7�s�#��N#
���;��[����#�T*�Y�A����8@�68(�Cz7����
�~�a]x^�Ǭ�)2�b�r5��6.p�:_���7Ǻ�[�Ǉ�`y<�#�Z�Eī�z�	�t�Ioi-�^����R�����Uy*��{�C�Iu�B�'s`�r���M��#7�|z�Ghk��MxO0����oq���w9�fկqgm'���,����d�k�_�Qc*(G*�{=$�������ԍ�a�Á�`7��Sg(������x����h@ е��N��$�\����&�l�E]�'l@�����1�H���-qw�k�͘�YrG�ƷԹP�C��/#Y%g$�.[~鷊<Tl?����H�H8� �i�{��ފ����o�rf�����,s�j;?H�mN.d��W��@�q���u���q{`�{<b�B ��4~���H̺�c�F��#喇C �0���1�c�V�f���x�ٰ/�dd��0Z����>��F[q�ek3��������j�݈!B8"lK�!L1�!��o1�a��
xD�eH�=�܀%3&���!eb���w�;�?��0=�������-�i�kwIP'��jz=f\�m&��I�V�����t��2l�|��M7Xtq��9|�^�dD��b��L�v-���$h��	P|2A�I���[��և)����Ij����hG�J����P��p�*�b��i�P���O�6��j�������%�J�A���J����m1,+�gA?K��nߎӺY�K��8I=oP�<&��@����ט~���;K��Rh���`!�R/C�4�@n���q���¦����)�"�+�2, [���8%��5��mV�]l���t��Gl�%�N�����c�m�V��lf�?��鮁M�=���^���7�ƤWW 92舥�g ��B4�C9^��?�J�3������h�ҳk��MF�*���EX w���E��["QM�,��������$8w���^���?X�C���i�I��L,6�a(�k� [��P+�������-��J��/���ajx.�n��X�\d}���Zz!5�a})�Ik�ou���?k��	�Y\�1�xޛ��l�We��櫜�<��B�ĥ�&<�w8�]6
�N�f�T�r~���J��K���� Z����̛�KP�(V����.�7V�>��?d������4T�k1%�X�3��ޥ��8ϰ��� 1�����j��j�6o���]r1��N�޻�]���)4�����̨sb��E���m���S�⅁��TA��.�7�*��s]C���ci ��g�6�,o;�AZ7^�S��-Mj�c��زظ�,~ ���O�/t����?�2��/�z��{�؃Q�ł ��'� ���_ātRB��0 :/</��4�Z�q�S���kK��)�1�4+��x����	a��i<I��[�_qX^�,��WG�%2���E��綅M�����P*�������fK�v�x.�𧒮K 1,9��+�mi���w�0��b��J����Z`#����Ŭ��o��Z��ATt��&?@�)���?CO
�Z�)R���q�Z.�[������L=
�5��)�A�K,�,>gѫ�y<`k����#����F���
�T�e_�T��	j������H�
y1`�/r�׵��Irn��ԿO��a�,	G��ۋ@�w���H�b�T�Af���ڔ�(��s,E:�伆�"�"�G�~��_o`��n�:J���9��i:�� ;g��Hmy@+�hy���9Go�Z���*�Ooas��J���B�B�,�k�e���E�^θ�g��D����g�f��!�v����c�p�^��t�Xf���1���+�C�?%�);!�A�j&�?�6v��)�6��4E���1u�m/�-�N���'���/8 ��_�[�S�Ah�~����jg��>؆R��tW�k:^h"�~C�P.Q!��j��7�`tZ���~�=	?��L��5���Z�Rj�UT,	A��#������XA� ���)�A5��D�M�	U�v3��]�7�
�j�n�ާa�vU�ȼ��3H) j9|���_8c�~���~I���xH�e��� m+З��lO�4f1�
���Ʋ�E�A�B#g
�����)�����:݅�l��=7��h �g����i]�8yT�$������fd�2�?�߃��r��rVG���P,UdX.R��������E���*B����Ę�Xk3鏿�O��ʎ;=���kR1'�
nn�Hl�8{��~�������v_3l+�f* �i�t�a�xaCŢ�.CH���[��l	����й�(�L>J�+#0���c��])6T�ń��3�Ď�7�n���5�
[��
?5��GM&*����Q�0��e���3�IX���v�I�#G����ׯ�bjs��
�ԃ@HU��2���ݴ��-x���$*-����x�2�N@�O�%�MT����<��F����aG��%>O@6li ��yDQ�i���R?����Z�0X_U�����C���������9:t�����e9���'��1=�ݒz�N��*_.���$qd)Y�/Utѧ���Q��N��A�����i�� �Xw06O5Gg�d f�47���`m/�Lo!��G*���D����Oㄽ�{pz��E���ٲt��c���%�NP�ز3wF�	���M�y�:���YEF�omb6H^���5�*�#u�wLo'rq�ͤ��;�Wr9��[���Md̣F��BW_�zXCYK��}����Y�΃^����h�8%��#a�,
�Kx��]�u�_X
ˊ{�2Pm^��޽zs3�¹˷m�����|pdZ���T�k�{rs=�8�>��;%jo�Xv.������:�g�0Ji͑�oV���<q��N�j��	Ņ�vqQ�Ƶ%�Cn:s�QKǔ[�{�)5�.�|����T��R*!�Ok��JPݶ�-��%4�|�c��%p���2��M3��"R�/`�mW�D�	F������s��<*�b6x�S!��-��yE���-��2�3�àQ(�������m쒕,be��Jk��ʱB�o���e_L�^i�VHb��2A���I��0}P{��>8&�<��v.-ѝ\U������j���"��f�@�3�?@mPk��q{z�n��M����<��S���r�VLIَ?�6��y���M��6�p�
�6�)e��#���F#
B��{�@> )k�|��-��ǁ�N�!}j㦍�g����4x:լQzRk�"�5�	�e�U�#�� 9��3� �ұތ�Z�CyS�S~���a�+��?�����l�K��[U��ƶ����ĝv�:;X��?m{�}�8*v���t��$dy���38��@�O6�-�*�-R� 
ڌ�9�! ��X�7���^ې�>6/S��͚���kDd)�7}]�qk��}��T���Y�2"@�q��AG��ّ`����w�z���~{ �3B/'=�Q��c��muq�8[������5z�3�4i��}��/�y�3����>�� �ɦ�S=�ys����W��IR�O�9���jFPhD9���X��Nr�ݬ9I���"� ���zj��&F�~��}��Dq�����}��L�Y�+�����EL¢*�-Bt����Hb���6���=Ai�x�c���A)+�t;�B��N�G�8s�T:���O}�Eԣl`��XD+���C�7	j�R��}����9BM������d#�ʝ3��)=B�<nD�|��!�;��#��j��ӌ����$��1���Q��]����E�bμ}�y�"6�(רV�2d%jHf����&��b{E)m�\6�/sR�Z��������QD�<R�@�����������"�����^ɐ3<=)��V~2^~�j���z]�e�S z�n6$�D��F�@��v�̃��c��]��x��"����E�����<Mݛq}�a���;@O��@١��(ѕ��׃�7[�>˩tY�~�T�Y(���G�<�������yfx���%-q.,ϝ���G���$dW�tũ�v�����
o۽���PL)�_���� ��#Y�ω�$K��-i����-����J�����<����o��=pJ��E���h'�Hx�!����m�Sk���V\1?;"�����(�o-�8<^�*&� ���}�"w��D�F�ZA	�<�}�m�Ĺ[�j�S�� Ci��I���I���޲&��6�)����I�|.tvA?�U��u���r�{!z�����i������f��&����zj�=O�_� ��o�����j�8��o��{�N?�lVYhڏ�m�g#�A
�'4E{��)�RHk�^����m'����/	
��04.����n7G�H�j����kX5��X��[��jKN��e�o��|{R�\�e�����X���P��I�a�v9���V�7��?6��Z�M�0�!�G�����4Kꊞ� ;Ѽ	m����,2�m�F�S�^��m*�L�S���ϖ�ɒԿ��n�Ek�L(M�7���+�/A�5�A����G��䄣���RT#I-�]��-;��zR�bA6�9�F���bYS �F�0s�,�O(m�i���^�SN�d�J)2_	���*s'�M␣�� 8_�٣01�d��հ� -kҌB��2\6�H�@3�N��?Ov��:Y`|���F�,1v�0����4��J�2f�(�=6�pB,řg���o'���4�֋�Rҍ�2]̕�ey朎Gb�t�rM7N��r����p����K�:  ሜEZ��0/h� ͩdGz
�iCr�S�@�[��I"D�b�YŽ|���uv��냽���]&r��7P[���>�%�}C�,�eX��O�
T�:>�1dV��]\JGA��M�eFpO���@�n�>˴�]��B+��£�̅�