��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�����X�V�W ��t�6�p:�Bc�B�Aj��
�J3zv�K)�`�ݾ���<Rh)*Q��+�[wB����������vY���ôn�R�O�%w��
'̟.�D������Ӎ����&E����G�;r�$"��n�p}rv��T;�[9��/>2����|ը~�]����a��P�Ǧq��(�d�	�O��ٗ}�^�?�FʹB]����A���k9��.K.�VU��筜W�0XK4$���o,�d�G�ϱ*�J���"�!^��i�WpA���Y�S�p�C�B���r^��	
.P�kCf4�ߞb�*$�մH����_i���
t��(g2�L����!10��k�P��E{�䛺O��en(��z����ވ|���&s��l��M,q�f�M�>wN7:F���X�K�p(S"3�R��t�󒽃���M`p���jL�L�֔Bɽ~+һ��8`�%+:�?�����-a�e�.Hxc�������+��K!b���;KKp<x����2~�D��;"��-�ota��Q�����[)�-�x���q�	�o�["��=w+�*~���p.c������a�����Q�tdK�5^ً9�0��8�b3��4�ɺ���n�\eK�V|7vi�b����	N��4��Y>Hn3>�0�B�q:E���G�t<����8��篠�Dҩ������G����Z6�V~�U}�b���ԣM�χ��P�H�x�ڤ��T�g�G�5��E9k�A
XlH�g��2d$�?'L�v�)�c���J�Z�Y��8~_���,��������9�ؔ2����@9�Ϻ����a�<�0����y
(���SЫ�.�Q�M�5	����#��<ˢ.�AoAV(�2˯���*��=GAKg�j��Uh_;�H�ަ)�۔S�Q5� @�PN�w�cf��?����{d����޹���_̒Iz}L_܊s��-��nXc����Y�w;�v&`Y��]��uq���[Y��է<+f+�f����^X�����-����}�������rb�O�o�t<(��
K���{$wG�smf���+hE�8����G�f��@�9�Х$b��ϳ]}�)4�w[6[o`�sB>��Sʏ�+�>F� �N�g^�+��fƬ"�V��b��� <�gV��F�s��Q���>͙����@�+�D��V˩�����(`rܗڮ֌u���q�/!m�����T%�Ȏ8t�w��Z�/ಝ��z�3��u���#���i
*;���������8;��T�V&��F�5H�׫���~�+���@`6�⽽��%"NTD;!�(s�6*@]NoR߿,,�d(�T���"H�3qy0)Q��I�{t�'h�USa����J�RT	����8u�?
���gDW[z��@|��ϐ�m~�@���z���G��Fg��2'����yo������۪er`-��ŀ�����W;eO�둡}ʳ���
�G�jW!=9�6/���,a�0�~��V��ǔ�[R��ҕ��u���i`+�s��W�sqjO�n3\tE�-ގ<�#����G�MC���vc��5�m�X6��!��z�O��Z5{͗���=�Z'Y�-F���?C��yN�cPԘ�3p����&79D^vrh0��X��Ϟ2��R�lR㣥T�R'��n�.������a�K���go�eV���kM��U0�Iq��`���C�����G�ս����o��j�HD��ᨽ�3"
���h����j�'�v!�Pc�cR�z.����AV--�L���\R�Ҏ��j���h;�3�G��{��gV�����=����%`"���Y��9O�[yv�A�{�d�c:�G���z�d���*�q��X���aO���X=�!A�G�D���t`Llf��{w!r{���B}r���M���*�ӂ��xD�[�/���.�A���2�<���<���f�����Rb}���U_\�r� \��}_8�ɴ���rЌ��%�$6��oO�Ŷ,u��ΉVG�>_	���ba<I��M�����"�3�X�Ƴ�.�a���.���Jp���(��`.D���B�$��#7	�$�[�:�l�#��-�Y	���e���b4�h�>�F���@��3A��h����;��݋�RBt�"[��|Y�T���z,&(_W'�ٳ=-x�����?|�o4-Mj��l�n��]HY7)C��������UP0�%b`���<30���Yz�1�0Y��t�=�ƶBH�MtT�6�1�]PGw$Hl��®��8'�W���?�1��<Y� ����}���ǫ��gc8OK5�O�=TJ ����l�h:?|K�utP'}e>1[/'�]hK[-��K�FEFxͩ\��tF�:�35}��J�F:*Abpq,��K�n�)-5�.ɏ#�o;Z��,�0zi��.���8Z݅Y���Y�o��MR��ys�7D.�Ag�lޠ� R�7^5��jñ[�]
E:Cb�E	o�~��X.C���f�w��$��ȝ�!thv�&t�$�8�eP���nd,����OΒC�+tKfg��m��[��荥�D�{�
����Y��|4����M[�]��2#��d��(L!2<^����y�;?撊-�E0�b}56�S�/��+$.�4��L����M��C�ZQ�';ٶ0JьO�-���'JLq#�k��Ƭ/q^����/�ʕ��|M`�?������M��U��)���֛
�Z��j	��oa��@Lxs*���-��T�?�%�x<T�)�v��9�,2A��/���T�)[�	�#N�뱪Q��,���ށ���O����'OM�⬠b�U�4����S�,a��Z��&��(����4��@�Zpri"��"�
��M�эćG�1��ÿ4��S<�h���i|����D�<[\8S����L>Z��^���-TٵA/�їU�����T,�xc AX�_�~.D��_|bͿ"����w�#���(�";RS@:	��:Ph�H�33k��/�W �H)Kk{H�Voܫ�<�����DZKW���A���w����+ғ�mV.Tu��b��)��jsۂN�ޟ���|�3��jz::��*ڳ��	��w*��W$d����vf���j?�� �f4��'u��]��2�+i����Jh����Oeaz(�D�i6Ѹo�#��YV�x�F�ӣ>�Ԩ�ȥle]r��%����iR��!=H�c-��^{O��VȜ�Ve��Q/`�Cz1����KY���'�H�+�ۗ�෗zc�a(& ����
%מ��k}�J��i��䟧�,�5��4��A�w����"���.����\H�ryL/I�K�9��h�<L�,dG�������/�{�wm�M7w�53��ЀӐ?��91�d��U�Y|��T�d����7�;��P��d�SEN���	;+k+�v� ��i6"[;����Fj��ڶ8^GEC��|s��x͈��Pg�"���\�W[�>¤2S���<�7�ʝ�����:'�t�YeFc��|��0&
WK�~��3�%��]���W�X�#�v��ZQ��D�Ya�r�	
��_�E�8�B(�}]o��]1��?Yq�ls*8͞��u�7��^���7���l�P���VC|o��̃M>ÊD��P��3$�3$���;V9��^0��8q���M0�5�;x:����6�S��dde�t>"O-T�Zǎ7+��Ld����A�w\�xէ�We*�G'*�Q"sPh�����8� �i�t��]���g��4�G_�}怷�:&��{x��>�i*_�lm#e�LiZ��)�q�4m>Ԕ��,�³��,+�\ uVJ=��Z>��:�����G�"���N�<Y��4����4�ǖ�!�B�x��cSO�?G����A�JN�u�G�s,��w���A�x�2��vU�Շ��=�'�u���զ���\3�`A�q�S��<3�z��0����K���c!;���:�4�:�u����������_�s��������H�kE���*���ݠ%���§F&��[W�_,�m�����SA�)r��+2��uxt���$�eaK��黳w7l�Ґ;CN�"���c&~�Ľ9M����"e4��XN�5��b�5����&��3�	�w\���S�5��Up�Ɛ�0p�բ��s�S�X�lc��$��Zr��-��]�c2�=8c
�醏i���g�^�|��BoP(iP>'��iw�FtJY_"�W�fM|�_u&2,lM�7�Q�d�>�@/@�;5ZH���Ȍ�z�+�x~B`�K����:d��Ԟ��YY�"𘁈)�\4Z���91IY�d��BC��i��[�%�@�mN��R^B������=�I����V~W��g.]��	��5��-�	�(�|�Խ�ǚY�2�d�4h�AȬh�v"�ė9��,��ӝ�ɜ�F����|xW!�M�St�{
}��/��"��/+�����LEڣz�����C���S����R����K/�	'w�gdZ�񠂲`���}���<$BE|i"8���U��n%V|�����H��t���."Z���K1���kX��"���*�Xw˷Z�>��
}j�E��.^R�?�?������J�A9PӇ���#l��3v49�pI2o��*�G�/=�R|��M��f�n�B�%�
}ݗ/d!����#�� N �O��r��@J��
@����*p��ўV/��!#�C�|G��	�R)��~-�,��l��1'k�H��{�o��㔗d����Д��(B�9�f�}򩩭H���/���+���Y���v� -6��~�ը���t� �& �i?e�9���ca�]H�3��.��C�C�5P�t�GE;JI�:ɳ%c�e�%���q����i"X0h�<_~d�\����m`���)���r�c�P0��i�7��X����,%�:WNo�z29�Q�
*���������ך�[��Jj!u�2��c��Gɫ���jt��|FkF������p��Q�8������7 ��g$��[���L��=k@��
<�'R��2�jh�0�����:<��h�Pa�~�ۗ#��Mtd��T��X�-��և����(^���[��ǳs��.�R���#�䝁�j
B��F��JRa�b�Uh�z�%���������w�.�bbU���G�/Z�}f���W9�X�HW���)F^�_�MsB�:f?�$�c�dXT3���"��m�P�T�͕w:'VAS�X�#�x�'��M� 0�>Kq[����b������b�t��(w�kV�
+pHǜ�B�ԡE���m�M`���-h��hd*�ܢ���ﶽ�I��4�h�MLA�FY���u�<J����F%TA��L:#���I/9?�A+גf�x��I� ]zc^���5#=ٺ�y#:1=r�T�˛:P�wa�L4�œ)�uȋ B������Oq��Im<ܳ�y!�?���P��+*nk��Od8�Xb��ѯ�P�zx��l���&�\��K��4�y�J��m�(#j�y��|�?	���V��s�'q��l0��8����[Taз�7��>����c�J~�����ș0�|��=4N���(�����_��P�Ј���8+��q�l�t��zb����oWΨ�̱0�od2��}�Y:v܀8_�PkdQ�F'��,D���H�a|�����	Pp�:�p�Q��	�.��ܭ�QwJ�Y:l�u�{8�Hv�0�]�34�͹��W
��U��u���M����g6Hm���~������|���}�Y8�x�Ŧc��Ǎ'&� N~�o��	��Ln�㶲�&���<Fk���J�GUJ���|x7
�-qz�h��_\7 �D����K�����2p������I�	�;�����a�2VW
?�nu��J���.%�wfWZ�eXI(��@(���iDF���T�O��0~��!E�np�p!��)5�;#Ne?�N(Rb2�w���;�6�;ɽ�t�@�G��=x{l��S� K{���<Ş��@��GR���BU�w�(e�f��53���^@�05,��	}��NƠVM
�~��[�+�#�T�)_A�3uv�5~�+�*D�p��Q��݀�qY�c����a��'��t�����2T��T���E}Z��_e�;���dT2��7V�K�P��V���z��vUB��O��4�ZnmJ4�Y�����-�~�g����Vμ	���
�ٸ5�r���_E��޻�/��Ne��D���i��ɒ<ѐj�Z`���/0�����9΂�r��T'��,B(�ƒ���&b��3�,C^O�j��+q.5ku����#3�l$γBi�х �[��'��2�fUL�_��S�Ha�*��&���|�*��Q��DO���ɱ���yP*^�S6U��4�A��e�Q��į^�h�9!/��G�l��"O�Kp�E��8sf�IK2���h�:���R�b���dV�y^&	]�T�b�w��=`����ݕ��D�]e�*��A㷟�\'���L��N��d�Z�����y��(��U��#�_@T�x����O��҈���$�w�\��z�p$����z�mY8J��nY�3�q�Ţ��O��w�����v�'`��Q$��Y�3���C1N���KBTo��>�&`������l�~/*w���]Sj�:�c�a@<k-E�d��+k���	�F�JHe��_[��W~�=F��ϔ0���c����)�˴�wꭲ�A��1�<�Tu D��\���f�U��_6}6�����;�d<½:��7��o��u�qd�g/3*Ě�(���.{>��I�s�t��ZC�'�-�M�S���Ķ��]��W�\�R��H�@}�e*V����9�����������+�a؆a�y5��r1�y)~*����}C�;�= #��$����=�!��/�.��ͯ�4�s�aO�j�0�V�6�4�4��=�w{�\���k��U"�ˏ�nt�Ĵ>QT;���sb�?��b�0Q�vVj�_��Q�lx�`u�x�|�g:3���������
J�=����5�3����s�k�?�@�x������1.��)��Wy����I���K�"j��5��ʲY➠��i��h-���XjB�ǈ���O��j����e��K���X����\W�]�|ρ����\�z��z!&05$��ʹ�4lh����X�	K���B^�N��w�&ٔ��1F��'��\���m�;Ό~wΩկW�4��7�`6�i���?*���#f"�:	��݆-��(LЈ �����G��9F�z��fC�R]�塖�B=�8F���|����f�����%�"=�����?8�|l6�O9�
�X1�p�v��28�ĪXv�M@�����{�]x�-�a��Y� ����$(�zN��������:@�R`l�Cˏ@Jg��u�����kw�֎)m!��v\���Cn��^���P���Œ��p�SD�&u#'���gI�A�Kz����'�{�[���8֞E=������f�1D��˧4���k���sOnb�Cyԯ�0=*\�Z����bg�4zo���S����6j�4Te%M����~u�ЛQh}j���"��Ud$�-G��{�)�B���,U|�o�`��N҄*��L��;F�H�Z�^˃.YR�� _��Jn7
��! f�-^JK
˨�9�3���ܝ	����X�����+yt15ߙ�r��LC�L��#���/���Y���B�(x͹�^Ɵ�BQ
��KHA�:��p6Щ�W%�r�7-�dTq��#:����a�'�=c�x���0+}�4�Uws�Wm�)�mE���,��}A��~r~
 G`̑�t��_RU�{2nHG�NC��j�8F�Ǵ�|jd�e!n�L7�K���<�8EU�,��R�~���o��2�[ٌ#v.��s�_}G�\�t�N���\`�L��T:J�]�9�w˸��a����%�7�u��p��qB%��m��k���e�^�к=s7N뗪�2/��'('�V�3�Wz��}1oN�^��蛀)�R��M#���I�$�k�QL���ˁ��cB'o���c!�����oC%k�؄d��b�{ ����>���y�417�.�IR����W\"��>��
k��/��J�B����1�s5۰�QR���A����.�#f�p���n#�����0���Y2��B�an� �&����/���E��T+e������7^0�������^�޿z� �>���O�fZ�1/�VH���zM��\��%|���l�4�\���^G(�{U�� ��R�v`wƵ�B�fv�h�#ӻ���hS'�ݍ:�KN���XY�=ȯTm�����T�@���E�#͝p(^��g�a��^-O�.�g�j,P��6˿�������x=�"uJiĥ0�O�	���0$Q�^� 9���i(bA�"ؗ��&Cw��}%��6��3��y�s��Eܿ�S�%nɔ=/����I�s���mh�Ky�4��׫s[(�^��=�ub�'b�(�KCJ@�8V8�a��h���6�	u�;��9��;.���׊�{M6o�j F����GJ��Cn�*<&�S�����#�u��������+&)	{�^K�Y���[~WƼЊ��|�x�5�B��X��Mc�Z8+�R.�`���I�n����c�6�w�D!aLU�xa��z���_���t?k�ɘe�T���k|�iH�7� �RܷS����)�K�րŇy�VN.�I�6R��)8`�`�`<�ʋ��]A�?'�uԀX��	��t�g5R/�keo��|�D�U1�P_�n���I�x��pK��)��q��?��h �>8/?&��^���w#u�֢��(��	z�'L�q@�3r�/��)�͘�T�	��ԜcN�=r��{?sv�X3#
�'�b�I�� {3�r���5��"+�9D��x2\�[�|��2a����İa��@�
4�jF�&5���r.�q6��-�y�Uz���PtYS!�,3!���@{�=��^TŜ�7y8�f�� '�JH�|����(c&w�J&d���5A5�^z a�;��z�h�#��k�v_R6�+)�"{$D���7�h�
�V�Va�Ͷ��q�B�
�?:�ş�V~�@]�Q�&�4cU�2':��m|M%�uJ���XL?��e)Kӓ��D�/m4<,�o�L�Y�Z2������\ A���˽��S��v!Z+K��F߇uW䠒NA��aFB�<�G�g���x;�����2l��S�7i�Oq��3s!��Uy�Ca��脅�;�@P�o���8ǹ²���q�
�׷�J�n�oZOsٶ��pJ>s\�|:�:�9��&Ƃ	0�F�!.�:zON�ʾ|��n��Ra�G�\�~#�9{rn��:h����a<f�xO2�d]^�d�3�&>�#Z�����fX(�5UB������8ΨX߲���HDʮ&J�tz���h�9�\k��R4/D!av٨zX��-?��t��N��?����Wfދк�bB�&���a��ˍ���f�~�I�9���88��zTty����+��D_�/�D�� e�<�2)��j����`4U�ҵ����P���`!	�#&�9~7ʽ)��T���M}k͉���<O�i��h��i���(���������b��5P/vS�CL-�(��%�o�x�@��/�e�~�_ H&�h�-G/�T3�O�����;�BBP���%��>)>���b.C흲���π�~��\�"�j��<m�\��>�^&{��QH"�Û!9�Rj��(��_��g)����c�b�73�;�� �(�	XPU$e���C-�n#���dCY)P��/پÖ�����_(��j��d@V�~�5j �s/oy ����-�HI�,E"=�Y���=SJ�j�����Fw6e̋~�U*� �D����h�*�"�����Þ������E�"/)�g�9ͩ�V��JBqw<�{NͯW|�ɐM�8x�aS(��%qN�����~��uY��P�XY�@����f)�/�8<w4�ttd� �3,�5��r\M�M#���A��]�J�J~��0LW� ,v��&�g+M�)�oY(���H�mϋ���:�s����;7pu�8ϝ���Bʷ�.t��)�hEy���V�;���T�o����Fg��G f_�ǁ^��A�lz6�Ǖ�.|�Í⦫����,F��	}��s�u�/��J|)PM���j��갳�=�> ��zJ�K���{����ӯHNB��$�6ɡ}?�V�){͔�̍*�#�׾p@γ�G����B�Qf\�fԦApO�;H|o'
��Q�)�������ٞH˕k�c,�-N�*+�����k9�F��=ǅ��;#�wk�'�Eo���F~/x� Tm|��Ƴ���Ws�:�n-@���R�)���`����S�;�0u��v$Y����hp���4,������D8�$�Bvm���������*-v��kL�*�S����W��ai&?*����	�$9�-�1�vHRp��'���-�U�i%��pd���i`��� 0��H��X�ɗ6�	y��)�W��f1X�1�TJn�m�4DO��oUظ0yϗ�$�б��T���Mj?���&j���{�bV��H�le����b����s��2/��#��Ƃ�L��������-��KG�g�}�d�zyD@�X}X��������UT�Z�#f�����0��cw�e
;����b�rG�	�cU��
�N{�!t:���z��h*D��r���>�&ߥ��:3����q����TX�!zS6�Mt�s)��U��q׍L��m:��B~�l�[`���*͘��ۊ%j�M#���\;�p�������K�p���}1����B�=�#�j}�8`�oOZжNF��B��H2��>�U�F ,�w��� ����*�P�G���v�"���KfpP��Od�R%�� ��B/�)t{���W��y����v���0)؄�7˗0��1XC$N�杗�W4�I��buzA���ɠ˱�7���r���0��ta=A_u��0��7����#��,�x`�x,~�֚��1�w�9��Ye��M�l(�4$��[��l�a����8��ϰs�$��=�V|G�]��6������"�HIF6�V��,;�$i��&`�ā��H�w��.%���F-^�,��|�?k�i���'�a��y$�D��
Uj�Zc��Pg��`���/��X�,N��]�*�qY]�^θ��ϼ���$$���\��8&W�˶��e] �Y�Ԩ����we�}m}��y�Z����!K5�Z�����-��,|����j<Z||ɋ�rh9�� ��=�s���M61\h)�ҫ�ch���d��[�����s��2{%LI�4 ��ٹ��Ja�vJ(s/n�Ԝ���{2�<�
A�@��/01!����@���N(%mb뜳vcrkw���h9��A2f�2c��/�\ˋjD���X�`����ݢ��u:��L �ｧE�		lxO-W�c��G���s<��޷�pdV��p�ma����fK�y���	`�L� x� �Vɯ�$sq
C0���=�ٹ�_6�UVg�ν���1O�����Jɣ+avr
�h�aF"�>2�fl�!1Vp]B�fn�%g��1�]�^�U�jP��	��J�����U�Z����öĿT���E]�����	����(WܻPDz\@���������>n���������g��#=?��1ߚ��$b�pͰ�� ^�E�X���Z�9QR�]EO��È�{��jh��A���5�ʯ�.���v7|!���$���8�&7NM9+=��#�2@bp[nB3�e���Y�5~	�A�S�PI��3Dԉ�N�	�{�m���Q�~�����i�*@�*i�uu�q��*XJƛ`��jy���7����N�X�Czfi�V,}S��SxK(4G�A����v��D�?#�!"ix��*B1����d�����T�C6>.ߗ-��7���2����G� � �+X�0�~��P��q�J��V)Q��w��["��#yC&)��d���&�K�|�<�UBp�rO��[��.t�9�
I��!��h3z���ʑ��>��+ ��W���_��3}���h/���@�L�i�(DW��jجM��Н���T�L�[��[FY
)X[؎l�M����z����z��R����3����R��9�;8�n�����4���,T�I�O��̻m
�g$3�@R��<��:��������1q�DE���ο@��疈�)�:C�������Z�9De��TͫlpI�~W�7�-RW���w3S��t�gu�$pkA
��f��]�p��L�e��"�?�_t_ʀ*�24l`�3�^��e�w��L""�d�Q�,�:��{�K���ez� ˽�%Si�Kld���D6���#��b���'$���b	#�R������	�ڬ��sMr1�v=��g�F���Qz��eBc�T��_~�	�0��)��>�.6怪����h��˘��F�>��.�dϬn%�;5.e��!�ZyǠ8�![m	
�T����Bs��� $�L��L�<T�9^���(>�x��2V���>zF�b��~x��u��OtyO�[��9E�/�M�������h��#��a=Vw���#e�/y#T$�;>�M�l��x�e���!���P���bKJ)o-bC�]��7��Y�⬰�G��}���q�ҙ���6'��7��M��	Ee���e���m* F�&��$[=�/�+}��|� :�f v~�Ru�Ws�54�����ڄ�N��2��¢����V�1�21�S�ڧ��4ĺ�
&q$����t�Ç,�j�D�/2�g6W�+�,���Al�Pg�x��$~�j-3ȯV�	�4����:�����:R�L?����.�faKoMI0 �Ⱥ��&�V���䯶�ۂmaP���y_J��R�7�[%�)D���-����1&��Ɣk���k��*|�$�����t����ĘίG,t����-`-��CHk���*
�۝E���� 
e�aT?�D^�4������N��D���d�����5��������/'�oC(�,V������O�b�e�<�/��D�W����-a�m�Ҽ��0��!�Я��r��+�B��P���E1r�W��[�d��[�5�`�t�:�����q�yEG�w���~��mS���뮫�O�:��p����8(E���h�4��&��4.#*�&�(k9�œ]����X��Ȑ�oe!*��!�Y$�ĥ�;d2J�= �����]HSEV���?ݡJ$��z�'U�)�3V��-�dh���t�`k��rRUʀy�����>�Gt�g��\%ij�� ����tҒpF�I��Ox0�`�~''}o3��y�LW�9��㊾����"���a-��ܬ{������T�u4��6ϖAV��w����I�!�C�W���Ň8?���2������b=�w�|�3�A������,d����vq�n?�}e,�2�|ʭ�k�2�ډ��Om����ӧ���Aa�0T1������5oZ���"�����.��qd`������O��HT�����4*渟�$���k��p1n��:�����.�"��}79���3O�D�J�����	�*$�8��}nٖ�:{W@:Y_Cx��[-�U�'��v5��P��O���K�ƝY&�i��[�|������.Hn��@o8�Sֆ�֝'5q��'k���l�].='�p�p��.���	����/[S�͡������<�ww�8;����;�d��TdO+.^��G\�����R
�n��9���^��7�0�����')�1J�)\��/`x��� J���pΆ�Юy�+���SeÂ�_d��P�uxؤ���;�9܍������;&R�)��nh�y媭,��/�F��������ɟ����:��e�kŘ���X�q��.�멕�:��OS�c�b��(�g;Z.vrS�W�/ō���m������J�L����2c����&�J!K������3ţk	��x��1��P~t�"k|�k�z�G�O�c��Ȅ:Mmh'_k�M���ʯ��#�;-  ���7�+5���W-8֋��L'詟s��^���j+��wH���l���y+�!�l˽�����ko�2��fu��u�L.J�8`4�]�2)Ѕ�~��C�=�;��5���(����ʴ��N�ur���k�I�e�'}��v�#���דU�!��RM���;J֮��r$fbb���Y�W�D؏���IY%*�mfeN�����JBx-���,G�2���*|$j��x�4"�_=-[8�yڕZU���0����B��V���9D�U�(��ʺb�% bU�Q�C?A�pU�k��*�o��t�)�f��I���_�:PS(��ԡm0��m���� E_]"M��?�%�U�f8��ӾZ|Ӽ�NCF��阑������X�%J��p�)T�V�Ao��(�J�!�^P	�c�U� `ېN���~���U�nw\INt�r��sK9I�|f��xp����61d�O�9'-���m�~QO����?����0K�QN�]<�˅�6�����Ue��������E�5��_Z�/�l���f���)�P��u��
M��h��JC�r��~v$�*¯%ѲQɆ������HLx�@	�����,�+'n��TJ̡rB�ytr2��h��SPc�W�J z���~��H � o
�.EwN.���\!=8^�^�G�i:7����j���
BM���]Tk:��	Y��q��A��N��m�ݯ�w�v\�7�{������k��%�#����ml��M�0n�R���I��W� ۗ�u N�hy�%uUZ
IW��="��@S�VwM��(�#�ˏ���P��0Z�/�չ=�F�� ����=�V�"����B{��-�I��\5aN�XiD�\p�?''{�+cQ&j���S�r)�q�c���e>��g��� ��#�?@�QE
F;?�����6ɛVNuk��,|����:�<�$U4H�]pH�_�b�C�cJw�W�8�+�I�d��A�0C���N-�#η�@w�\깏��Y��Tj��_�9Jn+b o�� F\���?B��tx�K�����7~����d��#�Ҳ~�"2�'���|��EQ�A���$Se {.���ڛ�Y: s�R���h C�F/����E}{֢��}x,)�V�����a�r�.�/��(0�w�7⤺���7�׽��hDŘ�v7ѻ:����ϊYÑ�fY���$rg�%���X�j����R,���;R��#ЊR��h������=�� �y���5�
�7^�����ZB"^��0 Oe�ѿ�#&�����s\6pq�n6���T��A2Ln������c�*����h�����6��`��Q�U��ͤ ���F��-(�G^A����D(e�!��D/�y<�Y�X��*_�;�8�d����ؤ�s�PIf��ift]��!���9��R�c0��, 5��9-��hvO;Ho� �@�����IZ�Q�x�=W"	ӵ���2P��D*W���m-}x%��:�Y�[�� @$��ǔ����;��X]˧�����i���� Aa_���6ˀ�XV�+��.��*\��~�u��9�d��34�kP�+�P��E��A�sk9E0h��L$6M�TrY�L�0z�PK;03�{���x�D�����:���b7I�T_����l��aʊ���z3���g+�wT_ޑT�h ����-[��!ik����?9�[j��ڰ�j��?���Y&f�@��(7��h��B
p�v���3$=���o��>=��ũ���'�G���z �<����\p�DV�-d��ŕ��P�����JRS���D�E���GW�twW�i�%#{��6��4[Yud�������}�7�t;v�:XCma��h@��x�S�m+�F���X��WO�e@�: (�*l�2���jf/��iް�K/����d�RMۋ�*��	��i�@N��i�@c(���mne���%�񞴩�N�x�Ѩ�R����7���p���L�ҫ��좲��8&�l��Ž�m} �F��;����.fƲ+�x,��TF�3��� �!b]u���S=���R�����Y�D�[��z�u�m�E_�/Q����#�Ǡӣ~7]���-�V�Z��\5^˕+�5�����_A�s�8������S�I��XkNn@�H|J���z�X��o�x'Qx_܋6�(��JH2{v�~�1�+��8E���JӅ�iC�~,޾"�N�T�Q�>=��#�5�r^��Ii����F8��P�hq7d��� ��7;+�>Ƴ��]]T�_y]V�'�u���+u���)��D�e�O+�Zr��y�	�0+��ǥ�1q�h��R�gv�ؽ��׫^�zV�\ݢ9g�c�Oj�ĥ��q���^Z>�D����N?W�X��E�~�1ZiO��7�A�Ё�[��2���S�˱���]X�7J���1�?���ӑ�q�P��[��&�Z*�}y�ZBd��i�5㇣sZ�H��k@j)��M&�W��1�!�87[��A��C1f�K�����L*��+�,�U\����j�K'�R��Vh���e߭�i&�(���q���+u��n�4-_"�a�l\�W����5�ض�p�ѿCG�w?2lP����;y�1Ke��o8��?:2�+j΋�z�	��}g�g�)�b�l�d�?�y�L�������=Nj�qF��(�a�Ks�E�:�L�����_��
�
3{Q��p����&��a6|����_�	���nK�Η�� "�{"�& x����u4U�+�7|8�e���vM�9�(�O:an�����o�D3�C�u贝�p$;/��Ic �d�����nOړla��a��R�r��"��$S�����rN�!�����a���O�/fr�D]i�0�_>f&�~
~���V�ٚr�������$0jk=�.�v�T�g{���m%�d��	ηэ1��|����̸����v��������~ӿ[��s/�]뺧&�߹p�\�@�ՠg�ugLXᅶ��S�u۰c4gr���u�߇����_��`i�*;pu��ɱ�мq���8����y�hj2��>t�||�f�f�)=n?fz�W��'��=@,%�H���J�j2��N��z�kK6E�d�#Ef���4�YM�J�a��-6#���f� I�t�#�ZR��C�N5���m[�m��a� ��ou�~�����<�/\����2#�2�8�?�ߪ����S�����dn�1;
�>���7�"�PN����@1�NX�D�0���iPf�*�"&=,	�X�Ϯ�� N9F���EC2]ޫf1\��A͉��:��wy]��/�CrEuQ=S�l�&�(����n��PX�5 �����!UDW�h�*�ϥy&���0Cb�+�%Y�Gm�M#��0kro�`��-q�S���z�<;���r�.��m����ET!�춘8��C\���ګ0]z���N���	�-]�����%(۽>�8X+��Y}S����OU!$3)?�78/��'M��9^���en�j�Du��[�oN����K��e�ŭ
���I�P��L�h��jª����	���^���	KT���B�2�Z���S�Ь���sS�� ��&/(�S�i`�4G�S�[H���ҥ^���x~G�?�Ā���o�KAs��P�<��)��|-棦��ly��?��C��@�i�!U&�EQr��w�Ҍ`]�z�l�2�F��R��yH��ʳ�5&�I�)̣���"`} �nG�:�nЁ�xK�[� ��lE?H����R�t<T��4��J6Z簢���?��#�?�M	? Q[�F��y�R?����y��'��2 �cs�-!֥鴯�����@v4�̖��c��\;4��J�V5|"�Q�c�a��c���/j�����H4m��$;�����pBC�%���.3�!ZD�����C�%(0ɗv��%a��}𯆵~O�c�����~1P�ׯ�