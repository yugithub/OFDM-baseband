��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��R��g�p3����Apǜ��p�~��!�XZ�1 ��z��Ey5KT�Y�T�cy�ϸn�:�|�4P�G0j�����0�H��
a˄z9��Ә��ZW8�|�C�F�`�'�/	��;��)E�)h�h��L�ߦK��j-��9*��	0��d	�����*=���ic�����<�R��=�ec ��X��=�=���m�F&����/\�'23�!A>�d�`�Нpce���և���_'o�n�ߛ�N�3?���ƭ��S�y`�V�>��(�_�<��3 5�r��������qHf��D��7�"�T��+�f��Z�ih�(6�HN���j��z�h���.���i�Ȱ�'�� �V$������T~V�f��VR�O0=X�z�H:�b��d�6( lfmP�O�t����Cy�㪎aJ3�ƛ�}��f��6�0����{ǒdK�* �dS,(5���sV��K�1��y7�qR4f�9ps.C]��p�W�uY��~�V�����*�Q�����H!e�`�b?eN�5V`��Y����V������4uZ���z�!����]����������ur�I5��u_"G����w��)ߡA�Tu�(��&�K�d�sAQƜ9��>�"��=v�SK�2�ZId��Uy~���2L�/*���	ƈ��o��QO�[�Y�`w�j/ձ?	��kr���3]AR�j��g�X��t�Z�Z��RB�y���wY���>B�n�b�?�K�X��Tî�YB���H�r �S��؇�U����⊰g-��,2�jnTi;�+6ǚ]>X�qX$��-PN� ����ab����L���q����X��.�>*��p��e���=Y� ͻ�s�_��^w�K�����1l�zإ.D��!��nx9^�b�����/>}����;����D�i�����ArY<&c,��v*�Q��	�0���2��3Z�4
*���{̭���R�F�Y|\+����\�S�+�:������û�y��J�ďq� <�iV͉;��v�8�FK�d��#�
�(���1���[�}�
D��[<�V
��o�}^�9X��r���Ry�g��(l���l�F	CV���!Pl���I;3�%ݔ����I�\j������s�+���(��\ Y�B��v�סR�z:��Y�wfq��~TD}���wM�-=��J�m)�����n]��7�g;9���>z��C��s1�]� ��%�ܹ.���M�߅�����85��m�^^�t�?.����u���ӿ[�>oˎ������{��FI����/=@�B$ڲ�5��]�T��I�>O����P�Z�K8?+�x)tDu�Ʉ)�W�f��P�.��&��/Ad��[��f���PWr�:�����`S���*�P����91�}�n/�v�Ɠz�9	��oK �>dj�C�����?T�]E|ΗO�п��>��Q��m�L:S���ě���X�dl�1YrB�_����ݜ�Б��M�>�esuM�b�(�T���D�����������m^�k���}r����~��9��Ԃ��.��$�j���Wǖ'�S��W�}�e�`��v�@~�Ν�i��7�]>j��Aa �6�����3���3�7�@Y(���J�k���X�N��#��q<@���\�l3zT�o�= �g�v%z�$֐g�jkqś�7ޟ�����o;~K�r�,3f]��G�풟��_
]��T�@V)��`�ݕ��U��؋�����Rp"&��.�>���)=�!��|2#[�#������������_��t�d�D1��-l�Ou?&�^�_Y��>mzA��9�n��vm�&����vJ�,05b�����m��Ƣ���o��[}9֒\|�F���l�� �I��:x"�9���ZZ?������o�L��H�l��Ů����Q��@S���AQa$6��D(!	���#�L=��Z���%j��D��� �`��\�~a; ��9�K;�M����:���Y��y�Ɔ���eQ����v�E�g�,����M��m�x�s��L������|�~��!�Xc�*_�%E���U�
0ʿT���%U�cf��uP����`�6��Y߇�m��l�Ƴ`���:�4%iB�LU�$�X�E��(���NPU���cub2m�*e��j�6=�7�<lR	��	��Wŧ0��U��0��N}�:�,o�y�n���9"�o���G�RVȲ�9�r�j�&�6x��g�6ض��ƫu�89`ʆ�����cj����4��?�P{gbF�O��HE��zx�!%��q�!�_��6�]���K�osöG�c�/��9X�<&� �U�~&g��㗀Q�φ�s��'㪭�v-��_�+ۡL�@Wz�2x�P}����PR�D���z�����\	��чjiCr��^�<�8%�,��mnV���/�?��\�X�Ci<�oIENf��h�����K���w��7��3�ђ��q�b���l;)�m��(���:���,|�s�yي��H/E�F蓪�ї"�ڸ�?Ro5���FSW��J���lԲ�p߱˚�!��h�'zko�#`�3&i�54>����{F�k�V��@��*Lw�!!����G�܌����Ѻ#0��9_���p�]ibu�;��(%9ęJP���4N$����
)���4��9�����M�:� �ב�ȴ*��9BaocC�-R07�k��@�7��$yމ��y��=���s5+ۉS L��4� r?�%vm�����q��X'�%�E���+l���!��Y�csj� ހ� ��V�/��/�z�ʭr�8d��
���^��#S� 3R?AS�.?/������̵G�n����7��.��;8l��G�ܨ@*_T��ͬ��6V1��>wsu1H�2��#@�y.�=�20DH���h|ɾ�e_].��*O���Y�6���6YL���ߛ$��aVB���tC��9>�Ō	������<:��fxgȖ-kB�9�f���>�����L���H�q��'$9��F��vR�x�����W(UV�w���Ki$����0Ӄ��=�A*��Y�ui[�31[�b��ė��&��,�T����k���uo�b����}杏I��s�/!j�'L�J�H�S�����Q�MΫ౸�����ڿP|��O�m� o�.m�J=�+/4c
�}g�v�.?����=I�G~�t-O[��w�ɞ�\��?'��;v$�"ǋ�Q�VR�?E������