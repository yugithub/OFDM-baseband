��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x������jTe�)�D�b���A����1v16�|,J6l��)~�S� �B�`q���(]�s�ˠ%��L@��z^ߴ�E����\>lt܀��|��>Y-��=��v�r@@����Q��2��^ԭ>=h��^$��f]vY� $za��"O� X��R��ȿ�u��v��\@��
��^(9������U�M4�~�&om^���O�|�;��9J0����E�{pY��W��AHgI��o(�s�����SL<�9K�	���-R��_�l�gI��9M>�5��׎m�C����E��V�e�C�FU���n%{��
]�^
;{*�>Ԣ.Q����ǿ���_�#�q�ƞEE'+E��`�H��/d?���� 1)�|鏺����$�������,m�����~e�~�ň���jeU �62�D���=������v�QԾA �:lj=�Md��1��q��Z
�I�JP'6���<]�+���wMp�����M�^/ݣ࡭�4�SY{��D��yU;���Ԥ�a���`h��G���RG��1M��0���}�'����;F

�'D�����VᷜG͙�ں9QQcc�D��><|7�~�@x�}x4����,���Ls�{�U���g�?\!*>�z=�}p���+6�qf���R�72�$�F��`��پ����Y�q�-�
�9�pai��[��<��~�Q$ՙ~mI8dº��[߇ ��9��6�s�	�
�&���F�T��b�Y�El���)�=Ln�]�����Xg+�̬�� ��p�����ߌ��ٓ�R�'��q�5�����ń������j��dVyR~7�"M��O1��g���y|QD��U�~�,�-"���=9��+RK�x�c�롂I�>�l,,0nK�P�5ո�H�1�����"���2a��5l1!^h{�b(���R�f��$%6��Sj������$����>�C(v��fH�m{M�(����I�����O��N�������2ߌ���������` �d
|l� ��#O��#q�4��x�qP]�[L�i�.�E2L���|r�N%�Is��b�����&D�m�O�ޛ'�RM�S��m !��>�h[���u�v�CMwņ1�;DQd6��<Q�"n0�;��TrA������<N���e���d���0#��1���j+iwh
6v�ᜒ�^��9�&]\�<�X(#D{��Z�%z�4
��~#�G#}%�BN��k����A�X��Y�zd.���C��� �_�m�D~]L�1�:G1��v.�k�
^�)[��-�ѝ�Z�Wfϒ���Axѡ6�IC�*PD�U�����a95eք�s�h^��&ʷ�  ��VMN�j��9��X�{0�#/�kݙ����@�����4K�U���j>����t�K?��W�0��t����]&H,!��Y���1�u �|� 4pz���0��Ng=�c^��rGy�4�\�뉣�^�5J�X%�pr��~V,���԰.-\?�2�s@��En��k�t�rU�����ά�ۋ��8���,��t)��R�S�]T7����H���v�ͧ�K�Ĉ��mң��-l�V���N�g�u�S}IP~��F�J��DJ��I�z�E�@�-$����)�Dn����A�f#�TUu�N��s�k9{�(O�ύs,�J WU�A����@�<�&�?f☌A�!Ty�*��X(�}<�۵�K��t8zb)���X�� ;Js���q��B��ǎ�z%�U��4�l�A������U�c~�DLs���}�)�� H(~���k4�͛�����뚶*+�gTH&����`Y��v���Q��h��6�Y��ѱ�kqR��Q��h:Vo#�H�:<MaR��^�.LG�k��?6Oߕ���w�k�Nz��iY�E2�V�R�dm�`��^FL�G��w�����4ή����3�Q���RO�x'fee-7���#9����װ	g>4Ŀu�O'�3�;Qy�"$<#	A�+˞p%}!������OZ��!G�릳׻!q[�R�H�T��ͦƒoq3|���#u\�5� ߴyr�o�,B:���y�3�^��$��]����%�;]��<�~?��H=��ğ�cr:����o�	�>�; 5�T4d�j�]{'�tB�1��ez��9��l�`*�g�[����}c �M��.|�)�=pI��(>����ו�Z�A\G�=<��v+*��͍M�$.S]EE�eg�y0�t��YU�!�xqn�	�IK8\�����F[|��{�x�'�$�~���?���7�Mzm�J�N7��̟,]qQ��Ћq���r��{R��������/�[���wT�Zmʅi�v��t�1�aF	����bd�C�2n��ѱ�4Ќf2m�`IHH��XA�Q��Z�����C������͒T�#C�6�Fݮ�IٍAG��C.O�x����9��zI�����������z�٢�K����R���K��o���uU��Лp+���n��8^��3�K��4 �&�K�,R�aM,5���kCBaE�7P��]���/�(/�?��p��!4�I%��@�3�Z37��Q*���d8a;�#6
�D1I���\A��R�#5hԶl?T}L�ɳx�(��b�tȰDm?�8�j��:���5��mX���$k�ά��Ҵ�w)���X��Ym���P:E��7�V�l��\Ҍ��^�aҕ(�A�ԟ��i^�۲z����9X?xX���
��,����0Q���#N�C��?�}\$�&䖼����A�y��B�C�|R�g=��$�0B�I8w�%.��R=8V >�x��B`�^k �j_YUVbL.Ϧ3;�����A�ꦯ)�%�i?ӢJ
!{�n`>��ų��S�z�Zظ��(�ʤSո����q�U?�r�Q���W,�|9��x�^��,#�?W��� 33 �vg�І�pȡ��[{i_�C�_��ݻZ���T�����("���԰������2�΄�OL#�i�]�Y�'B��7�3�PiVfi,�}8in��j
�A� �'��և�yҳ��l�唨ڸޗk*�Ԇhy+�����t���v�� �����I൮�nMF�'��޶N�6�$>�uϭ�Cn'�	�@�u\�G8��2#�����o#q�e���3�M�|�ۣ�8���T�����<f>@�}xe�|A�(�ݓo��R���B�$ʹ��Ćd�_:���a�x��5��Zn���c�[����>Pad������a�F�h-6��ۋ$�!�Ǟ�M�t@_�΢S��_ĝ�Uw�
(U�� �YD�z��jP�V��K���l��dбy��.w��$��x����+0�׈��,\ٚ~_�Q{+B�Ӡ| �oX�q��_
��1�.ۗ��\��q#�?x~������v#��[F�2l�����8S�n�o�o|���|pe�U^F��(,0F�ۢ~�b�J�V���R�Pǋ��T�����冂yu&X�m;T8��i��E[������H�IBJ�=��I��Y ���{� �ʤ�~K�8���,^0�Xct�%c�Q�Ys��6I�����m\,��S�*qx���}��#$~��yl���,�#����$^��d�K�=Ȩ��0�O��d+w���Q�vuVg`:'|����b�w�S6k�^���P���K�D�6G'c���ORyn(ф$h��F���?;	٣~o�g1��[�;V7�M�m/&�l�ٯ��k����v_D��'��<γ#�3� �����y2����jz���QP����*��Fx�.!&ʹR/�˯���.߮�H��l �������RC�@���>)��7_��]��?�L=��>������X�_�d��|���.�;��IZi�z8I�q��/�6B]��K���;�����[>��bH7꣩1u�i0�>��e3-���рadȉ��m������.��"5rJ��K&��t�U`���9���a�w�y�o-�E^��"|�zI������z-o��>�l̓{�s*���h1��C��%��c���e8 =�h�z2�kV�j��q�XP�5t�7s�v���ߚ\`�A��d6���g�!c���;h�:��K
2�A�Jz<�ِ]]�`]�sU��8��d��-�0��֛�b���P��e�87<��Lt��������>��V�	3B�g�q�r
V]��Q��<b� ����3>���b�#��6�P��rA��
�',�z�a!��ڏ��&��w�&Xy~�ɲ|���4�\`"*�th�m	�� wy�(B�y�b-N-�-d��`g�w�������as6��&�j��?}���<b�SJF���\w+8xb����=j��{i�."�bŢ=�Ky���'���6r,!�,�Y�3�w�,T���\���y:�a8Xɫ�&�FQ_ƙA�Κ��}�#~�&��{!���;M2V$�����$[���dRTM��)"x�a��S�vFڋc�����r�.��N������
/����1���.��Jx#^��Day��WQ���r��\|� :u\a��8��ѐ�Ž?����E/�>,)g�"/أХ_$��U,c9�m�"�B���r�1�3q���j��Q�Ȉ���ZH�Ebi@�ðJ%�6����1=oUט�S3iK�/8`Z�A�[�Pb	�����������Ks�B&���ƙ*蕞E+������@�6PZ~�Ƞ6ˣ	�:&�^$,��ER>��`�!�R�<���0���rR�"���k�䔨����ӷ�J�s��?W����뾐�e�~B��[y�C2���lѾ�C3�x����P�$t��_��H�P�n�L�po���
�$N:�ib�!�c}�p��@��6� �R�r��v�����/���NY<ȶǾno)So���E�l��`�UZݵ��n�8�G����v�����:n��:�N$�V�� �����|��摁�\�^��ν��j��U�sTDI��чp���|����]/"��$���0����$�ٌ�5����?�o�)���7F������+���D~=b���+`E��3]��Tp©�$H���H͹�ڍʶ���������0`��pf�zu
KZو���m���������S0C��[�	+*�K��L{'ԥ"(.O�Vc@���<Q���9����$F�9<q7��G�e�=d��Lʤ;a؝L�Dbh�ˑTЀ�H�aC#��s�E'�����8`�G���. |2��o��������ڷi��&�h�N[�xu��x�y��v���;##�spq�"��w����߈�MⓍ�
�����Pb��v��D�� N%>r�m�"�iڸ�
�烘\�qzs9���a�J�_�oF�l/�h1R����t+;����ذϬ#��`�Y� |�e�Mw������w����*���!�`V9H���nў��x`�3z����������Q�Ko�tX�4RI�Q��=��K;��c<|A0�Ƙ\�Dx��W J�}&��oVA�*-�~�[��\��1����1���vHƞ��/5M����%|a��J�`N����[����Of���(#֘��5J'�r�fu���T)O���̈�n��Q9�B�xV(;82@�k�4�K�5j���v)�ty�O8da�]�T3�{������R�+/Si0��%��{�T�V|x��K�/-���1��1�u��~�,NChv0E,��׋�~��R�cZH\����[f����$z����5���dΠ��}�S����な35�H%��M(:sV�|;�W�DϾ��Cn �GY���Ƕ��x�X9|�%��'R�g�J����<��_���\�C�4���A�_Y����Gn�}���v���)!{7�^d{!�juE\�)�b����W~�2��:�w���:/f�q�רIw�#��b˲B��/>�4�6+=�3]�3ҽI�W� �&-�.ö����_���ߗȧn��^�PK��%���ã-Ko����Z��/�Ro9�ۈ��W=���ݤ��R�_K����_�=ׁ�5�:g����T�2�g��&x��g��'�9)��}'��'�5����^��bN��@���f�r��r�#��2G��`yH�S����s2@����=�|]���d��$�`��/��;ny��>����5��Y�:L�"͐Aczv&ΰxf�M�;�:���B�}�d��P��N���=��p[m�s����|M���p{��ez0�zVC�񚊪��+Ӟ0��Ү�g�w�^Ѭ� �R���^��Ev܈4\��!�a�=e��d��|,#��)Oĭ��m�6�2'E�G�-.Q��
V��r);�,�E�.�@ ,����x��)�T��5�e��VG��O����L��(�#�B)A��~PȤ��Q�-��p��{�;�"- �g��y�5J�4�C�~��Q#b.���&�W��X��#%���q&��_��_�mF��"i��DCP��U<2M�ujɳ#��dзJ��жdW�`o*���ቄ���0r��J�c%E�����P��	(|��`���PW^ajB�k�C��p���lC��Y-HYCJ�P��s�o�X���v|��P9|�gQ��YT|����`^�V�8Peb�ACV[3��yRk�JP�Vs�"BF�j��	�y1��o��<(��̽!<P׮��b�?u(��(k��m>��j���G#葡О}�2��X�D ����F
P65Ny	(u��o&���먀%���z`���
�*|jqu�p��>��vҰ�Jg<x�u��*�R�-jD�!�S�	݋2���WM���6��lL�ucⷎj�0�
�n��~z:%�s��R1�Ǔ��i��BB@��P��a��w�����)��N~�3�[1��Q9{���BA�T�b3n���wq�p�<W ���KIߨ�PL�`ir���+Y� "y�B_QՕaN�� 1�k��<��ҩ����W��3V��*�mY*��Q[��6��7%�	ג���n��ݒFe[��ϫ���-:�<ż��zpЈ�%}s��(O�g�m*u����a�NW<��Q��l��$�j=f1�Ub�_��T�b���H��;��6�Zc�n|b��5�¬gt�aV-s�<�&�/��Y ��n[�l4t*k�(�2M�:�|����@2WO�*�QT#�Ǹ���]����qJ'�G)W�|�_�=`��{c(��_j0�󝜶9��^��h�L�>��&�13�d�h�3�b%�o�6���l�U>ѫ6ޮ�se��6�r`��<L�V�2nQge"�s��"���6�=_Df�TLY5S�/��� vX����um�pn�_��e�4ڭ�Ku�*�)�A���~�ֈ��^1|Q����l��x����Qa�W+�Ec�$��y#��@��[<9�6!���g`C>L�A����Z@�����[���OY;i��;c�� C+�O�>^�K�!�ܗ��9nO!9Pv�.i�w��)�������f�ʁu�`1i�k���1��DW��^��?�gC`���t��6ʱ�  �ۣ��Ńx�|�ow+��Q�#��<��k�p-��$��߄Ʌ
;݅�}�C�ó0��$�P�n:�2�W'�/��'�e-����������_I�>�X4uKG�s�F���$�p�cY� ����p=�d� �)'_@
�㬻A[��J��[�D?�?W�71d����%2>�S�1��@����7�#<��ƍ�B�_f�+��#�arX(�!F2�	������3�}�#�pF����3�o�ɡ�j�a��B�F�kn��х6v,�V��u�m����Qڹu��#Ǳ��kni+ՠ6��_�F���-����bx��4u`dɻ�N�;\2�lI��gb��d�?�
�n�g+�ĖV�Z؆a���8s�R��H^�g��"D��k��XeHѵ�/�Nh$'S���<'�MS\�����u�ӑ=�̽ȇ��	�#@SY<�JI�p�?���8��.�,$����=�m�@�Рz��@�A�-��'�+Or�â�üι8`���E�:��V��$G��Qd[n��8!2���M��Gz�[ű.%�p��0p�V�\�pەpy���Qd.�^*Ȃ���-�Ꙋ�Y¾ɤ!0\u!��*T��Fֿ�דUBt�k����7���f�
B�X��bU��+���#>�l��ˠq��FR���:����'�~�c�"cV�'ur����L$�a���I�h�0��2�a�69���.8bV�8čg�`Q�#�$�ʱf��2qC�Qʔ�d��e��;�,<�ǌ�C�ҋ�O.Ê>q�����_��a,y#[˱�K���b�ڎG2�ۼ�d�%Zm�_��ㄆ�6~�Ǭ�����]��'�u,bN'.i�J0�Zʏ�����+wKJ�/�;ڰ_�W����۔�B������q}8,F�k S!b��[u�.���@
�����1E	��)�4b0�������EtD(7�*c'􌌂��D��x��K��H��Ұ�"�����cF��[`ra.�}�\~��,/d��!�{�� ;���W������hn�|�O�~Ks