��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ���!�T0��'���Q�0ŇJ'���2"�z`���^l"l�Ρh����Gs�e�����DJc��к��w��ʰ!Bgz�x�maaw;ۘ�p �U(�� ������(��Pϖ�����d�"V����bk���M�))|=��[�K�Ö�uY�LV�`�}�^�$҇*�`�{���1�J��ir����&6�a��Ks�H�}~Nr}��w͊���+���HA�X��m����y��wUY���`�-���}8,���%ӱ<'F{mg���  H{���)���l�
Z���և���^��=	��)+��
�X��kJ��}��V�|�@I��^�`0�:��٭ϯCz�{1�Z��V �G���öP�[�ԝ��|�S�'b�C�ĳU���\���y!$��oaA�OW�TΑc#��@h{��4Xs��lCfB=�&��m�fp���=8v����j[�.��?�AH��;m���u�����\����x��\��	�G��k�t�\�:��sp�4������K�H��s6��$�Q��f���r�ac�}���`��ɮw�;�kUl�z��u�=,3�b���*��L�I��QPci$9T�C vv���[��W�и��O2�NN�`w������#:*\����+�td��Ji���b��03��G�L|�<�w#���35�8�xl�KA2R�8��?�QT�(�՛ B�Ry�v�o.�O�o��7��k�\����#5~:�X�
��,<���M�F� ]��p�3Ш	�� ��

8�b����^�3�ߘ*�@�x�I�˴�{�e�\�>�H�??"n�C&��|#�-G����z�i�w\�F�v8��/�����l�Ϥ����f���k�"L�O��r	A���5��ڟ(�!cn�8��D�H��{#��^T>������d��5	ԁ��q��AF+��#81�`F<6��/4Y���|JF'��o��j����N��L�:Z�����%;���\EScix�e�5Ӂ�~�Q(�7�,��n�+#���W�|��#�B�M1�)��J�t B|{�2Yq��=�r��!���I�`���!�i ��X:U����x�b!����]�Z?�VP�>Q�Z���K�/Y�zJ"47s�]�}j�/���m4�Ton������_:���F�z���j"Ρwn�!O#��7��$Mד4�lج8%��ɘ�a���3�q������Z`nq]y6_n.7s���$QMw헢�&�rE�}ԆU�����,������8�7J�Q3�Q1��i(�ޖmV��\�06�c0q��_`�8lV�/�ұ��=Xu�Ꞻc��]���6�^h��2$�[�ҙ4(����c�SAQ��m���/w��aQ�%��"�g؋R���;K�0�K<CY��$z�������:��	3�0�-<�9��Rx����!VM��ay�7)�~�m��,��tP�:�b�g:=�6�<K}8�V�2��P�3JƖ���W�ȍ�N�uOR6ō��jԟ �J�5m��MX"o^Y����&���8��� ��JN~v�lJ�MA��b���Qa�\��M�R��
rx�u��(��L��h$�^��j��}A���ʨۖR}7ZL3�Y���V�p��ә �n;Q%�7���,`�.�q8%?��R��}T��4��T؇��>��h� 1*O��]7�ѣ�猱
���c����9�+@:��+aY��xp��~�W;̝��,�j;��mZ�WE����(�-6l�(aˁhw�ʹ��I&��9M��^.n-�D~�$�����ϗ��#�jzp�خO�P���+���Y�%�W	y�^VD���շKEE��?]�������q=�j����~���&�H������#��i��&5�,�ٖ�N����`&�Z �����Ne�Vj��O�&tZ�����
@W>M��^���G�0�e�o�Zbo$�����k8W���h+�]�GWz�������r_���g�����o1ߞ�Ӊ�LQ�m�:U�}+�a���v zٶ=��$�麣!����X7�\7����T������-%^Y����ə0K�z��u@�f���G���~df�La]��]kF��Z�1�=Й�$������i(�>>��%�Ɵ=+�(	��!3�e��_�M��Ֆ����>��jƜ��5J*�k���F��~�h��MS�3��S	橡�a�N,��^Ձ�pV��ng��� q�~W��z��X�(�}���
ݹ�J�@�Ly��=����|xe�	�$�JB��f�l��E���3Ҕ��7�Y���¾�G\�w���֐�µ2uǾ��
�ʞ�Z�<��Dq�����=СNC=��6q$ ��k���;�
�.���ß=üJP\���c>�^�4x ����]T<�*�Q�V��|b�/I�E�t��S�Y��R��:'���n�,��c/�o�A4��Vf*��in�}��:`�W�����n�y͜�ӵ�Rj����S?a	!�E<��RD�'i�*DV"�Bi9"+%n��jmAy���cM	�T�n+w��<p��WY�����N��TP�2��i���"� ��ɺc���#�'v�W6���� 2�<�R�h'!3���X���� 1�WDߜ����;;E@�J�u��8O$�탛K�d��?=�l(��:g���q=����P��j�4b8ZR��X���T���(�+�7�̢��5����fY8�����ȣ0o�8�H�!<�R{4��m
��T.�--�v���
�xU��X���_O�pi"f�9�\R�N��]Y(�ێ
2k�8X��ӡ\���8���I]Z�j@6����Mx�^�Z"o�*c��7o!߂��$34;��J@�Y�Ow��A� ��Җ8Jfq9�?� "��ծ�E�����rbC/���1v>pl
�r�`�ŌόC��S|�L-��Ԏ�|�8�$�v�sH)��d ��D�9E ����.���_`Ⳡg�u��V��MsDh�`��yz�koVmVf��LR \�«o���9���d�/q���,�}�8��DzJ�{I�鯩N-i�F�:z�r����ܛ*[�H�{�g𤿵\.HV�4R�7�0��ެ=^\8��6���]Yc�}B���`��d��0}(�+�x<M��7��:�F�C;��S���f�^=��!���D��BSf�]>��������D��}<�g�*�!f�˯�b�\U�=y�l�E��6��/b��}�y0)���V�]���a	j��m�O�N������3�����e}�ռ�����6���[Y�s��3s#~�4�Y!��j^�S��M9�`������#2�F�+�[S}�f����y�~{Ī�#�����6��R-��=Ԧ	^��Ucva�����q�6��EC	��zw��Ir���c�`;iSp���G���Z�F�DpmӻIQ�;�-#��۬߅|W�1&�O7��+��z�=�٘�gf�N|�����,���؁X������4���*V{�L��.�{��R�����B5L�@S�z�(�gp�@��{���u�;#�5v�H��_�ȥ9��v��R�P��⽉��l�6���或p�m��JE��;q\�� ���1i�a4�P �����fOi��D��"<!�kZZ.ϼh�].��T��_#/u��i^j�� c1���o��bSU~gӀfޭ�3]�}4�C��b�&o�T��&7������f��n'���wE�(�'(W��bF�m�q൓��N�^���oK��ƨ���=�}"vf3'%v�1��&nݻe��*�}����\��ީ�}���m��c��I0K��Q�c$�$�lnC�,֖T?��&Ӛ�^{X�<��$Q�j͖��ȷ?��2m�I	Y&G�~�A�4���g��bwnXΦ��o/�Q%����$�d�",��x���@��޺�r���sQ�>N
w���� Z:.n�d����}#�R����s%�(UJ���We��}�~9�ߩ����^��o�䠔%8r�p�yk�üK�<��Rl��yn��@���SmN���y�h�!Ybp��^�/�B����>]�b88��TR��*P��%��e���BQw��l���:��_q�N�V)���\ф��7�!T u�y�.iI"�g!P[l
��v�v}���Ys[��"�~��M��G����F���Rl]��P�oU�w�^P�\��.
�{��}�;��\�<7,��a&[z9�N����k��]~[��3�%�M���@ȼ>�U�m�X�1��$��d���8#B[(���S�� �.jb������6#`�;�5��r�j�]����]f����P7����Hj,Y|�md\
���AU��W���4W��S��h~���
�.J�4�ӻb^��B*7�ר]��m���L*_��A=��Ľ]>���Kje'�ё���/l�ĹԎ���u �"��!��o���k� y���-�w�i�ۍ��f�a�V)�R���4?��G"!���l�OC�_�CA��p3VT!w�Nna�oE���}8�c�<��uͧ"ep@a!�x�:H.w�ح[�3��D��p0fN趾j�T�K^65Q�9	�t��ά�<���~$��a���������=}�X����{+#?&��w+[�B���c��x>y�����</���ỄNٖ�ʸumϛ�X����ﮍ7R-�b�M�3(xʤ�;���7��2/�ه@��?
�����zפV�_����I`������"B�^��1�n.�=���hHC=�8{q���,�X�����1m�A�U`~�˜�%j��8��8��'W�s�~����S�Ȧ�g�~�+�k�C�i.�4|�"���+!�����z�5�F�W��'��I�ɬ�Y��1ʪ�J���
&�8K��!�x��^�B��t�[g1��3��p�F���/�G!>���~|�Q�Fp��e���X�25��xi��՝ѕ���C�]3���R������9ْ�1ui����Ų�T�@_�~��`�j�B:�΁ɻ�uϏJߋ�z�Xz�~�"�<�ޘ����S�1sz�bY.�X�3����d[x�s'J�X���D�+jAM�谝�A7݅+2iCG�>lT}:@���yY ��&d��#�;���hM,j}{��S���Z~�F�
fhÇ6�ȯ�����h��KU� ++�4����p$W�Zx�#?�zΊ���шT�/���${(�A�ʨ��Ѡ��u8k�~��߉�,U�-�<a(��=uF���aHf�--�j�7��b��.�?q�-�pAư#�ъp�ْ�Գ���A��9����	�r�|��oY�#������J#�>�6T�4���{�K\
�/�; �b1� >����h)MqɄ���?W��>uf"���}�����aK�u�B-c���e^N�L���̡6�C�O��Lb+F��u�z�K��4�b�B��Z_�����a��#3�>�Q���S�" q��@�mw�/��%��e�$!A�(2z��'+��ժ�c�TC��i��X��1���j����ď쫄b�Ҙ֌��)����I_(�����������.���/nl�XS���l�p��u_�l���zw\"@{���3�5t�^-Ea�t~	R.���"��v���{�Ջc��Mq�Տ�(�5|�S�
�U���[���-Dt4c5��ݽ��7]�^Ԭ���#D�y_����ы�?c��7Z�*� 	��1Rt�2��W����&����$Z�SEdsJ[����߉v��T��X=��#N}���q�N�Ko[=�%\\��/��IglV�_���M�;*+��*��!GVƅw��ӜY�&a��Ұ�]�vX����^��߶W57}7ܭ���?������i�.��1��z[�3  ^}`���J�/��a�T�TB���M��N#ܰ��s�<H.�)>)hMzfǩ;��g����>X�j
p�w6�J,+��B�4*�f�3���⁇Faq&���5��4>�g�$s��_�n�P��29�ȹ��p˜"�W�+MςK3����f�bX<��+	�SKu�1@��!���m�T�9�F���pu�v+?�do,>�]/zz5��8*l�Nlf�L9�eqj����0�mRݕ�X�%j��o.2@T�~�B{���7S�G��톆t[Q�4D�����z���.���,������-��a�bV�lj[�t�<Ƀ���;�M"�!z�>b ����1�~����y)�i�D=��� �V�}���Z�ۊ�
��l�#;v��iq����i?����-/0b��߷�/Z)GH�"% }��{��vw�r(���[$����m�ؑ a��}u���b���qb^nh�;�*r;bl���d�I��w��۸���}�9���^O\~:3]SQ2���������՘�7y�b�똑�x�$� �h<%lRWK�bTfZ*	�X�oQ�vBqeJ=�%Gq ���r9�}Ҧjm��`�%괪��V$>��џ�8H������ �l��rF�yFi/���l�����S����&w���v�jX����>֐�<�H��� �q��Zٞ�����Y)�J
���.�h%Md�q�,A�$e�2�H�8C]�'<O��`a�����W�d���;�/&�p��ݜekK5A)�<�/ ���AH�I��%,�!L��
1AX߈,끔wܢ"߾�36.�C���,�M���L�q�$�a/�vV��#Ҳ�L�}�z)�N�3⍱vR��LQ��N3����A�m�T����>o�dyt}����㸣��Ѳ�� ��*�T}��"����z�NI��pbİ�U����e���i���};ot2�Ϻݩ����z�z�̉4��x:֖�G���H�z�^���S=ځ�o�~Q�8������LS��˕v��z+t�;�?���m�B�(0���:�S\�ס?�:�I'��\'&OS7�F'Sþ;S�s���.���˗8�;*?���D�<v�RW�(��ܟS"�������C)��Ubh��~)i�Y�Vi:��ethG�t�d���9��'(���A�-ty�;saF��W�PX�.n[�x����媎�^c��~��<rqJD�Z��׀oC427��m�>:S�i��q�Y�b�ISh۲���+X��j@�3�7dl- ����� �U���@M��Z��$jM/��889v�6k�ϳa�$+��@|���A_B�ĝZ����$,�/��w��iAg*�ƺ1DSx$Ғ��7��C�5Ϸ�����3D֠�'�mWLV�ky�Y���~�\r8��J��̓�P���(B�<�*���~7��]��=�E�&Y���d2͏Z�vF`iv#�g��1��D��2m����K��U��x�%��ڦ����	4S#K��T��ˍ.��
=�OϺ���GuA��&�rN���V�}�u������IjB�aѸP LBX�wU���:s��lw��gB�/z���_UՑ�i��X��1E����"�C툷��\D��Ӆ�&�?�n�"���ꭳ�K�&��d������~�L��.dv�&YPty�`��s��5>�-PE�D�-@�塰F{�C�o�O},7ZJ�ϧ*>���*���