��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�؆q/�֜9Y{/jl��:�Y"S1�pck0k�j������ ��.)�hj�$��v�L�����"�pa�B�f�V�Pa�w��|�a���yя��:{�O�o��\uL�����ɶ� �#�蝢��_[	��1 �q�U�A�x��)]O�~&tk��f��Η��}G��f��}�F��{W&�U�k�ގ�m\�Uqn��Ɯ?2d���Y'�6=�S���M�Rh�⟣<yCh�H�<�q8m�ĉ�w�b+T
`a����s�HyP�.h�z�:�?�q! �8(�x���-��Z����?rc��O�<�{Q� ����oˋ��%�r�Y<�m�r��`��	6S�"w,��J�spu�J嗢
%  �x���77��,��U�W�K �q�
��DF��R!;GY3���=�\�4��1=N����[t�D�/�4�ծ<}2���ҩ�(#�(d�yw~�K��Z7�=hYbl�G"_���&Yڨ!�]b�kq,��o�ʹ,��U�
˹7Y�
�ue)�3
9����@�L,�;ʙI���h����;����F�@�D����xF��������5���Pc�vH7偑��}�Y�(��XXU�^2P����Ѓ�5�N���,3
8PB_��l�t8ٙ��Wv;u^��=�Wpe�C��t��Z�6��zx�f�6v��@� �ݕLo�u�+��6� !�Š��i��B��d��E��O	A�%mCvt�~$���Q�P�W<K>��eDU�����y�}��$~���V�Y�w���
s�_�m��ap; ���	 ��H�����c�ԏ�$$�s���?���񱕼�����F@�`N��C��4��6�㹻� �[�]����H���i���j�4�\c�;~�sr�[�H\"@��7\t���x�iZ
���+�����o�x��^&z�@ӳ8�@�Ӑ�T?����=��H�#�.��º��J7oy]�t8o���=-=��D����Ű���AG:�Yqo�^�U��^ d��2�U&��<����_�c	0�������Q�ue�.[�Р�n'��fk*�/2Bm�NZ%O,��6%�_����]�0O'�'3X�D5,ꨄ�g��X��O��<#4	�M{ �MN?#Q�
t<8�w;��W\9����Q�����x\ZMc4�䜅���b�1��;��K�,�'�@��ҕ�萦�<k���K������
�*��Bq]�x��-�5�������e��π��t�K#|��T/�T�P�)b;7�
��?O�m��������h,�̌o�E�*�,�r�~d�:�9��vT�T�>jmD�Ø3w��V��B�w��p�J5H�zjnE R�h��2���s�ڱ��	g��?��FLM���$4��i�M�q��c2��{%�ajd���uD'|��-�ޗ�-of��P<G�/��=���>,шï	B�� Z4�D�.�`蜬	O(�n�(@��jʽծ;s���d.M)-�:�i��7vjn,l�hŚ��y�yE��V�����F�CX&Pw-���ě��L;�I�g"ު�H�͢��}u!d�dY��#��Ov��\-�nk��������<�@�|s��)��"�;���_<�Ξ���1<+SB�9|�A���K�/V]%O�'b��s��c]_*��L�&%~G�Mb�1c_�H$��;�d��S��dQS	�6�|a`�C�8֖�X��C���[�ǆX:q��6d� L{kj������w>l�G�c��2
���^��W��/jǳo�g���(�ZτɄI+N:B��7*�Ӯ,G�Ϧ'���;򸧵����ר�%���!|�5�K���e8]G�Y.4 �$�疤��R�y\zJ�����S5�c�A�+4���ܓfϟ2#�X�D�:��\J[�;|�m��Β�P�@��9x����؝~��tG�����4+���K���w'���U�8�2������3�����^ˇɗ1��a�t�v�>�ͱ��˹P�;kwo�����%���?���^y����v��
װF��R��n4 �|A�h֖R��w��$��r�1S!^���R��( M �Z��-��ô��cp�)�#%����6(�8�~�i�Ts��VB	H� � s<XQ_�eb��'�VXҼ�D ��H�P���EL���nhE�?!o�:�v��4iMO��[VM^:��ثT}�=����q�;���?$f�`��P�ؙ?K��Z�k��`��TY�zsuޘI1�"�@z�I:�2�+�����F4���ݵ�L������m'\����µR�0ut�]��K߿kI�r�E?����?Mo�x�}�35E�w��F_�p�7;q��� }a�m�\7��@9�UH,{��t���V)�����O/19|�� ���$���7�p��+����S%�4��Y6hx=WN�)�P����"�. Y���� �a჌`K���w}�f�~���v�t/���m�Y���������2T�}]܏⒠��<���4')����Zm��I7z@�"�xNɆWs���o|�R�ϤO[������D�����B��]RѾo�ڢ(v��i�H�3�+��+���<es��0�= �G�%(e߫ti0�R���PtX.r��]l�qo ����l������������C���Ԑ�Kϑ�)���u�wܚ[Uq�D��<Aj%{�;���s��|U(C?<�Yit�}��(��g�mwV��>���A͔�j���#�^�A�W� ��4��Ȁ<{��;�,ڧM�m�ɧ���$_e�	�ؼe�_V��r�@����߉��[ ��\ή_"�Ύg�K����L���lr�s�z�+�y�Z��ʩ;ً%�s�,�|��f��p3���p���ʲ��~���,�R�}����DH���˧��gNc$a���`�v�]f��W9�sp��+�����&�h�d�Bܪ�hd�"�� �&�l��0ՔT =sT>T��aG3�}��ђ�+�I��ƿ6��"c��\�yp40��E}X����ӄ;��&qӤ�X�9�W�y-Ϡ5Ŵ�����.���P��I��$�dF4ەdi	��:�Y��]��yT��w+~�����F5�n�ð�g���(�/L�q��G6·��l�فM'W�1ʸe�x������CmIٽ�f�B�7����bۻ	��
��Y�&?�o�t��/�ܥ����ꊋ�2�I}ݥ�Ln2�~$��_:��ϵ��"�w���	�9��6�������G�{�r�"=P�H~uc�7@�����qG3��y7��1����H���w��H��fS�~�����O.C�]%;x��؇�sm�!#.�R�W���2��y�v�-}��κ`wbwM-�s�L�"��r�C��#l�S�76����9
�&{4q��ά�f����_�@�mb%��=��
�-��l�i�V�D7�����"đ5�@�\�Q������Up@�rî!��]�C}�,�Ը�u�u@����}a	�x�qB:d�"HB�t��7�E'aH9�c�ŀ�A0��2�-�@��(���	�߷�n��~�2D@��`��L=�&���&9[C����M�����wn�e�Ry�����E��,@�!iS��zu�"0w(�4��%-47�;�oR t�3�A��+q���Lr���sdt�9k� �Nu���u@��0q���M�?/��w�x����2@@6Z�;�Wc��Ǻ�MeI<�x �\�M�z./-�"�pI��&�����_�������-.��i����^ړVZ�w�ڛ�G��O�\�P7���WV:l��)+Mo������[S��̿������ޅ2����V���wj�_�2̄y ���z0 ��bfU��v����m�P���+M������^��EZh�_H�����U��L��	��`[��[<���/����M�^If���Z�%(�>43W1���xn0h�jÜ���	�3.K�"��F��j�%�:��g�M��[�X��
�yD���Qwl�ٵ��>[���D��^i�L��Y�r���{]�
���6�(0��

�H�^z�m��Ri�`�(��q�,�ҚIk��q���T��&�l�y�^��ڜ���@�|��
Ȝ���m}|�[V���j�}X!� �s���O�@u�oO0�sؐs�����HJ:��>`=�����{�Ҍ�ܚҏ5BT{����'�m�PM����d��yr����}�jy��ۊ��Ǘ�>U�$#���5�қ��R���N�{UP�y퇙?.(OY��R����6���8M�����52D8�8 X� �F���Mƿ:���=��Z���x���A��&��X=���C���sÕyJ���]9���|vY	��eG��H��q��4qKA�jXV�+-�j�v�7hĖ���/�������+_���K|��WL�d+K��}+[��
����0hu3��^wO���=_=ڢ�S��^=���Y�;��y�OE��K�q�K�Kc�����,)̀ÖL
���������Y�u⏵{�M {N�2/���_�M�.��k�q�2Q(�*Ibt�r�xr�ŵ�6�"��1Ye�ߧ�e&�c��#�'�Eܩ(��g)�,�u%F]0�;�ȫKG��N7:$��6pg��sFY�7��G�$�ک7�%~�����t�ey�k7��~I�bY�?.90�׷��v�+ t�@|�O&��c�t�e��3��� �s��=��d�i�����yo�5љ,�&ZR�����&��&9�5�m�p���:���f�[����X��/�
k���Y��*R��t��+������?�	5v��%{��|��b�Я�u!�ĭ�}�����M�N�"䎁 >�GMN�����xhi;�2w�_ת=u�B}ܯ��
��OCo
=X%hqX�	i��Y�"�?50&1%���a��4�	
jѽ�򁔭F��W�}HAR����Y������rY���5��b��@z
�֩fY����y<}D��`3t���j�抺�5L��g��-�wn(�*ڐ�T�xW}��})Qr�h�S�(�U $�+X��/��Î��%\��7!_hU�'7X��R��-�H��x�8�S�d7/vޠ͸?�7(\�Ӿ��g{���A�T��(�{M�M ��+Q�>rQ6�?6������J){�O�_^;��Lf�Zs�A�-W"pK��ۈ3x�i������e^����#2�`
gb2}zt�`
����=D�r�b�P/��y�6��A�3Z�(ĂG��-�FI��<����t��0]K���J'��*�72�7�v� g�a���@� �7�A�����q�p���6�F\#�����[���$9��ᕻN��Woߕo�s1}h�G�5��c��m�W�.۸�_�KdG��Lz�c�I��էTz��#��S�7���ju��g�%3��9˞|����`�e���&oY���?E�Z2�`9��Zc���.M�����f��,��UV�~�K�g�S�p�����fΩb��g2��퀮n$˱	�m%��I�RUnj��}�&0m��Xnc���,���"19�_��Emؗ�0�hЅW���!�Kt��OwH��a�~�U��~e����ؼW�~%-}�f�+t(J��W����)���$<�GRƹ�ŉ�*N4�:!�K�J�S���l>I�`3q�.�;��{�K�K���=��v�֮u��V�H����5]%��I 7t���6=���*X�ue6I�1 ��C3��\>�d�9�=R�.�]��xE�� �"Oi�CQ���`i�H������j/�A��Y�d �MO�
���&0�~�����2,�����0���&2����,��H7C����`N�
�2z�tꎍ��7Vi�H.}��.q�Ғ~P?�Ԝi-p|<	e�A��+<�{>��X6������y�*�5zn��9̺&R��qu�-0?+�g�L��8GX,�
�0�2�z�xD$`̯�^ӣ��7�0�.���Qo$5j����5�s�od�ɐ��)1ޞ�J�8d�� 48R���#,�Q�X�M2�΍�HB'��+�-�)~�zK���[�"C�d.�b8cP���K�$�?W��&�sن~���L�퓽�{�<l'Of��y��.7u@"р��
G��A��
9���	f�Z�f�ҕ����u+3*?�?����usIs�m �wQ�̨�R�����r��?����N��8x$>�)c6ѣi}�O�뻭��PZ`�$}(27)���)���}�����e��O~�[o�6��+��G�|+Vs�]A��cd���b"s�w*��u]�� ,����t���t��+N3,��Uā)<Oe�V��ݠ�B#�vv�$�R�P�K����87J�=P�%D<���x�W"3�`��6�/w�n��I�D���1���h{���Rq"l;��C�Ӥ�6������Tx�G��NS�5偗�7����S� �.$Yr�D����������G���/XDY@7�5A��yD����x�B�oz����	kD�y4^��{e����J�'i'������+�˺���V�2h{�sL�O�(���BG����Jx`��^v03��n�ݩ&�<!'�����--(j#&��-�)_���B�sZZ�Z*O���FXW�Z;��_��B�t̔ӁE�W��̃�s�i<�%/�"A��Kqr�z�#��5�/T��U�D�CC�FDp��,��K�C��+��&�W����6&��w��)E����E# �_1�vϭ�����|����]�Q�����_>J�]g��Ҧ�=�J|��(�1�ZmL��ۻ��/|�ψ��w������Ux���1��'��qnؚ�������*M~��#�j$�K�l�*������'\2�����ƭysc67(��0��Ӏ��n�?z�q\{���,����<3j)k��b��n��N6,"�k(+f��l�	�e��@��r_���p-�̎Z
���d�P��9c��*O|@4��T�J&�1��İ�|�%�*�cr�f�L����?>��H8�o����f�>����])T��
^}�Wʶ�bٟӘ�+�K �U�rZi�F�'��7�&6+�ϓ��N��GH�W��)�CTG����ܞ1���zv�7È�zn�9A����L�%� ���k��ġ�*4_Ǯ�}��ق�wW
���V�V�-�t"[�h���0�VwJ-�y�M�'�-/Eʪ��sR�Cp՞�G��Amq16`�noM�� �1 ����AyH� ���M�,i��l�D�`�F�cs$7Ha����?~��t:k�a�"(E�Q5���4=�%.8����Oa��(��'fga�e�+x���[S����ZQmÅ6�����{�knS��blx��1�{E��X��L��^}�L.�ڄ��U��1�`X��7�h�;q�� ����)����7MC�Ӛa~�x�Q�I�l��D���	�,Pu��	��+L� �aU��m;?x�#�1��k�/0��Y[dxbָٕ.�K��ř��@����H��M�� r���z�_戳���{q%�CH~�ۼhs,�(�
qPt���0�=��*��d�"�����ִ"&�
���J~*�B��KE��2��q�z
1�'�(]�`���|�X�1%�7�4g�X���� �r�J��y���,8"�������-���c�I�*I����o�~U��SϹ�S����z.ghQ)�� ���Bj��ȷP`�˗MT�:�7)����~-��s{kT����x�V<^�rВ:��F�?UO���J�e���'���{y�L!֏E͓�`�׼����s(7�n��_�F�1Bf͒�v�K�+�(���ߛL���eJGKY���iQ}U3���v�Y�BrOs���f97p�ê��a679���d�7��S2�>�����.ݸmnz+��XrM�P�˒��=�s�>�������؈��
Z�(���,VޣH��4`�7�a���v9�����o�%��2ӫ�5���I�'q��]�*�9���*�gɊ�'lq��C�2
���sx�G�r_�=cx��;����;T���P�5�[0�Sع���;��X1#$�Be�qA�Nȱ�)o�2���d=ԣ�����Zxz^�q����������P�+Q��G��;3���~g���eZ�Ɩ�者���A[9ĭ(�R+�h��z{u�-����>��<k�S��A�����7q�w�0� �E^�6>�ډ��(�� w!mڲO�u�����'.o	{Q���_�Jc���.�wU���Bjk��;\��w��+�f�"��mn���W�A���|��@�LP'�N�b��m���X�S6�o�"K�3ľ�ۭtyu�y1rd'�����|�l`���-�<ƙ뼂����`ͫ��џ��W���h)��U�V.����LG�-ͪx�QJ���WgL`�@�i�7��yhOL�߾.�*i�&����Zb8�mΣ������/�⏡�����w��<MO�"2Q�v���ɡP�$�i5 ��ҖZ9�?W﨎��2C�p(�W�E-�3���4h���*^CV�Q�_�G��׍~?Xb��Lx��t��� i}2j� %hV@�7^3D�ޭk?�Y���:RâL�!�hL�p&�ïp�߫���`iTCS6�X��̰�CϑF�DU;�]�UR**t�"��7 w��{v̥A����n��|,jK�"�.N�*%#T�X����J�9�d`D6dASaH�rr(,��<���
{��;9�S ��Ψ�c|+�JC�u������$e��:�f�|��b���+����	�J��w��%u�~�Y�񗴒���q��O�R����؈']�������|���g��51�FdX�ޔH�h�ԓ�n��%J��3�`�~b�$��}s�&�d3S)�v[E{��,u�*1���-{I�f��oݮ�~L� 3�jcgMt�'�h��^��鰴��1e�dP娯�2�Znݮ�Tb�r����LV��uK:u�k��@K�H=�q�D�"B� �k��	RLt7B�r�t��g�X�]@�ץ�K<���)��k�"�~�5UPt��C.!�]V����� aq ���6�t����B��}���:��#�Lٿ��򸃭�b��B{�+l����Jٹ����*>U�cϱ�w
5�69��]�#d����}΋CI�<�ϫbl�[y��m{(?��m��:�8�or�З�W�.���t"�#2����qK�(V{���ؖ��e���i(�F�F�#��x��l�9C�;,)f��
��g���Zy��^�X0W�
�������F��� �<@i)�}��F�T�o��k��$�S6��4��i��=�cu�b��J��S1��q�. X�3G���W�Cί��d;B횙��CI�苺�A��7�s3�h����xc��n��n��i��p�'�RF����ECJb�Ld�0zJp�tp�c��/�7�*2�'��3�ì�Ŕ잩T�HI�ϼ���ǯ{ ,�{rj+9z�O��b6x��z�9����C��t2Nv5PYxz�T�U�n�4��3���W�U��_
�܎�w���0V�0�@�]f����z63�R�]6�9RZ�v'%��}�!(�a���7٧l��9�?��r��z)?�2@�C�h��7�K��� �^GS{���e����B�6Dc������k��%�C�PR��U%}���l`���j�g�aF!RrB��m6�b�}G��aG�׍�)���
>��}� �'�i��L3���'�:28=���q(Ʃ��� HG2���߹���@��G'/�6w��u�3�
��0��1$ӷe�p<�˨$-�/��:2��[��Roi����ח٤˻d���.��ia8^�c����}!L3�pOW�y1�ՒLx���a;%��tb��Wk�seAuN?u3����9�ud��ݝ��)�9�c�7z!s�c@y"��<��� ���9����ڑw��v8��ga.�2#V�/��뾢�>��˸R%Z���s�h�޺�ĉn��tI-��@���9�c�i5XS��[�4f��n-;������3<N�eFa���
�Ҥ��> xk�ϵ�����f@V��YT^�w��Č���CIw�ˡޮ��(P�Y�W���i'�`{���A1�%��	R4���m��a��s�'䂦���_8�y`6[�z��1����*J�ү����w�zϖw��>�F����I"D�04�<xEe�7/��l�.ەm�'�u"�M�P��+8m�D,; �0�d�<[�w��ï2�+�|��X�L#��<��o,ύܵ�9��]��@������!��2���]'ً�6ۛn�����[
ʇܯ�W 8���i_*��6*��8����������ȑe�1M�5a5����S��<c�}�Y|�]�I���I��f�XZr��0�5�.&������*9)�Ȁ��k���ou�(B@W�o�����T-R�Z&g�'�~��9O[٦�k%�n)��?5�l���:\�Q��Y
[���eb�b�S����pHI�(;p9-�B�*B�RL�"LԈ�l�|80��n�R�JZJ�#��R�5��G7����W8^H!XK$bz��V�p���s�C�@�bN�Ǯ����je a1f����՜�'�k�n�� � ]��tk������.��,��Q��B�Mq3�9�*��;)�҆Dg��Z��o�b-�ҹ֗�����E���j����Թ��4�ŨZ�
��ѰS���?�||'�m^�	Gq�֥Y1 _x�N6f:A jW5�ډŋV�/ʎ
�B�ܭ'϶�F5�٧�&DBv��}�������l�
xCf�n���5��T��7C3.�^^����r��.�����k���Z����^�a��jX��~ɼ!�XR�UwQg�'P���,��"��t��_��}�|�+��h�x	R	7R�\H�R�y���ZYR3ơ�*�.�<e2�>0բ��֣�z��{b0zC �%����qz��d@�f�!�fX!БY��Z�
z���m����&g0%��t� өhV*�Թ�L��
�[2��TY�:B<�ǔkk����	S1lJ��8A���r/����bU�aK#�`�^/FG ���k��4�f�ݟ(�Y��kD�7�Iǌ��L����JD���E�����fϬ�DT��&�����=
}�<;�-WK����r��vΩP&.R�mv���<����JV��?�U;�@���\�*=?�Ck��i�`� *Y�9�=ދ�������ԙ�	aψԝ�"7����q�+d�ݲfx�O��Ұ�g�
n� �����'�N��ޘZ�D����q�[<8[_�&PFdl}�/w�j�iO[���!C�4��C�la�҈�mvv�6L+~�p. ��� ���M;<z��މ?��$�paE놨a'L	��P�L}��87yʧ����'�k�d����D���$�ٛ���~E"�\s�
e���x��+߃���1�����UF"���ߨ��cn~�s��k���t�X-H��	�in)�6c�����i����3\�x���Un7�x��#�`EjK��K=�b�����SɈ[3SF.ĖC ���	r�x8/�3���ڕ��?3�v�Rᾁe��T7b�ױ�!�����xK�K?�Pz{@�Nכ<�h�@X��'�C�/�>}CW�HTp{�e{�#z�A�\a��g$Ʋ�my<g;uXY�Mf1��>r�������^����pO2�D:H_L{�&�)����FLY����\��ҫI����Z�e���g+/�n��o���h9���f�t�<j�M�c���օ�Z�ʟ\��ע&�k�x�B�/ƽ(���8&��?�T4�(on�K�J)M���ΐ�P�񏤄��t_-�>�k�������F���,�f� <nVXA�D�M�5���gdH�s
K\o�E��M��:���!�1�����h�	���n��u�^Y��a4��޷��yg/X�_c��c��QK�X �)<�tPjcO��W�*�����/��l��`���zO�-&bJ݃8�Wu>6(�\:+�X`;H����8�Hv��yM�C��{r�N�ܠ:9��h���6  TY��PA����y��1H�%��}C}s��oU%��sLd��i>ja�M���ߺ��?�X�����5U�.2oq:�Ŝ�W�Q�kО:k�h*\Y�"?]!��:Jֱ����/���-�֏]Xx1>�ݳ�ɩ�M!��S,�ӭ[H�,����6g@�I�ϑ҅#�E������	�$�#��ǯ;i�;|6D5�wo�!:]۾$xɳ�ůs��@����a����� /���MS�����������<��������-j�J`aL,<���2I 7�O�-K^2��;#��I�̀���ږ�"�5��MA�V�,e�Z�&>@�����.���%ݷȗT2�ЀDO��bikJ�s{�tYtg�gm($�6�?�mTA~&[*De:�AU6�)g|](lAA���p)�[�mӕU�duMF=�����C%�YD�5����)Y�#��q����^�f��>��H��Z���6���E,����� ���$R��J�'�@O�P{�c]QE��҆�������FZ��tk�h�#.�ԑB�F}�	�|���Mo�G<%gtuA������П���!t�.+��F�����L�����P�dV�h�TҎժɒ�|Z���뵭:�wz��$��	���<>����$]���������5�����Gp�C��C���f�fA���_��;v�V^��Y�#JX���3�B���%����ʭ��<��I�l8[�+[6�Q/٥�J�=���e���UP���P<0�=E1�^CѲ�H���m:v~PU�ÿ����\��]|U��b�K��b*�𲇸��f��x۱Z�N�Ɠp���)��8��* U���2:�%���-NI�s�K	�`y�3�L{�j�^И���@k�a�!�H����}�� �����V=���M���������)��aqK����������'$k9K4�����=p�HurQ`�D��ԏ�(��Wt&k��_v�l�OBFM����h���r-p��`lLؘG�w��L���r��;�.'��p�x��`�R�~�F#ꭻ�~z�)]���Zϣ�!��rr�'!�U) P��n��"B�kR�{<�>���D�#$�X����m��ZJ��2 �22�0�����q^��!#P�^5�\n:*���x�p!�X����-S����F"�X�V��xr!N5�ͤ�s�f7=�^h8�à��I9,�r�49�LԲKWL/A��#�,r�-Z�-AV�ԁ5��i���&WV�W���TQ-`A;��(h��4>O�dn���N%nq�	�8�ԸP7�0�i'"k	Kh#�Կ����M��73�X�������)+d;�w��U���>���^�M�V"I�&���"�|�k��<c8�<W!y�e:<@��B���\k���bV�O�/  ����@|�%�D�}	~�\dK�JV,��r��c���+�����T�����[e)#2�$^�%E���aEW��&��M�v��H�E��on�#a��,��>@�%*j=�W�CC`	o ��s:��Y0=U��x~O����8��_Yi�?�Z���O	�=ۺ��8%7I���0�
�`$��@�	��L3 ������1cq���[���$�f��B94AaA���Bn�%�s�E�kWh��W��6�Z����u�k	Cd�	�9��?3$?��;a에nc�,�V\Q@�A,K�A>�^��=K��hih]�m�9F�7;�iDBޱ4��^$3�O`�G�S�ʊ63��uaWM����U�N�K�0�{[�@�`Fo�M����B�����]�7J��D�an�2�y>ip�ǵ�Pm�3��|B��7ԛ��~Ϝ���92V�X.��<�W�l�vQ����N��_�٘��Ӆ�����[ �l7�J�~U-y��$F��G���D��L�n�Z���˯�;�o���S��'xR�����-�S���^;�1�� a.�#����Nz{&!�>5m_`����?1
T���Z���X�R;V}?��F+>f���W�3��{N9�x+�������%9z0"�l�>�d���������|�gCGv@�w���er�P��^���X����O�N=�8��W��3_�Q��桊�'�Y��x	%}�|X\d��t阧��ʊS(�u.�d'��j��9�6]8��{We��j��%�v�T�ri}t=�r�bw��31
�u�0PY�۞4䔱��G�i귕��P�י�i\�m�1�S��|`dc�*@�\�
 �-2��ͬ�1�N���Q�rQ 4r�f�sܚ"�s���D$�Io�$�(������ME�\=y`�*%����[Q��5k𰫲�8P�u���'Y�\�b�|{�Դ��RV��s.'z�ǪϡE���;�t9�*�"'?Kֿ�dR)IS���ң�ා��S�1>���&�_9ͤ�@Tj;�a�/-�@�!k��Ӝ���1�x@��m�*��ST�e�l��������r�Ɉ�}�y��$�l�qM*�/o8��-$u>�*�(a_��>�΍Fψ�1�#6�N6?�J�r��yO.��;���&��6�6x�oܒ�T���~V��'@�ɿ7��ڐ�2����N��{.���<%��"/g=��0��x�H����Ӯ�1��"��=hq��m�G��Iy�X�B��-e޼d2����h#CjX�0a��n�m��b�k�C���{ϕ���_A�)��K��P�#�ƶ�(��i�A�?�C��qd��� ���=���Ab�xh���)L:��`�g�H�r�>�}���(I5��rD�L��$�ڭ��3�ԈV���2���2�˷Uf�9B錬�;55m ET�'7�q^�[�E	z�*�fdE�Ò�>tۺ,�߿�
��|6��眄��s�,	��i�aw��ڹ�#�Iv5�}:�?��$E5�$��Y	��p�R�)S}�E���᡹ZO ���*~h���7Q�t�������~�En.y�T�|A�"��2ZݍC�(y��m4��]	��O��B��4�?���44!⩖��Sz�j���߯�tuI~�K�	�a�K�%��lE��%[[6�M:P	�چBCr�a�{�m�v�S�D�M�x',��KWOc��}P��`�gD��S1�1�OA`T�3��@9� �W���
)6��>���hX���H�\z���S�u�,�(��Pц�Q�w*FK��E�5g}k����\�JI��Е�tw.�`銌L��������ӈL>ˋ�0��NE_�."��;��Do��9?+���ny*�)�>۟���mS(ǣ$��W��r=f;[^ �~L����+�B�����&z4�J(�E���[55���(�;���(�x}������q��{�ܹ�K�9�"D�H �K(�Y�3{V32O�dLi�dl����C�{�C����6z��]#��C���9����۝�J�� }q�	mҚ��Q�h�!�g�'�� ��Ò�X�Q'�����l�l*Lg> N	({�:�*zsd`KD�T	UjN)�0�v��-	��n������Ƃ6o+�� �B���>?C{�����g�:���㘋�5y�� ��C!u�g@D6eә��b��bF�!��2��s��m~��-�l8\�R͒i`ɻܖ���( ^0@G�~K��g����.�u��;nf�\��J��Dek�ݓ�EK:͚�xA�,L�>��8?��-���Ot2Z﫶=�մhH�t�vr��
sOЛ{�Gfޮ~-�
�Y�dC9�B��ݳae�I�{d7��d1"香̓I�,�FW�4�3A��~K�z�n�M���K)�@?o�j�J���ِv�C��e��P��)�?�2^��@����O�,؀����1�(����Jh�A���$:4P�6��i���1�iN����U
��<qv��N�D$
@C>c�<�(�
�W������^�����pA'.���f���kg�ڟ���
���4��[c��4���7�N�$�e�4����7��$V�r�&c@�//�W�j3w9����+�3�ؐ�����K=p����$����z��[��?݂� '��V���'[�p�v_�U�w�2��6~Ա��]�~-r�!������:�X��j�P�8�jg�y�2����C���h���82�	�7�F��攢�[0�%�w2�L��_7j�A��U��[�gy�d�4[v3IA�J�'vtđ�>U�G��H�0rFH�tK�Oi�I�}c��{�&����v�dفD�ZR/w[E�oTF �[f�y�A�R��l�3���N*��{\�����w�4�b�T����Js9��]�/Z�Q(��"�R
������S���X�F��%UaH�j����'�^�>>����~;�HwV˶
4�����v�?�Q�h��O�1i��su�����V_OR��A����(���)�/�fL\��K��e�_�����㤥U�3�q�l�[}W�E(�}���Ce|��c8A�9~�
�8�{��-(G�.]4�Jy��57���%o+���%�U��)���z���۳.��=��TY�Ѳ�'Ѭ!̋<~�E�g�ʝ�҇��^O�7b��M�>�yㆍ�]�-���$�Y&�r�����]y�Ƽ�w������nT.;���%���f3�k�V�jP=T��+��]��D�H���@��L�S���-���hWZy�+c ���k�!i��;��YK��n�O�4\&WZ'h>��II+r��P��H���BT8���f��2�,��d�ȬJ��@V=���x6���*3Q�IN����2����;ƻ��:Rih�a&Ư��u�a�x��R�r}���|���pc���F�F�Q��W��AD�s����ƜظNt6�Umh��Sא{�a���JLp��᣶��6n��E��*x�E�Ș<@��%����==8�aD-�)������	А�{:�hG%�oʡo}��g#%C꫔���`�J�R��}�S
�С`�2C��;�������2ߑ��"|W�F�hp0b4�*��R��Mo�%�X!F�7:ۊ��Ӟ�}�:��*1eS>�l_:�IAUP�!0i캢�ʧ�*�E��'p�z�çδ����KR�t��wʺqq�r��Ė`!�F�+�MWRy}<��3Z�t�> ʜ%kA�0B�uC����r��a1G?h6�d�2��Q'U���y��h��G�����I4ׯpX��hPs�5VXO�S���[ck�^����W����O�������o���^�c���G-��[ҳ�����D���פ���?1��4�����~���x��MH� �\d�;��b81�K�ڞDi��d�战.JB�@۝'�[�/����VP�S���#�NN�&�B�"��ϊ�-nOR���r���m�4$�4�D�nLb�!��w���o�Ƶan�~�7\V����7�~�F8��e]�B�[R[���� �*�_m�0�*���̻�vɸ1��1q�/dW-m���e��	��/��6inE����3n@k�����c��jȢ� ��o�;�4���$�Z�'{��F�y�	�"թ7��{\f�l��%���y���k^�\D't��N�R�z��Af��T�)8�� ��KO���D�*���z�� k�<��@-�>i�/|�����n����n�?NȲ<�\4��a�*&�4�QD��P�%J6m�2F�C�����il���N闱2y��ϐ/MQ�`˹�mwzL{G��0p=w����+���+4�A"s߈�'�>z�����B�c�Rb,x5i·��ҵ�J�E�w(	?i�75����ԇ�h�o��$�үW��X����p*B��&������>����j�;tmI�
Hi�g"�_j��~�X���)�6���y�vg�&��Z.޺{1�\�Ӏ�7�:[w-9��͈h� �϶�S��.EJ�6h��꭭UM�7n�����nl+�o�N�G��zy\k�����6�.xkěx�O�'�� ݫѣ`,��I.t�B:s���݄/5?��[���gF�;�=��*�)�kc3���㍄:=+����GZ�b>� f5�*<X�l�맜O�!d���z��rN�+����E�H���
������K@�#ƺ�����\��

�-�9!3r������I��xFZL}Y#�E$|�L<M` t8*�y'�ў+���h\��B�����Ԙ	��"�$CL�6�F��6�_�NU7\�B�Q?E`w͕H7��!�_I���R`�L�fg����а�~F��d�]a���:鵀Y_M�I�.�r�����!X�ị��������r�X_��å~�s�M����tO���D+��B��.\���}V�����rڿ[����]p7
О±XK��Ql�{��g�P����W!lPߩ~������Y0�6E/�w��P�O�j�j�i��Y{#x�2�`����d�=	�K�/�s��o�=��E	(�B�+�$� I��*�p�+����.�u"�fu}��hf�I����R�˭/��T�m���R��<��r�f�7��n$���@D	�Z�Y�L}/�L�	�P��T1LA
�DnN��I����3R;��3s�[�%V�v5L�r����Oz�~��8�ZNΥkő��ʸx�i�-f�R��q���*F�T�`߀A@6�q��N��\��cŘ�c��U�f�_%Ӡ��o�Aa�z�e2^U9m���sn��Ԗ~��-�EC$)C|�Q������ny�a�8�ڶ{��l*�M�v���M~�j��_��٣*Xm�K�Z��ܗ��]�$�;R�qM�H�o�㘣��\�a�9�+�LG�Mb�����*�J�BG�X'EJ��]�3�{ʢ����P�諸�띇B �gZ��>�+�>ԁ���8{d��)\wkpDÄ�l`����7i� �}�_[��Į���<�ݲB�W��w�����nG��)K񿖅q�N�%c���V��t'�%�@��W3�f���ok/��y�R�����F�<�����;�~��o1��j�v*mBٰz�6�y'(?s� "�yR�i��D+��+�f
���NB��m*;Cc���<-���L;:���ѡ�L���C�@Y��#��r%���7}t��U[���%�㟗��ed)�|M%���MD�BmVd��g�q5�/��7`�Ii��]и��:�T۾Ɵ4�Υ�vbɝeycأ��
�\���X��=�+	�A\��h]߀|D	�3�i=���Q��Qďf�4�*���C���J�v�s?��GS���Ƙ;r(qS�h�!��c\Q�B͗"��)*����<i떬Vb�@V���f�b��K/u��Esj� �
�5H���E���}��N)G{��*9H��$��眙7�!z�+t�!���>R��rKj "=D�O�
����q� 5!t�]�\^3:�7oR]�B���	~;`��;����LP�8�'��ґUeR.�O�P�$�:`��^A)+��Γi�* �dY�~��c��n�3Q���$H%|pS��% �������3y��F��E� )�������9ّ�	LoR=�|%�z���jR��僧�����)=��:�0�|2���/�'/%Kon�r���\�o�=�]���b����W��:C�ͭ�)y�#d�M	����}Cr#���l�����?J�J2Q)��)�-D�/��T�;듈��"T�Q�~z�㦴��z>��>��tTz���A����HHjd^E�j��$�1r���EY����7d�yO� �����eh	��*��Z��8�-���r�R�L�ns�F�<�R��CX`B
k�	�4�Y����"����&|`F�+3��ۜ��cD����Q�]�"�&���P	��
�x���і���_ї�#PyCu�u�Va�岚�������'H���v�<s�L��(���qe��^dZ���ۚӆ9�yƼYi~�� Is�R�4�qd�"�r�$
��	H���J`vf)UY���	�3U���� y�qt�yA^�N�8���e�< C"]P����)��'*���p�|�m�۵D��A4�f����&3�����@������C�+	,� �8��M�7V �^Ǣ�g�m
�aQ^��eav�a�0'����}]:��Hl����j?� �h�`(�"��`�[��̏I���B�W�Z^����т�2ʳ���Ti�=����x��%��M���F��[JE�������˸&��Q�^]W������ONn���7G|��ǆSjI�c��V
�B��;�:��%jnI����	/�8�*��_&��_mƫ��5�<��р�òa��ӊY[F��k�]#���49�/���؃`Tf߫�\(��z�;*�7���#����P��n��a
��;�sD�����<'��{0�q��rG��{� $�ӽ#H��X�;�/v�@~+9-��ZPW�(9��O�jF�
1��8�7EY�-KB�~SZ��eQ���BԶ��K4���3�j�G50�����u�k�U�ّ��w��/�U��ZZ3"��K�O��}\�u��o^���T���#�هE�ȓ���dayl@� Y��s(��Et6Q�hv{DaƲr�B;�*�q���.*�鞩@��f��%4�΅����Z�}gn�.�uKF1h��h��O���,���}�?��,�{��R�%v�*�ls���	A��m�&jj7�w�s3��a\�$��EQ"U����i5��E@���(����,X,���I�+�(z`������4:���Q@X����i�u�؞�,�6zW�cQ#��C��"6?����#9
J@�M�Y{��m6�B;�yh*�DN&������wZr4��ɦ'��������$�d�dz �_���'ۭ	j�]�ߑ�o_�σ�a]x�W�݋A��{8�p'rY�Y�TΎ1'���J:_�-�KI�$�Xf�3��K
z��X-�ûXb��A�o#p3�s�xk�:NѮ�r�i"V� �%����4�Ky��P�5��P�[\e�1�k{��F��%����<���u5 e����W䔚7����-&��!E�&
�K��D��Z��]����i5|��g�F�	���@<�ȯ����I���n�XNy�,{�c>�~W���^D�f3;z�L��gDb@�zXw]�����Iv�g�c?[Z�&:�ޱ 2��F��������2/��TA`�8Rܰڐ'R�M���kJ`d�f$���bX��������������5�b*#��D;�7gݿ�+$/��}�nQ '۱ؖ��:��ol�@u�������*d�-��y�	��hLB����/
^�C3SM�9�yE��
:�h5Ga�k���߄4��'h`PmD8�$�e��Դ��$d�Nd���;�L�����&�F�i����}D��c�2���"Pf���@��i�Z�Z���zS��3��K}|�����97|Vk�U�\�S�6�p���t1Ųz��x�������OS��dM� �����6c��^��dc�#�Y��x�6)����p�g�ՠcn��A�)r�Q��P,&-S0*��{���8uG}�[|�U��h���h���3-Al����4��0��>/��v�Z/,��B����<A2G�¡KS1���AJB��精/É�W �8�uIy�K���r����]0��ڡ�E?ppۖ�[�bK�)q�ğ��\sUR<f9x�����/�c-=�h倏L	`髢��*�b��u`�q^|�Ԑ���C�A��<�܅T��ǙR�h��6��)L���x��;	ߴ]X����ߡ+G�L����]�Me�;B9f7_\�l�-�"ZV�9����J���3pe�A��l��X�h�c[�NE�f����H���mŉ��Ơ3��d0��������Z��{g�pAyd���u�#g�B�Ï�����;){�y���i��L�|��ENZ��k�YS�:���"��$g*X���܅J��s;ݫ���Fg�kB~�t���Wy��%���\�V��,���	\J¨w>@�oW��Ӛ38�.�BM� Y��(�3)�%x��њ�p/�8@�)�*�>���F��p�%��dh��R+�-��֚k��f%�=�<o�j�p �:�p�L��r� �]Z?d;G��=��Ғ�$Ax�օ+�6�e>�u~��Ý�QghjCS�%��d�� ���O���/�:�"�Ϗ�֞)l����/��lcO)HG�3�^�J1����Ɯp\����tk���������ōm�͸m�<�E܁�O��4�I�l,���:4���3�2�Y<^LxK��Uqu;�h��)%�2B6IL��ҋ{�\�@��z�����*����H+vA]��E�h���B��>�(�|hs��%���W0��5�!IZ���Y��I�݋-l��L4\O�xvtЫx����P�cH�����"���(*��9���� }~�\�[���〧t�B��-J�\{˃U�D��p0�95m{U���滩Y����̘�&p�����Ղ�oqf�S�UW��W=��I\�f����'	�q��`N*�*��~�?X�7`Z�B�<4B����럴�����ۚϓj��aLH�J����r�WԽ��}^�ׯc��C}�}��a)����i��
^_W�>z�@7_�S
}W2�~[�8ޕ�o�������B-.�����$�ێ��^(���)b'��)�(���!5<�������?��<A����}v��[����3�f`��7×_����U�U�w�BNJ�+i����>cr��@�<-O�΁���DV�@�G�q U;�K�8�w�h;Zȳ��zc�UϨ��]�����ĶL3�ʟ\bm%&��Ѐ����#O�*'�H�>������r=,�~�	�΃��s�.��v���/ē4S)x����]'+��z���@�:��Q��	^Uh�ʿ�,�,o�$��@$Q��&�n+$^\NKd���1��b�%�?�r᫇��P�	)�"�GI���2�W�	5���w X\��2+a�)3��R�h�Ad��xG�8�&�0�����O_� ]0��<�.yRIm�Rg3(=�A�.�l�}�MW� �RS��m2��KYa��)�_��k�؟��~�&�AZݹ"��7�\HW�Y#K��yӬ�:
+��Y����C�% ��J���t�ӂw�KA^�do�B���v�m�o�i�X�O�`�ENkBl���"���&ql9���[]�(���R|��eC���S~r ��b��zL��׸1�)M�#;&L��&C�^w�U��� ��R�:5܌^�zX�X8:�Ķ�YniUTM��oQl_|��+�"nC�%���ߦD��35�z�Jհ�%�FP8X�aL�o��pY(�#~3et/)dVy��r`B:L�pJ)Tt�<��2��o�K�w-�;�Դ����7��+*k�Š&{ `'_-,��>ٲ�"�������E�`x��-H�V�+��sIw�ʬ�nVm��VI۶���De���eQ_���F���a8&�|�ʫۖ}]|�M0��-�k��X���-I�pu��u�K�y䜵	�~��1����/�G�A�����>������Irgݍ���+���7�M�5T�뺲���(&�b��BI�,�t����uU%/K��A�k��8'1$3Y�������P�4�w��5��2gd|��)
���Q��$	�ˉǱ�L��wF�] �i�+�phV�����L��T�[ U��<�lR�WuI2D���Rq��?�X,�^_!�,�jk��T�~XU�R32�hZM��jM��ߝ;�ePv��gf=����w��o�י�|��>��}sI�n�ī,z�i�D����� @������k���z�_�Vl�F�:	M�7�WZzZ�Dz�M��y��	��L;��-:�fؚ���:�x���+�L�{i�ʏ϶+cj��.Q��LXh���4�?r� �<&��H��[�9[
!�,tH�!��	�[�O�)�Un#��ѯ]9?������"�VG:�5��)j�4��5�M=]��
sD�����)0��gx~fj�ǩ���R
Z�^ŊuIČ����6�o�$�3�Þ�7�s���p=�&%YS�(X���l�NҺ�0A��*�2I	B� �4��Qf��1�NjL;T���tD��j�]��0@4:��Ƞ �>��P�Jw��I^ j���� >��h��Ѫa{8�#6r�O<�7��,�\���q��P��>J�ԝbK~�ղ��a�ؾ
!+�R���틈h��0���#��O3X��Ⱥ�}QA��|�'��P��4�7�+`�="?f��=/��[v���ߪ��8jLD�	?���=�R7�������n�'^�A��Df���c���
+TNL��}���J�F��e�/0;2n�w\�K]�!�Z�J��ǌR�F�h��O�����yщ��	������Ǭ���%��}���q����&$WI���dd���Y:^�z��2hp�b���f+�"��2���>*i��ܯ�N����e�= r������{�1�8�(=I+�c��^ F��j	�.kPE�pm s����J2�e��+�㱟��|J@ӄ�+�Q!."����:���s;лN��)�/��E,s����.b�{�Q�2�E��/�T��R��Qgθ�I�,,��;8������H������b�����$�hi�j��x��>�p�2�c���<�L���H�'o�e�D�S����0��c�����\N���:&}\�Z�(&n[�)�0�#�Uk<��@�Cѷ���_�$����L�Ex^X���ϝ���oVE�SQ[|�V7q����su�k��^]b��s~A��\��9��`�#� uST��Q��9]|�gm1�	G�\(wwJEdx��l,n��YoX�7R�{�5��#��[A�)��Xְ�lZ��~�b�r:��;�"8�%
� }�8m�&��"�P�4��?�W�}���� �O �%U�Q�%)m^L����ls.�M����i�P�E!$�[n�E} �"ÄYB���������	��9L�#!�&cR R��*�����l�`��J�.��஘�6��Q�;��s��y�w��}|��0�8�*xc>v\�XL��&=ԆL
G�l�d]��7˯�N�<XA�NH	�m=|A�8hgJ-%s-#l�1U�Q�qz �i�O�D5�K¼�\8G���5\#�hN��,|-��x�:8�>��UIC��1���iB��|Y�X}���~) ��1��?�ϗnzG���"b(�/k��σ2Z	�oC[��5��˩����u���%�D��6�7��:@e=��K3p�,L��\����jG�����Y��Dq;��� m��Y���.Š��E��V��}�߭��k�7d���q�b�aՇ�@k����>�ɡ~�񃼵ۿj$\rR{9$�����	����ٕ�Ӝt]�~��"��pI^4I��I�GK4�q�q;��a:}Lk�lǛ�F�~pyw�1�
iי��!���R�+��t;ќba�����m�Sz3�B��4��}c'm���>��	�����q��Hz�z�*�=��K������P*�ܨ2V�R�a����מ\���p������u��5jm�ЃDEF/,�~����蝻��$Y�����b�O��
� Ĕ|�$>����wn��G�lx�%�i;n}A�R�T��M�M��>ۇ���ՓY=Z�����5����Uy���:�UY5!B^��ҋ<���W8�N��8,���,u��6�!AƠN�C23� N��}�L�RU�%�0��Y֓��4��7����̵Ov����ҳˍ�z@1,��J���W���FF	�h�-Dx�ۏpv��;6m�B���z��k�mIb>=���/k�YJ���Џ\/;&ξ��(@����i�N�1��]���:�4�5y ِ�l��!3>�Q���\�F�8�#r>&dS��bmS}3n�P�T;��f������Q�\�5٩�3�k��3��W*���"GKƳ�65l�޴�GF�K_�G�q���h����);���ݯp�u�Jg(�'_y�����M`#���`܂��������>ܑ֌��5��*	���X��y]��ިRH$A���@��q�d	��"��C��f+�$�F���Ç#��H������~��0�J�T
cn�F�K3��P	����X�^m��+XLe�3-r[�������G|7���hP�� e������<��c��)��C��Z��*���;�������ϴz"��Uɇ����7�{oI9�i��ŭ�d`��_�Sc΁��H�H�rCA�:��͈G�&�V�V�x鑖�/Z�D�ֱ��W8�.�|�l��4�$l��5���So��D��6'>n�؜�6�m",�512�g�Z\X��l��lZ�:���1�l�-N��Zխ�:��Y��O&ʉ�ů(��(���]7M®Y�����A��n�����	�x6��	�����֎��gU��u�#���\�q*��Y�D���|0��`��l��Ѯ��$$�%��W�O�k�8�z,0o}��:7��iY�R{��e|Li�tyR-xDg��<�]��7<��i����s����-�������B��lF�|��.=t�IC�ٿR)�t���^v����0���49���HEd��&c\"��G��i���q(�@�SL1G��m����mC���71�/N�hE�[Y��T-	]�i4�{>7��.i2O����Fv�i�3Ls��/�\�PFE���¼�+��y��K�k_>�E�z�\)���.��{xP6�G��v�V�A���7�� >0�����^`���ԥ��;h����"&��(�����m\��ً�u{���)�gp�밁���CTU&O��j��B2q>��RZ��#�s�x'F^���O��Z���,�X�ж�as: f($sa��@8�C��.}�jֲg�A�c�WT���o�Pgs��̲�ԣ�h*�-�cv�j(�㳅'lL��%ps\[�Q�˧��2��7����PO`��?�D�L�4�K����+�j��}�9$bT��G��qk�:C�C��Q�,�;M�<�Y��iԏ������-ňw���k��@�UY����&��#J1�H���rt_ iR��՞��8c����dsy�˥rҭ�������~��!��p<�Y ��`�;^HL�m�u4bl%&4M�7�*������Z����h��h)��1���3Sg���^�����h���Ě'��MF�����݉J3� Mwvˏ�U\8��\k���4;'�T��s����q$K��F�}Y޵W��<WZ-y3��J���8]{�2#h8����O���GLY�"��Ԥ9��_̸gS^'��9-C�M9�q>�[_i�0Wl�XW�F-0���/���
Q`��;�{\e좦᳃g�y%T�v�����M4�=\�;�*��K���W�G��hT���r%�;\�Q&+��xs��FY��垖%9ޠg��МO]k���Q)ZV�[�/�����h���˨هW�A�*�9F��7^A�J1��V�1����l���������4<�/�427�@.q��2��B�0�`�S��:��$,��%�ë����ko�KԄ�W��fE�c��hD��<:�̨4D��/sb�1����C/��c�1\�k�d�^˥���n�(��b)�8������jd���ޏc5� n\ٷ��6B�O%����*���ɤ��$�:��"���[���KZ�"�Pv�x��Ȟ�i��Or
yT���Ԩr�F�8l���#�V۽�C�#A�-ͷHt���j#R�C�]���DL7x���f%j�/�P������>8iJ�W�V7o����=,c����ߔ�e�EJ���  }�o������ g\[v���J��Z<xY����oY�%�>���]{&�[��mF����p���&���jOH)ؒ|K҄�DSz��nJ��w�{f0�޳cc�⼏�yi�R�'d1K�\#���=�/ ��)yʟ=��~�w�0�u�5n�a��-K��m���^��[u�=��0B$����H�.q\�������m~R�����&�<Fd�rrբ�2��V�&/���k�Zs��w��>�,��t�(U��Hh(+rM���'*������z���O�=K9�Aܙ��QiN:��;M��}zL3wg�hD	�'�G��I�*)����f��[���U�O��
&��c?9�RVQ���W��0WV��>WW7���:�mf��Iz%���z�	�|��0��a�67��[��3�]]�5PG�J
��~/R9�E<X�\+G2z�m���?5;��I�i���S� 8[;n��.;�խ6�T������O���&�m�k��Upny&��u�Y��rDhM) V�V>R=B�s�+�k
�_��etXܳ��� ��x������r���2n|_͏�1ؓ����(%<����:���#��qk�i�-�3�d]���~���R�n��H�Ҋw{-5�=���rsg�u�i�g~����M�$�XS�v�gh��� ���̜��ܓ�{�=�� �YG}��q(ߋ�Fi���&��=�����?��.PZT�W��iX}�p��\����WB[o�J 	��ợ@�ټh~���Qۯ����]�91ʇPc�*e��H9�xG�S�8!���HU�,U�n׏��Iw��	K���Mg��;I��"C�}��Ri��ktS��u7A`����� 1�]q�PA�y���E�hL
iŔ������χ�.����O�[�hu��0���M��>	�ԕ�k`�S����V	6q�K.��u���^��J{Hx��������n���O�PM��QC@�K� �����2�]���)�U%v��i�s(	7��`l�(G#��nu���7��M�&�k�lg����+K��ΑQQ��Y�I}$ �1��=C�b{�,���������m����3"�����v�H����w�Bǭ�LS��NiF>��ke���I���b���si�o苿���% ����we� �]� >X�|w��P����G��\`�� �"���Z�,a�)��9��n������@}���W�!G8
QJon�&���CyZ�Mi��,Ku�A���B��A�j����������'�qfp!������[���\c.]�H����om�YAU7C�']~���.E-}w83���xl�3p@@�����u�`�ƙ���Ls�l��Ҩ�Z�����f�L7��C����'�Q��O���
�ҋ�W�����`E`�"=%�M�3x�~�*\���]�U��r^��D��Mư�g��� tO�L:�2��4Hl�Q�A�;���@pqb�h-t �+���GU���Ba�r8�n�`%�ܙJ��:�T�ϡ#9�R�\c{4�_�!�P(�u�F�EY��mo�B0d�X��O��
��>Va)d�o\#:����$�C������5�����D�ST���ݷ�C܄��P �r[\�զa�҇k��D�:� � Du���x@�R9*�S�n�e3��QGq�L4��h�h-}�)R�d82���gy/��;!�XF	�fA����:�T	S� � ��?i���cB����г>���~���$�a� �3v����~�X�g~m�5�l���/ �D"Y��L�� >�BY� �J�N�u:hn��	�,��|���r�{����i��Ң\��A�����5��7C��F2�m���Xߦ���䙅}|h���zP0ʫ�!
�|Vk�[ +y�DN�'G�`�Y<D?�f�(���=�FV>���Љ~�^ ���3yY^���<�ͥ�I@��8��MC����]�J4��]Iړ�O�m
im|ۋ�������i�v&r�a�䀀pNC<X�|�BW}��JR���=�e�lWs�2���wrm�
���ᕈ,<nT�\�E'��e�X���s�!V���T��ҭ�Y2 �5e���.��ܼW�{Ƹ�1U�S�L$f�*<��誛�ME,I�N����������U�
�Q=���q*D�����Qͬj}yC�! HaCЅ }<:��9؞.ȣ����K�t/_[���C���@��~��9���G�c���tOv ���&l8�� �&��Q��	�_!(R��,
���?pO���� 4Z���K��`��S9���0f�Ij�l^~D�at�9ɛ=>�������s�6Q�d��T�"PD���|�Vl3����>@_���^�`����=�n�<�ƿZ���F�a�Bx��� !`
�B+�(b�&��ϰ�+wp}b�����z�;n=���?���u�S��UO}���%e���sw���	��&ۋ� �nG��$�j�z��c�"��6�AN�B�H���������l�E$�6S��g4	��d���.F$����A��G����9�ؚu ��5�*rba����J�	��1 sT����5h�hP-5|9�	��b3�X״���	G}%���0��&��Q�2v�Gy4�F:TN,�L��"'���w���(��G,�PBf�kT{�@/�����d��G�2�S���O:�ײ9�.:�"l�.��g�&8xd*u���]��GZ��1�u���ױ�-Q}�# T�>�lអ��X��Ԯ���+ʠ�cvq��xͶ6+4�ZoMZV0�eYp���0+����)H�җ�*��e)ߖ����ɨF�r�St���6jl�T��d��`�0��0p��n�o-
���s�� D�/5���ג���j����i$)Vqk*��C�@�)�)�i�J �7�Q}��5�]��f��ز|���(�z5�TD�ޠqw��,�H��og��� |��j�҇3�Pv百��ns.��R�Ϣ���]�,���Nj�׳"��*$�0�Ԥ�	%8��)Ϩ$W6���B*{�~�3򜌵�6���tIC�R]!m1�qr�P.W��lI�������G�9��C����d�`S�2LTk��F`�W@ʧ�[�P�|M��\�pKj [p�����-$���z�0f��w�-�T��A����I=��`����1&����[��J���;d�����|��o�+�q���N��
���4Y�[;t�¦!O��s%$��
(��� }X������g��@~��s�JW�6�Nց���L�[a�,�"Mk�	�4��k)Ek�432c�֊�.���3��b��o)jM�d�Y\V��.Y)'�S���ԧ�JS6�'j{���K��-|���es�o5"��k��B�Q�7Y�X���|K��F���(�f�AP#��ͪGf���y�6����+f-�ǈ�V�&�9)N7zz�!���}?�A;�O0�v���IM���9+�	nw�L�}�ʬ`�(?r�&ǻ�4��[Ηtt���R��Z��LɽMZ���b�6�A��J8-%S>��.��b�@t��K�x�ԃ	���"0f�u�,z=�5:=��l�#X��#����[�	��℟ʻ|�R#7�)��3e����h�(gzا� $E��	O`*��x��}��Dg������+���}2�n��S�������o{Y��P8~˱��3SQ���5R���W��٥�h&B�K�ny;@Q�"�Mؽ�)u�fS�砤�c�3e��4��u��c|����y&�p�O8	Ò2��U"�Y����3^��5q�ͽ��Ќ+���w���E��UW)ٰR��ڭv����q�f�l�S!e.���Ո���p&��l�/A[��Y[_�wƭ�F9�c?Y��T�+;�K�C~�b4��+7>����~A- A�� �����*��o�bB0��wK����q�2im֮4���>.\����1D�v6O��AMu�s�<P�F��xΉHȌ�Z3#�$�����z+(]Ȯ	�n��u�63�n	!������r6�� d�7����ْ�SSa�?�`�'�5��!/bE��>�w��QTp���t ���N�� ��2/����ظȸ��o�e)+��F�KOI��+��E�%m4�Π��L��]�9O�+����Y��Ř���=�����"���ōR	|�:R��`D�Q��v u���\�Е�}y�8Z.U�,���N�B��c�hN��#L�9�H�<|�݋���Zu-�(Ӑ�_g�Et�z�Ţp�S� `��o�JI{H���BG�J���w1�Dh��U��wx�1���|��M������,�_�N�X�eYW+�у%�{�d��-s����I/��xy�`l]�b?^Uv��2E��I�݀B{W��>����s�ǰ���U!|��@گ��{��_�4�1�Aw���u5o_ }�C��1�b�q T��
]��bEW8SM��5hO��YL��)����t�U�ahs�8S(���6�66��.��vz��3��s��jξm��W8ឺl_q�Y��4��^!Q,8k���_-�괐S��gK�Dſ'p�i��̋�[LOu���:�}:��~�n��9ˣ�
M���ɢG,T�c_A��ܡR�Bb!�`&�<!�0�٫@.�!�G@�\�����T�>s�����l�q'�������O�F�.ߝ�2�����C���ʢw� �T�&����j����*�1"4U�����%j�$o�U����N������ԓ�*�U#�*&*+�SC�lDlw��G�V�
1Q����W�Iܼ�\E4w�ˈ �Wޢ7t�𾧨R������~�Bb{�bn�Ѩ�U��2
�V���uv�/�B�w�����([�D��e1�;�X�
��&^���^�H=��[g�v�&���^L"�ݶ��	��^]{G
�෩<Y��Ԭ�2�+F�p��>��Y�wr�fb�~��m���:}��4�QF L�C`b���yF��D��f</����k��^�2�q��F�QDMF�gf�w��{����CSa�زyi���C���WM��.���r@�O+��k���	�
N����C�Ђ\�<?�ǳ]���՟u+���,%�^Hْ��Z�I�΢>���Y��@�͝�6*��>Ψt�B��{��6܄�h�4�4�
N�Ty���ڡ�ى��d�\����C02C7���u�!�pE�=���y8��-��u�#�j;
�b�O�7Fo<+�]-�`�y*NC��3@u���#ָ��Efk���~����A��X�=*��<�P8����`��ܯ%x�Xv��d�Tc�'c��!�k��LQ�%�A�HeBSPq�ݕ�O}�ǎ:=Q, ���{~�$�P�Df���ȏd��jI��B�ˠ,�M�G��٨b%*.o��#3�Ѻ�g.�tr��r�<B(���
o�z�}�I�߁}bv6�G�Cٗ@�����؝�k�H�9�M����*f뙝�K�)��Q�_J�1���{�uY� �	��sc6�2�Q1E����Ȍ>>�v0# ��� �
X�	�$�s �kL8I����|G./D�K��	�C9N�~Zr��*���i�#�ƒ�|+�I	W�9�ya$�w�������q�@�W��DJP�ڌpv�9~�dy2H��GA6fǧa���dy �φ@Sab362�<9�\;���8�e����Z���D8FP��3��+�O-6C8���u�]}�@��e�N��Þl������P���,�ny��A��ɮ��C�@�u= ���йC[袹\�jP�ح#3�'y�"��bV	UAL��֥)%i/M�,KK멃U�ݓ�2(���ݸ�ũ2QU�l���R�3x�����A(���~v�?~�hkv�mxik�K+�c�dP�g0���+r.�\8y(=f����z�
�gH�8�L|�1���VK��c-�w'�}����7�;4�y��!	�a<L�(\���k�P�Z�HN����ѹ�#Y~�K�Ӓ8��#�En�s�z>�[���k�*���z�z+N���y'���kOu
S�2����o}�,ak����)��&��{����V�u�� �>Q��{�Aq;L���V7~+F�j!���`8n��a/l�-�l� ��A��m\�v0�a=®��L�pei@ ��M���ZQHV#̝t#�����L��~��n<�����w�芹A����H�I"�Q��%|�/e}�I���[̠���F���ԅ�������m��s����`�� �ğoa�ͧ��TR�97�D1^��Ȁ� �����ΥV�s��!������곝��*�h��qN�#�d�5(3�\Z9����[�t��e��N�aAt23�н�N�L�,#���������ʏ�yG	ĞN�z�p�d�]��sg�b^��9�j��=��ɱ�~���T/W��
)p��Y�iۛm�C�*�V&oR����w��� ��:$�NV?2�*�5��A9��~H�)n���;�F�HBV���t�[B֎*�����XةJO�~Q��Frao�5I԰�wU�ƨ"�,�p�+��0��p!J�%M#�T�<����V[[�biFJݎ�ܘ��s��֏>Pk�<#��^ ��R\@w��2�jjn��w�}Ɔ�V��# ����BH�����Z����e}�7�yOw�J�;x@6�Kq,����pkE`�o_��s�0�u� 	�;��igH���.m�ɧ5��Qi��S4�`W�s�uK~����:�}@�����:��T�E�G��r��ǀN�V���o�$�B`��5��.2;�!Di0��)��(b�3hP���O,
2;	��&iK;p�?��Z����"��śg�(����6Ƽ�]>L���ķ�揂������ke����&��ҮFhڠ#�3�IlyGcb��~��P�2�ϊ등I)�x�31�+����(=0\{�jS���hk��v�p��eyُ~#L� N5��N�'�U5;C9�g@�&�j���V�	ch�w?1�g�F ��b��!���<�g������U=<���f�-��%�%���l�2�cHO�l 1�B��3v/fA��&�ufaY˧ʁ�0�i�\!���5F��w �6���	���ou�p��Ϳ���I}�� P��O<=h��'���@yLڬΡ�	voaB�x��1t`j��~����am��Mso%�@<�_�O�r�dpJ�rO��_��4K;>/*�@H����x�RI�P�I�Kǈj_ӻߜ�n�����*�Օx'���,�J~B�v�m. )3�ꡆ����}'����7�w�k��������ʨa�6J~e�v4�?��XfYǨ��ߍ�ȟ<E
���0�x��5Fb�9Y4M�o?�VU���4�l&��#i�*;ֵZ���Z��A��r����O��W������&L7,���~���o�����M�W&jɁ�ڏ��-��4�����3�j�+u�.�♨3�)�V�6L�L�1c7��c�����h�9����/\��K���������C�]�݌ǾL
EQBw��m�EW����3���8����tȠI>�a�Ӥ.�����R��H��t	8|'A �)���OW(�&i�l|�RX�R�h��lF�%>�� M}V-y�۽��7�~����Nx�	#@"q�t$�}`]��n7��Z�w��9����L�f\T,��B|06���S�s$�\��9V`w�K�Qǿ�p;� ks ��ýR�&��fI�p~7�)����;�X}�SU�"��m5X��dk�x�	���K�Ito&�����'�Gʺ�a�v2��W5��=s����\������������ʋ�{埏tb�	�nQ�I�k�z��vן���E>�Ui
Ap\���$��y�����%<GO���۾u���L:%oo�����p�׶�M�@�暬1c���>�6�t/�'#��_�^֛����&��N��;�؄�b��h���?]n07��D��ඣ�.��&>��;6ls��EK<��̾f��[:�SW5o��F(F��'����A�	����F� qZ�r��ɂڂ!��>Ԓ��i׾e���f���EY�p�^w)m�K���bUݷ|s�ńsew�^�ǪG�ɛ�����4�J27��� 9�o2���{Í��f�_�rO()�Ŗ]��XW���ۜ����e��y<))/�=_���d`L����C�p��Ҩ�;�ZH�_\��7^��t�%K7 �u�-rqˁ2����lBe�Ab�nr.��/��G�f=p�xNK�Q?hG'�����6��ަe�2���b�-����b�t���VL�8�y��{G2�n���>߹��S�Q����7 آ���ݮ�8�l��`?Xy�euۙe;�C/��U�d� �qzA�|�Z��l�m�/4��&�{��4��_c+�괈��ʒ�3껀v�
Xe�a���a�oSF@��5leh?H)6*|g�@�3��1��P�	��r�|�@��;���b���'J�[�>{�WB$��Q�g�7n{�q{ �</خ)���@�zm���+h ���,x`�q˜JSrAPÓ�@����泿݀V!�� ��l�_��K����V7�Y�H�(q����\�Dr �;�i٦h�P�L!���!Ì�T��邵�o�7�8s�;(	N���u��"l"�5N�@�8�"��[|쩗�S	՛ש�\?\ʤ������-�i�p�w�E��րU$3v��e����^\�}Q��p�S��n�;Q�I���S��d���[�v����������"���ԡ����H�oY`S^H�����l!��[��H1%0�y��7�r���**]�G�Ӌ���~:�L�w���}��avx3ph�$��ʁ��l�֢�}%� ����ś���%V�����	��Λɫg�fOj{6��ʴl��:~M+� �uC�?�{��  �O3�m*��1'b)U��g�d;*w�c]����[��0�4����`ҡ$�0��sU(�V����ѷY�c�xڂ���Y�� �G��� ��-W��qb� R��zP+�ᨧ�l�;ي�!��y�ChO�ӯK+�;T�%/-�_�gj������rg��`��3go,gDx��yc��N����Vd*X���O#�:�0.������A��^�F[@u9��/s�6�,���Qx��$!�[�^�J9n?���㧠hp*�u�xi���:43cZ5& sF����2j5l5u�#u���bܡz�v�8�]��#L��	y 5��gs���-�=K�Ee�