��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ`�2�N���³)������t�^����`���H��۸'�U!|F�lu�#�4�v�Gd��R1S	j0)�)ۉ�v?I��0�M!�7(�@�٘��"�j<��#��qG��#�0򨈀�\��m�AJ4������9����å>�j�ͧ�}���^�M`z]�,����}�u�ep��{��o�?�A���-]��H ojke%냍��`N{1[� �z@}�'MA\�:����Ⴔ-�E,�0�3����z"e�mgc��>|_u�0&;6����:d.�-�T�~DҀ(W�\,�E?������jE��V�Kn&7�TT��V��}a��8��^��|F)��]Tf���G���m���&��#Yf5��]ayj�~���y�G���zlK�]�8��UE�����]�i%��e�/Q�M)� +KR�,ϥ���I-�w+�uZ&(���F�*� �GPsb_Z�Y�|0ֹ��ç6��<���}x�N��C�Ol�/y%��R�;^�b�`Aު�0�s�i9��}=�c싯	�ǒ':���M�4�(�^�k�����,��Q�{CA��J�
�u�����]h��UB�5e�EMDz��.��yr����|7S����=��6��$�%n���ϴR\�_B�(p�_�� N�X�JM�-��������4��mA��#���-���x��2�~pdcY*�*Ԙ�^*��|����:hP�g��Z4�{B�c�5:.U���tL�t[�Zx(wCN������a;�$-�G�ZP �R}�x��_��&��Tw	�D�:�Q�ʒG|x�6���8[�sC\��Ż�*$���"-��4�P�4U����X]T�k9>�� ]�']/����)�g3���[���0}�@p�4#��#�1�w^�l�h��u2+_K��"�/\1�'^�s��{W��>��V�K�Y@:{��w�^|��~��J��;�0%ë���H�����z�R�u�Z���Ɛ7�� d�^�DS��Sn'n�\;�o�'m��~<j"b���(��lr����8�$1Ġq�����D�8��]p����ʂ���`�����.bWJ�:?���<n������t�`�C�aI���}���Z�i�I���Zۙו&d��e�x���Ns���l
�$�'O3��~�6��ǂ8�L��u%��F�޿��7
訮/$!:����Ss���5+��b&]���4@�[v��īH�FĂ��!��θh�'��0�C&p��aa��3>r�:xH� �;9��߬gǑ�xUq}Y�Sav��A��m��a�2΃1���k}���WwZP~�Sҋ��w�� �5�v�����H��/��%�3'��P��[@^���^g&����ej���d���!j(�`ڲ"ɛ�"ץ�:3p�x��D���3v����w��<�9`�"�
΄�$�*|Blwr�P^#��