��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ��Ul��?������,��m�M��t�E7\ ��7z��-6�#��<`UJj�I\9#��zW�x^�k	L�c���������1^T�%O�b�5̓�#s���x�R�c!"���aŢ��#�{��vw��7������U���s��bۍ�iG�l+V3�եՎՌ���o��Dr��s$վ?��F�|)�i�*+c
+Eb�
i�`j�O{F���{�䷛��w���tx�L��腣�Q=%}�!��;��n���Y�`�;��rE�`��^;��,�����t��W�)��|�����N$'[�xiA��	]���$�6�e�����p��ʁן���#���0H~�8<7bE-pk����;q8h#�U�;:}V��T|��j��B�,�\����%�湎�p$�61�>K��z��� (=�����'}�C\��0�r�d�?NcR]�G&��Ih�j����΃s�$���ZW�/�}���u&f��#FR��<H��g	]��*λP0���0�@A���e8w/�_ls�S��n1"�Z���eWVC?>��p�
����_r��S��ip��9�����u�w�G��!T��/��X��W-ؔ��]G��-��I}�9�f��]�C��~�4�j�q %���1c��T�%��G�ĆV�l"�q� ����&���{����&C�z��`r��~J�,����ƃ���>��Fff�h���e֎-��'�p���H<h��"�������I���v� Pԇ���@F�79QY��7�kz �?VSQQ}����4�V������;�#��}�����k-Z���㷜��f��\���fu�L���-������$`���ʔ���/Cy}`_�����SA��@��pj���"ۦl-��?Ń���cv���C�������:�Z��O�:V���&Y��h׷�ǃ� Ly�%˺���x�!����ʷ�����E�2m!�@��2��M9ql������j�X��H��S����ϧ-DvOx�;0��J2<���i9*J��l+_>+q1P��z�6��@ϥ��5͘+�"��%79CC�2��E����U⹣]��|;$lk��p�<�щ�|�������g�}�0W^ش�T<�xMP�HrŮ�A[�P �9�`Bw_ε8��Q�HF�h�Pnߕ�H)F��E��l��u܈��.TPx6W� P�0/����R��<��3c���_��`J�]沐Z#��}��$�f�Sn~����g�S�P��(�T����(�P�����`	S�!AR6��c��}���Z�t�ku�H�Ķ��k�p3ڭ��)Z-�?O���2k������ed���PTSW�x���!�qi\ۋ�2�Z'�ߢ���9�~�E"�R�D�I��}s��6�v����AaC�c�G���ރ1��6��]#�۲��<�.%r����W�r-����"�Ś�{������Lɛ�[h�� �w�\,�������4S�fگ__28΂c�L5��P�ݷ�㟴�4�W�C�:>�������C|N8>k�=��'�����v��v�)4�,�{b�/��8c�7�E<@�����I�e��R�q"���*������JځE��X�+bGDݍ7F�9tg�E<.~�[H�d���ā٨Ъ�r��($�m��M�@�A/Q)�g>�^t����`�wvR�?	�F� 
/���4k܂��4�������˿J��\�T4?�$P⊍I�g+o�f��@�:�Dl6�$���.l�+z� n߻^��@�+�S��gcn2P�q��Ƈ�+�oQ�0j�de���a�R�O���$�h���	�H�B*@��X���8R�a7 
�iup.�eN��\�Gc��������W�}+�:�W#FN�7\-�r�y�v݊cG*��j_{�#�\8�\	Dxb�:�g�CI��5�]/�9RG�|X�PfƇ�2b��H"�6��N�p�|����&T�xd�g��٥E.1�,.)
�ܙ����������h��V���=a��#���b@[*V���2@���E���Q�q�&(m������I��T���62��}�I��bӽ��+}v���d<���m?1��&�|�@�<*�o������;����%zE�Or�Nc��hI��a/[���x��㚝�u����������J�rT$�Հ�� r����B�Y�n�b=�]<�,7��-1�ƿ�S��K�v��9`7��&CM��u3kΞO�D��0�����r�3���z>�s���YR���E�sάy��Z�� o�H�k]�曑��)��М ��p��n�T|�C��b�F�9�gTI�E㱬���q��Gܘ[���GdX	q���C�߄'��DM�2��ӻ��LҤ3g~[ю��Js�C[�����;"�D�"��r�N�
���Us('� K��5�@�����J��SB����'�ܖ�����,<5K��0�:@�p�
9��h���.�Hˑ�r�3�[����샇{������ҮRF�n���q鈎��n)��6�J1��J��t���F(�|��W;�4�by3�WWX��*�P���I���i�L�V����u	���R&�1���ӦW���
�%��.�%/8`���W]h&���^ڿ�Y	8D��!��~Ԓ��䲏�v�yl��2��Jl�Ad[tUu���xW�g���G�	�鷰��n�I�?���9�J��L�q��;����N�vCP�]� yY�77�Њ~w�5�g8����Ď]C�Tݓ���Vt�Yk{��	n�qFbm
�nF�dr����3
>U@�(�Z���޷b�����
/�o;6��$��i�=d���� ����q�2:�+���|
K�$ڱ�:�������C﨤�ZO�U���Κd��'W!+pִ��>$��p�,ei<#B�~3H�#��jf��m��o��"��^��A�&/Z��m��k�e�~μ���#Dpc�r�ך�4<1D�d;���*�I�Nv[�L��P��L�k��!����c6_�7�JN_!�XT�@d'a�/\g���$�<f��
���{_��J�b+�g����.���B����h�����%^���,�kq,��PnGwo����p֟pe*��+�_�s�B�|ΒR=�u�]��k�},��s|�}�*Qm0xL�5[�
�`1���{�̠؈ӕ	�.�oU���;Bt=��P����������ze��̯����ڴJӖ+�N ��~d_��_��!�k�������d��.̀��K?}�Z��5+f�φ��.�~���C����z��*�n��CBF.E�!AS�#��`5��"��A;Ƨ��Ӷ\g&�S���F����#U���VQwp#�����֯>wE�	��s'�nz!,��<�Ĵ���#���V���m��IW5H>�����2t�3���>��3�JŴϑ�&n�g�{h��`O��?�58�'!k�?��p�j]/pg�>�(.���`S��%����F�*�͑w����O�5�B*B>���������7V�A��ϫw�dAK8/�w�m��1�m�:!`���E�9��|�l�G����ωXl>��(�ݐ�S�f�z�P�@��rb�����p�fv̥�ࢮEn��L��{i���l�0��7��.�%��<����E����>��7@^B5�F�-j䴍�I���930
J�>y{� _~'��
A">�KǞ��>��F���>��U�������4��4��+�f=���ы:�ABj+ {�db	�����}��;�ɿ/T|QvO�
~K�d�[�u�N�K�Ծ��yp�x���DI�ݠ7���Җ�>��p/��R�|mr��I��*D�.�]�~��Yѷ
{;��CIa��As7O� �a�ς�.��z�s����ʞ8O
/O�ira��θ���=�{������PB@��H�U��=�����@�˛��WWPm= ���������	�r��s����8���mf��
��U�o#�Q��Cۺ�Ws��B3q�X}��~�Չ��z�89��Q�:q��f�]3{�2m�7�6Ip������3Τ50�(���}��wf��B����u5�Lj���6�S�������4���x�STJ�/�@(A/P�%�3"@Sc�ޥ�2�;)E���
M�Hx�BT�\_� S�P0��\f���I�C��?KOy�����&4a�G}��$�Ǔ��[g���Q���x�{����Y^�s���
gn�����0��p���#�F{3
$��f�&V��h|UW�Z��g�6)���=��o�J]B'�e�ks!Em�����<�M�ˠ瞩q4�7|�ڱ��6�A4�0��\+^�������5Xj�֗�0ђ5�&e"b�o"��>Mjw2�TE�T�+WG��`-8.K47����Α*����*4����/ZL����c���l�Խ���������ɭC�ѐ\���.U�+AcT�v�����}W�ݏ%"Qqv���Vv"@���3���8G\�����Da�W�i
F�⪟�q;�Ƚۇ��(1?��i֭H���xN�V�:����/U\^:u��
2����G�p�b d*p��i:�.�bB\N�Y^C���񳘣�O!L>B��;r-u�L_O��^�[���({\�
:�q+��e��%Nq�AS@J�-�Ѐ�z`4���3����t�S���Z�y�D�|9��kF<��4�-�!'� �Z(�!|�(�ȍ�!'�`�ٵwG�ѧ�K5��`K����#����;Ml�i��v<�P�����Oč�|(y�Q�&\�I�op�������U����: �m�����;��Ah�J�%���Y�����,�ZE��Ni�Ӹ@��G���"s�5)�h��1.�Ϥ�T�p��8�]$Fo(�\��ͻIvd�8GV.�},R��RT�[C
�k��P1܊�S$ƌ�Ϋ�+��.6t�x�]��Q��G]}��)hO�yC��q���#R3du�f�?��.J���(E���Ƣ�j���R۰>�Z=)�HT?wӾ)��v6<�w����x(vf�J�8�'ۍ�4Ĭ�.�&N�v���*� �4��#|�:�}�>D�^���b0�΀s������x��[X&:fDb�UӔ�5G�)�%�xrv�VJԦ 	˸-�OF~����)ȷFM.r��#�{b����䆞ܓ�pjQ�V��ҿ��<�"�k���ź�8Pi����iojWl��<�K/���b/冊�>��m�l���(fi:��f�c��9�X���\�):<X˛������$4ՑUxK�o�aT��Cu��A��=w�����9r�D�2��Qφ��{k{���xVf�˴6<H�3�]�m%�N��r� b7\��s{�:O%�:��Q]y����Av���f���RR�D� E5OH�sH=ȉ��n
�����Ho�Q�b9�W}��G��	p�[e�+̓Vg	˾���=�F�ruo��x��A3:��_[����-o�@�O��ޔc���s1A�"kwz
h�
w�~}�E��x��h�+R�寕���J�#W���'�woS5pG�=ѹ�F�8�S6\�D:����#�D�P���-�Ejv}F���SUՠGE���h�W�����=��a�&�)���S�'�F�&��ְLT�K8���ay����ԇL>�ݥ�k�q&��n?aP��r���bc�|Mn�v���7�PN>�Y�|�z���@�{tyy��D���܂%aӸ�=��k�m+��_��z�D,y����%�����l�����1Y��4�ƱV$��e�f���͕2� VH.�p@���4,È�Fz1O��9/Y I|��o\���2c��T#��]i��5S�3!w)��j,���ο��<}Mn(%�l����������2������*�F�TCb��9�k�e���s#i�n�j+\u��v�������c�C�ä~��9a��c��Y�밌� 	�/��<��P��>����q#����U� �ו�������h7��I:x�L�΋�#J8;�t,�d����Q$�d�K�b���M���G�3��q�Ѥ�@���7�������ɦl���N�٫��?��4�9v$��\��l��^��q���Q����3cn����7-�� ��h����7=��cHU?Gr�'S�C�ύ����Hyk����*6�HX�}3��KK�W��l1�Y}��s�&6t��J��ʹ:r���Ĥ�M��w;J	H�'�X��r�kN�	��,��K�E:�(:B�I�k�-�t��)�727,Y|�vbA�d��0�P������wi*��*�Os�UiSJ����H���	�x�=��9Yĺ�`�C��턡��G�J6�R_7��״��Y�����U�2��lŎ �d��bѝ���켆B��ϛ!��˱6ޓ���Nm��<@3L#A[#��
΂^V�f�w*ý3��6+�F����q�)���W�M����q�R����Qo��5
b��Lq"��o�M�����~��8����[�IS�_f���>��fA<�j��ـ�� ��{��{h�Bw�|�C�/���P�����ԑ�,7n��b��BZ���*W�F��\Q�`�ڈ�ᇝ�tfa�^�'�,�Ⱦq�F�����G��x`ҋ�A���P��]/�dp�@aV+���1��I�^8�Cr:�
$�m�oy�X�~i����q��vg���sC�����$����W�l폔"t�1�|Ne�z��p��l5?+o��
T�r��K��:���ߘC��=&q�ar,+dF �f�ƞ��]4�I��k�����w�� ڔ�v-Y ڈ�*͂>0U�p�U�k�����6�������/3=����;��zZo���*����$�5�F:�<��嵭��{Y��;�U'Pc7��,����h1ڦ7��.����[�8�|/�Y��wf�ц��M�́�B�+��
��]C�V���ᵚ�2=i+�/iDR��t`�b�s�����U�Q�{=����?��D�ksg�a��xd6�^���d�����쫼M�f�q�@Mඔ	��j7 U9����}όl"�r�s�����pnu����D��WԻ�d�j���g7��E.0qe����܅�J�)J%��#�(F�W��!��SL��@� �~��*q�3�c�#1V�e_Z~����ljuy��k�]%SEN�I5�n��vv���� ӿ�	�3��t1�ӧF��k�Q�����b ץS��Ll��㒙��4��b�@Ա�g;�h��]�O,�;N��tS*�܂��P)~�Z��>"�)�lk�	���ɟ,���_��U�Tu+u�W���"����^�8�s�t&�c� ��i�`P�*|���\��3)�L5n�i%���h�][�N���=\A�m>���f��n���q�~�AR�i�-ott@歖@� �܀�|F��:���N��5s8�b���d��\u@�&��D�c4>��K����R��c��>�R&Rur�kZkDg�[����r?���q[�<h�+���8('��1PA��fN���Y�I�N~��0���l�a�x����c���O5���J��K�����8f�C�8��?y��;� �~|��!R���y��_�gh�O��I�r-�ƚ�� Q13i�Ojު�ݾ����*����xVԬ�-zv�)m �['�9�T��̚(��Ђ�µ�T>�	����kI�i�6\MP����v.8mD�����7���u�##}�Wl,���_"wX��|���U�Ї��
S|�T��!h�@����U^���2��m�K$�It߶Z�ӬD�s�5)�Lg)�-!]�@����h�=2}2Ps���"S����
g�{�A�ڻ�m�Ot$� ^�`�MZ�BX1s�2v�lB7\u'��i�Q�/I'H�U���3�5+���ʸ^�r	�Gg#�U��zQMh��oՉ��񛂿��}�Y��T�t#����	�(��˗��i�<BR���I[Di�v.v	��J����H��7D�����e��h����Ix��ڷw<�?#O_2�d��;������9th��P��i1qG�&#���NI�I�A�f@/"Ǆ���r���&�[Zxo8@2(���Ŝ���Ŵ5(�B�	�26��?X1)�ӆYV���g��h6�b�м��[O0N���h`\0H��'ʣ�����km泯I��ؤ�@�(����a�������ע��]?4���KߩޗHY���b�DGGU��	��ݠ~V�fG��e�YE�)Ѱ���m ����jPk������i��C_��}:29�He-eܾ�9�ă��x@#��gY��7��u>�q����F�y�A�β7�.s�T2��y����5�����0����<�^�!#�i&4�\�sS(�����q@�Ua9��_��W�4|9���q2r!���y]f\�%��o+��K�����[쫘��n��UW�
�iE&�ZI?Z��L-���O.�]u��0���m@�7 ��~G���e�~a&l?�J?���h)A˗�=��GAW�zZ��#�T�����e�}%1�4�G��Y�>I���*��.�8�hp�ջU�;�)��>�-�.Ё���L{��� h�)�� a}}��(�R�x���2g�Pஔ�-1ԜZջ�8�'~�BRc��Ӕ��Us,��z�N��0Ĵ� ��3�P�X�����Ѹ�<�3r��We�w��DV=P�~�ș����B�U�֋��YH��58����d��zݘ'g���X 	��p�1Z��Ge�����}�I�����/oz��<�&	o�@XK���<o���I bB���t�qu��(�9��s4��o�H:�y��|U��o��ZۀP��\\ 2X�������*�me�S�w�zVV>�%��K�n��G*x��Cy�J/�����wF:�r�bG/%�,���Pry�Z�t(�r���|uX.���X�]��ܲ�{�����g�Q�ʚ����ng��}x�]�}z�lGi�Xm/�`�~K-n,��i7�ԃ�֍Uv.��~����[Ŕs19L���U��Ҵ�Յ��-�T0�( �TM�j��@�k��6n�"i����g�K���]�MAx�k�W�tK.��U&+�M��]z�8r�p�Qie�(��_���]���$܀-M<=6(��
d~��s�?���������4�Mz��-um<�+�ռ^Z+wPW�N�,mvC��d-@�@&�b�'TV��C��h�Ȱ��C8A�#V,��Xp������������+%A��G�C��mW�ˎ����y�p(I�&�i_�=}�x��ևUk������Ȟ-7��͆���.V��u��)`Z
�"\�j��u��<�S���\
:�/F���m��͇~P�df���t��O��f .�쵗���r�~پ��F	�&���lA=��!����se�y%[yI�1�r"�1�S�r������+�>�nҬ��C�鵚[�����_��wv%��L�F�+;�򐺁PII��p�&��/0�!���I��D�Q��a�7]T�N�G����BX���&��[����̧�l�Q�����l�Ĺ1+{L\@�F���U�_x��< 9
�����g����=Vefx�T�Ÿ~�I{�ד�,k)ׯ�}>�َE��a�5����%px�6�S̃��g��F����ៀe?
Uc^��$֔.����R� z43�� �TC�!���F�����1L*��Cs@��F�^I&� on���,@f�_ ��	R�>
�	.�����%���G�����ʬ⽄8�^oRtYµb��B�c�y�Ñ��K�P�_��K�����9�q���O3~A�����%��A�:�&��&�'��m�9H��d���]�-�}T[&�9�Z�O�a�\�[���2+�GdG�]�N�#�/���~B��QhT9���X��_Ϸ���Z���J����vu�������<@���A~	����f~��P?츒�U��?W�R��#Q���Gy0���zo`�ʀ^I��А�"ZK;���b�[�v�
��1���k�z�;}� bh�rL���d���^E�e����2�fL��>ۿLS��I�+uuNw!nҸ�5|�_{��)^z��	���h%�F�t�$=� �_��W���.ӳva����#p�!���.}�К8�Р"�h����.�@]�8�2<N87"��������%��N��F|�o�rV���"�7�C,��O

��ǯ��B��f��M-,�?�;��S�!��`��HS��2��z������zi`T G�ص�q������J�^�z�}�\��wZz�!HPCf@��hS��#�0cj�@g��T��/oo���l�����������7���
��$��5J�!Yq
ZޢHe,���lLb;3B�/���{j�����Vك ?��k�r �r����ș�������N�������U�3�%���<c��q�C���ΆE�J��Q��SJ5.�� BɊ=���!X��RM�8�6���,D�����.0�=���.�M!��Y8�=i����T�\ѧ����'�O�pA�*���۔��e�B�_��O1���y�}~=�|D{������S�{�:�ƽ�&;F.���^{Խ����%�dIj�-��#q:
�:������c=ILɑ�9���+�?dG ?̔��"���V9:������DN�a�!���I'53��J#�la�Z��Ѐ�w�p!H�\Y(�~�"p�4<�V)y���K��/㏃��_��:����Ƅq7(���ˆ聢�Rn����n������d���1��U�rB�l�DH1��Z[g^�Xgr3v\�����0-�L����hJ�0�(�}S%}r����k��ҬA�ei6G�A��:�.�j�,�<rt/��!SP�=hD��2�\�Y
�u!'7�,��~�����fT��kCb���ۼ�
�Lcܱ������A��
���DpZ����S�)����f�O�f�^�z�6C�]��6�J�رr5���b%�f�f�A֏6�����������C
�����q��z
�PqEm�k��3�s��a�����Z(s?��I��RL��
��t,��8J9����Lk��{0t[>n���$[�
IV~H����� �W�5n���W���h�� 5ڌ*��P��������"�����J �0��:���U��~{�!�F��k,&�b.�h^d��ֳD) ���x��m��Z��<`�j��v���1�^�Yf]�jO)�d�/���*/c��o�\Nak�aX�!���R�\��۪f���%�,!Ϻ����؃�v��m��B��i栦�f)����{�
e�xP	�oκ�"�-#v~�'m��k��303�J}��b&�V��ɪ��(��Y �l��7Dp��ұ�8M1���q*�d�!��8�Ƶ�D�vk��"\t\��#�n�&�A�~��E�L���_��3,-�ݭˁ�@�N���d#���5K�ȵҶ^Hl<�
|��Ov�4Bn� =��\w�c��6@>?���* ��\ƿp��%I�6J��� ����r���(��9ƻ��&{TP�K�HX�_���':�о�͡ڬ+��a���j��{���8e����J*�I����P�1�*k�d[=����s8�)\'��Kw��@�{�{`�T�#��.?�TTtZ~ �<��,�yJ�I�ut)W�dH�Q�^^��3�����!���3%�yb-uY�p�F01��>�M�L�?��ľ����P���#y��=~B
��~`i����|+�^��Mf;����C�f|�(���S3t�)	�Ո�v1o���h�K��Ϙt_���V���H!~D�L=Hm~���M�����\��>�8�6��C/��$��uw����Y`��FE��f��Z�wYlecEV�/E���'�{d�
T;%�����
A�V:�����ͷj���0V������T��D�SWucޙ����}"!e�&�Ƽ��	�P��!��"g\�H*)ߏ��|g��f��<]d>�ڳ�L�R�q`��H�[;$������bF��Eo~�T�_l˨�4dp����p��I�~�qγX��$���o
�b�ˌ��)8���d�-��J�t�4c��A*��ԟָ���p�g~֎{�����ѽ�)��ƙa��q�kan�V�.Bg��(�ŗH��A.��ɟ�Ա��u?�ޠQ�_@a1�}��[�D/�0���<>������>��w�0��BZ�6�m��dv���	OC������Mΐ�L��3G��|b��j�y'�&1F$�?ո�䃢��s�U ��E�F9V���������Kmϡ'ټ�3�M��MMp5��
p�Ҷsn���g�F3m��D�'M:��'����T��GU����B-I|\3���#D��?��7��#����yI�I����;.#u��ʄZ�<�xv����:����n���x�Z���/j�K��Q�ZXZX�>� �f-���xx��s׳Q��G�@� ��2��`n�3�NݕB�#uF0<}�������q}�Ozu
���`����"_yj.��X�S`]�+�Ǯb\j��8�1�ko�z��uE8��W��Zk�����R$��g�'�dhܝ���zK�h�^��?�7�bdh7�����	:�V*���̐��Ée�^�BQ1uȘ��{���Ey]�����N�}]���DÄZ��#��V�1]#�G�?!���R�����\I�ZaE�B���Qk��'�'��?{6.��[�ǎ������zh|�5���̈�O��fPe�IR�`��-���$cBЂ��~%�I��yl����ܺe��8�_��Y�� �o�2�>˓���9�,�B��#[_��Űe�AL~�A�B6D3�������3҅]D�o��ƪu�:~��@PE�Э�(�NU̇Ҳ`9~ĳ����)��E�"#SӢ�`���Dz�f��D7��R�"IM0d%��X�v��h����a$�Ʌ�*����g!C�X
������tzQ������rf��Ж2��5qm�� ����������a��I>� �fT���̂-��S�1m¯���^��T&���7bQ8��<�H����l�`�O��y��]��$�X����b�U�[%�n þ��� �L  ��k��d4
2N�2�}����Ϭ�=���f�Z�A��>5��	k�/�Bo7m���^�jHwk����+������Y�?�+/#�#���"wi�/�f���BQw��3���
Z��+
�U���3Jc>�R�5���Ct 9iƮ3��0�RkĎ���zd�&5N}9�@�r���StK��Y$�#
�f�e1[_�G��#�ϫ6PR����'��@��zg�&��ߠ�_D�**��0yI���Ε��͇�&��a��+vo{!��reV-!�t �$��?�WE-� � d�W��j��
sԃ�d�$-1gj�]�L�Y�J�X��DvK�Xo��`����O��J��@��?��i�UO·�������8�0���e�"�y�cX4��3?�j�\m+:��,Z扬�θ��+���1c�Sr�=]P!�fY��wd�����N�~��U��a����C:����!t�O��5��[NE��T������ΞΓ���.o�;�+��a�PzB-�nUaQ�э�5�oO�S/��~�a����.+)��U/Wk�4��'���$[V���i�@ɣVS��V��r�z���l����3;~�:$v{$ ��-��]>ց�d�y�0�E�7z:�
7t�����W<{
GaWe?��@����NG�mmB��QCw5��*E��[����\�1BWN�B�f�>�jgݻ�N�F&=K�9X1U��p�4(�oͬ�Z�%�������"�5��+�vS[��?cVY/KX�y�1 �\}��5v]߽z�k�;Ă@��O����3�0��v�M!��������΅=_Ȫy�8���t�n�Z:���H߶�l���C@h;�GgZQ�Ԗ�v���幫߃�<���>{�����n�>2�9�
�|��
G�	]�Y�of���x�URc���l�x��Vh5��Sf����Q�c\���p���!?��	X��/�)�Bp��NZa�α©:�IQh����E�%a\�P�^:�8*�Y��#38s�r���Ҍ��+>Q�䮎��{	Y�1ف^@����4,�oc�7�@r��y_�'ϝ��6/t�E������,����t�ֿ̽�����9A۱���s*���=�S���(�RPP�������+����y���cd��!����q"z��;���6jC��	�n��ߙ	�_�&K�hX%�y�\<'�]y���DT���6� ���唿,h)�\7�5��!��#��D��M��Z�)�*��u �{s�.n��С����i�<��:S����	Z�n���D�e�����QNI�I
~�I�A_P�j�Z�2�����ϋX�7�2I~M�yR'����E ��D�@>��ӵ�A���Vv9(�Zj�4�C���9k0z��֪#��.�h�� M���I��W�Y��C.| J��D��w$t�d?r�k���M� 2�D��w�D�8����Co���>�(S���Q��"��2;���m���ߓ6@��OiQu	iE�`Pe]�O׊��3�[���,е������z��� �`�����	�P}f�N�a[ࣈ�V1op:%���!D'� y��j���V	9�I���D��G��Qh㾠�-�K-y�;�>�t��W���?�1c�E'[\ �F�� 4��]YSoϼ���4�����U�H'�Nֻ��kcnY�
�̗��8�4k�eO����}h~p̺şIM�����TIc�>%��0�al5D+l7�o�V��M�]Q�:�@���=���g��މ�L��^�J�p�%���[+�e)?A��w��h�na��\<�oL�mѓ�S�J��V��N52���&�G��z��p[6Z�)$�e	�W˕���7�u]MD6�"W�u^'��Y�_Aڗ��qz>�Y뷯� �����_�,O��ر̐#��E�T����V�t}��5/�R8������s����>��ψyho��,�<TAK�+�G���k=��W���dݺ��y�:�Fp��-�G���s	�!sҫ.�{PUs5^�v�6/��z�aXQ�M�&�H��!Ip/��K�%�����M��o�`"ϰ��m}�7�b��N�	l�b�����4-E���a��]��F������	�d�<�TUA21΢m������y�`8��u�7�i7hb�.���4/���sR�)�y�O�s�n��'�]Ռ^5��fc�SOQ%<ǟ�.޿����T��Mc�zHp�����=�ru��&@�cp�0)�, 	R�1+�����X#���SO*�Sk�w� nD"?|�X��4	� BF�"y��bb����h�J%���ߓ�t�os"3�s�&�d��␄~��s?A/�|��s*
N�1H�7�?�phbb�}��P�����?2��Y�Sb��!:\1���2��N�`p@��`�&]s ���� H��_����d�d{�n���T�v!��e	�Ib<�/'�K�5q�3� �0l�*t� )����g���ٟ���t�O�����j�r����iR$��*��G^SU|����Z���2T�P���U�Tk��]ιR3�$��#���)M�1KW@� '��Zۅs��Nud�>��w�qr�qVivr���ݧs��3�N_o�[Db��]���|E�x�T7�����c�3}�6_o�T��!<��iH��w_c)����{���Ѻ%Kj�d���1^%���܋�#���Rk�1�;��d~�D�k��yfq[z��1�0�e=xd��m�,�D�c�ć2r����6D�G����6�b(�i�lɀHĤ&�TVe�����d��;i
H��JGX���u�8F^�"��Ko�
'\�W��8��CR�o�f��1B�f@�kʌ��ƔfFzJ�> [��
�g�aE\��A�q@�Mc��H(Ϛ^�a��� �؎7r�Sk���4�R�Ę��U�l8���
�@����a�>S�.�h(�P��ˤ�჊|�u�^��!�!kT�|����n��	�y�Rt#�ON<\��Q��m�H�U�#]17�Ș��d��L��TmԐp� 2��M���2���t�=8o�5�B�p�������y{�2(
:���K8�>�����^��TK�G����a�x][�4	2I�����g��*�������}�Fޭ�Y�T�X�|���URpB�݃�is��y���ֹ&�wJ�;�2T�����z�hy�D�vz`m��Mq�{�J���Z?a�dz"|o��I�z)�| {b*�^Hq#�N�����kV]�8�v���h$klVyb�Q�"Ne�1q��CX!���O�#y��B�6*M�l���j���o�t�����rŗU��^�,������~	��Եy!V�	�u�;/�����LJ��&h���Eތ���
Ev,���*�d�.�	!���8��$���ⶩԐ��Y�o�9N�߲�1_ֿ���m�3�/���	�ȣ�C��͢TPY9L��o_�/uW5L��)(p��V�����rT�U�Xw��6a"d*��ɟ�8ȂuT��ɼ���6[�`�YG�+y�ǆa�=�K�6ߘ�u�j.�ο�)v�d)2�V���c>Aru�E*̑Hܼ
����y�T�ׂ���bL���P��_�.�Lb�lK�:_�>�Q��G�:ir�`oF�ɱodw�ݎ��(�H2O-[C|v�w�;<P}smX�������:�k��Z��B�+�t,x�+�KI㿲��R许��I�׷�J���`����|�|u����k(�e27x������v̝YP�[x��bzsd�D篊�y��U�	ǃ|���>�nϒ� ���A�����q>�<��Q��|\?G*��2|�#㉆^�����F���<������C >{R᯽�z����F$�Ku)ħE>��a\gp�?��NQ�L��J��5�_���BvB)6��K.���cam����I����:�\è��ϯsg9�\�3��T�+�uЕQ6����y���XvU �Ί7�Me�Q����m
�u�ջ25�<P:pmqV�߳���K�o�)`��F`S��l,�L����^�F<�$�'��0A��~����'��+q�j�QK�Gm����D<�%"�A���84a/+����؍�e�n~�|3��=PA i�QQ�m�c�a�!8�ԅ��%�	L�7�Pv� mS����	��zs��������B�?c�����5����w�q�F����ņ"�R�Zm���_�{�k�j�3y?�a���Nt��T
������G�FG{kM��f	!�v���OJ�M�,�10%`��|�QT�E�
��v�;�Y��7��eU'���?�p;Vl�.��5��գ���F�g�]�9Ɯ���p{Gv-��4�Լ[0�WJר*��ڰo�����(A�v�	�7�J�խf�Z�{���Z����m�R�=�I\N��N�f˛���-��6}�{�p�ز�v�9�ґ��8$��K|�aH��;���#ݾ+��E/�Ym��A���֮���"˘����<�Hb�v�UOb�LQAtn���@��N�����>
�5�ͯr�?±m��(�6&=��A���ƑHw���Q!Ҩ�M��
N�RS�W�'�O�<ᦝ��C��r�	iwu�@&`��gͷb����ι&�A�b�e���e{O���HS�>���bDB��Lv�=���n,�h�׫w<�L��J�N8�db��ψ�Ib����@�}��|����sϿ���;�,%k�i�BX��ؿ���n�Ƹ�b�C"�v�{��*�v�D�-��	���
����&���nk#��|,z��8�B��7��Y�6���"	����4sC:97m��T����7�������q�Wj��wl4�Qz�����[$�v�g�D��'��ڣbM'X�e_b�����\l=o�B�@ lDM�k�@��N�E�B��Y��ʦC�N�YS#݈}I�KdlU�|c�*�9���@�����Τ55������$�r	#����P��A�����8�������$0@mjE�ё��R�y~�F�Q�p1R�k�v�����0�Y��>މ��m	/���)�����Z��[�T�����/F�`DM'�/ly����MQ�C�h��8�� �@�E=� ���%��ڻ������IE2GD�躋Uͩ#?�ەX0���g������,G�`��K����5||�[%wG��Ǭ��te�<�Q�,H��ޯQ�� ���@��z�~v�>p=���:�X�>��ɯ��&��#i�b�?��&��2�v-��s:1���K�N8��):M'���CƉ��<�s�G1���Wq�{O�4p=�� ҂&and��%�TC U^>����MΓ&�)���~x�@�D�#(~���b]:`��!s|qS)F��֧��Ҧ!�>���f��3K�&4���b��U����J�d�>��ȩs������3a<>˅��&��}f�L���6��Z+t�HN�k$e�QgFJ�=#�|��pPl���>�Xg=�k<--l����֌���(5�ו/
�����~�&�zS����:�#̔,{�-�Æ�(&�O�*w$6y(:�Y+'�����ëa��㉯���wF>9����b��U�K���j�x\3jʚk�2�A�����A{��l���	i�[��S9�ِ�Sq������rO�����7ٿN+������o[u�o�z��&N��\�h�U��Ҝ:~R���1"hY��±�@��e:#�P�[�}цz�a'rbf]�a:Ĉ (����X,�7��(�.t�"Nds|�%��ZX�_4��0���YZ�̇za���J�}�e��%_���rH�P�X.�S`�|k�u�
�T��J�ok1����_��2Tˊ��h�a$�&�e�'f��ש��K��.�����Đ�D)�>B9�O�����֍
������E���1�����\�2S��!D�s��sNZ��!whţ]���^�u0��c�h�f�Y���WNI��J��<B�L�Z q�w��Q8~,�%cۻ���,qK�]�SV����F��4�Q%�!x|���
�R1�,��U��v4��˖���/�v�p4|�}]�-IF�.� y��$��)��$|���X�@�C��|r��̻�WM _"7��ֈa,kw�I�>~�e�����1���O΋(-z�a�&p���rKZ�ˡ���h��Z�Yx��̺�tsd��N���E	1�����o�0sS��L���"(�h��&�W�N�
U��?`G���]FN��prh@�i�����Tl���H��o[��u��6Y �n!"� �q͉�e5�ˆfߦ!U�ҪS�uP0���pgH0U6|f�K#�- @��0�:����<~>ϭ�S"5O�N�w�(Z��%#�o��g�f�p/HI��Y�	�����v�|�R��hv#��GgM����ٝ�k2�)�Rش�'�4{d��y�J�&����ƙ{4P��X�~`�}��4�\{m�$�9;h嶏�!���N4G�u�s>�=�s	�j���}'_��rPUGĥ+Q0i�h��C1%HOtW�} ���Eh1R��t.���3C�Y���&�|��-~�Z�xY�R�M�������wyaD�$�B���G�Aή�m�{ 6>�}3 ��T�𺔠u��eZ��s�1o����^LJ��%�z1�ëf<�) ��;�S<0��,����l[0���~���>w�O��"�⬞_9�w�"��0b\D*�wkj��=m4����^vs,��)8��{ԑ��֤����:��6_F�`�U��=�sN
�z�՝M,��n�m�OQk��[X�/$-`�d�v�ו~u��)e���e���NY�x=f�TGB2��3�(���ȑ�xY֞ѷ�����:2����
�,�%a�o�J@& �[�zI2�m�O�c&�{��w��<���{Ǘ�EW8�!.$�ҟ��{'-�д�'|bIt෭2�Sh
��L`nu�tA��Q�Ol���ktp?����k%���L�g!,�_��ݸ9��)V�~�m^���(���m� n��<G1�H��J�@��cWLn�i�$�Wb��?&�C�Ly���.q��G����B��j���QI�������$f�0u� �G#��r�~��(���4�q���1��4->�kh^�}�9�^@�5k}71��?7b���]W��K�2r���`��؋���.s<��l=9�`�D��v�-��|�G�#��EW.�T4=�@�ɃF���+�d�U{_b˩����?�j=�)Z�:c
�F�-j�3 �]^�3���%@�&�W�`�07���8�n I;�p��H3H9�q�H�Q��_9Մl'�H�����5Y$wu���7����̈�^ԫ	�j���af�1lx!�R�ٗ?������Q�� ��6�H�l-� O�-휊�ѩu�C�y �{w�������P>�1X�!�-T��
iK��y)J�k�4�W$	[f��=+�����ωX��M'P������l�������\�;�T�V�hJKƼ��q�����4�#����v\"Bd?�v��h�$P u���҃&AY�'����	�0?#3Tǣ1�Hp#��u��@vd�N˽
ahQ��-�[����
�Z�՞�pz�}��\���5^u�'K��]�������}��P�H���<|V���3�S
U�L���-`4�cf�8����?�N�Q�M	��/��u*�)��┥dI���7�"+�!E �*�IU����}����I����7�Y�C�j"�{��;��DC��y�^������}�[��=�Z`�Q�EL*�#�@��soKڴ1��/�XQu`-R����nnX��V��C��|5��<M.I�����;��lƜ/���������3��b�#Py�;ȝW G�]�1D�LL���"��5����9�
�nHêEu�}j�Ϳkбi��cT9��pk?x��9P:���yPL�	Ӎ��u��I�('��(��/���-�r
>~¼hҊ�V>�g;@O���H�P�yʠ�/��6�o*bb�;lS]Tq��	���E��}���O��ˑ%vQ1��k�B���g�XmX@�6�9bK����x���Ҧы�����4*ղ�	�쟭\t@0�>�0���c�Ցޑ-��#(>���LO��9ޣJ/9�x���k�o��N}�0��j�QN����1�/T��+��S�h���Z)*�1�Բ��z>C2~~���'i}}����t#�L뷨���d+���;3u]�8�^ua9YN����!��y�f&>�o�Gf�D�'��h,$*�"��<��{�p��}PΪ���լ���Xk�ѡ�RӉ>B�A�}԰�v�/mi�<EՏ)�S�"{s���v]I=k�`^����E�����D��r@�� �3��x���!>�����g��v���f�+��;NWi������5����闓؟��]C>��_� ����U#yPG���Z���h�R5{T��� ��@P0�RC�.�&��X�mo�~].��7�����'��xjj�A�~l����?U�ly��o�mm���+ư33
I��B�Urۓ�Wou����S?,]%�]�]/�����)�\I�!ozߟE��� ��T�Krz�D-sn~W�4��d��b�v�V��V,�'�\>»X�r�j/��W�.���-%{u��>!�YT�X�;k��2��]�����mNڐX"{�XI��ld�<7��42���`�%�3V��)��-�Zԕ
���D�=�n���H��J=�g��%je�ݗ��<LS�J���[!��q)�^s\ۣ��p(5kU5��Ş��t1D�\���eP���i�z	��_n����{6�q��(��O�U:bՙA��ޯ�=:�J���*Ky0����?՛��%A�k;V�N�.�\�{K����@Iz���K�R+3EƄ ���@�ڵm9���+��ֱchex �qc
:,C�FV�	��/�f���������]Te;�n(�A�e��G�����/w��V� ����^,E�r�dc��/�j�n��h7l�=&��R���&�Vs����#�>WX�?CE����^�хZj�b��nn,�G����;��H�os����������d����6 �-BC��{�EzB��g Rhˇ`&�Y8���h�\�ް̇'�t5��C�@+>j{�G�n�rO�I^=�+z/�s�6�b�b�Enr��� f��w��%sb��?)����Ԣ��)���2��F.����$�z7�d�!�[���M�.��ɶL�0����~��������*&g�����O�O@�
E�}^��x���^%���7�g/�)��mV]��ڔJ����Zn|�o�nJq��6N�@�)�_ж�N���=09D�����U�J��A)c*����9:Pf�Cs�Yg_A�*�s恢ɻ6�5�����{f��qT�����ih?:2���~&#���rχ�h�ou��'h��i�G���|�TRF;YD�:8�K��p��_�b��E�/�[�k�tʃ4����*�"Ě��#����kا��w�gk\�:R�GȻ�%� ����9�H��+���K��)r�ɲ��U�H��6�\KD��54����uG�li�/{=gp���a�*U���o����q�s��ғ��V��5�j�+�2�#�e�g�W)����`QKם`)��ړ����7��{\g�*��:�x��T��bR�]"��9j`�fR���&+J(O�G�0�fk�s�u}؍a�&eT�$*JҦ��)%3�|��v�`Ш�a��7��6�;^a�F��_���]�H�."�x�`$T!|s�4�M�q�<;+���CƟ!�^rB��E6n[;F��cT[~�m�咣��{*]�CkV�~���h�h�u���o$�N~��[��#{��/����솀U��ەx��l�vM�6aѿ�t^a�|L$
���b��ܩ'��zd�->��T\��lkw�PN�M��fvϩ�������M�(4���0�PA�ޯ��K��b�PW6�o�&�v?��"��d����kpp���r=^�?8���3$��C��y���B� �DV�w���(Y:�JM�Y��W6*x�Aj��=�;��~�:o� ��PX|"=�Ͱ�)>�X�2`K)u������1�я�o�S-։��PbtŃ]yu��E��ձ8q�&�<�Mh�^��NwQ�D�����Q^Ԭ�"�	¿��3�j�'JZ��q,�k9@V��8E�o�~�vN�6��tE��C)'��]s��)���̘D�( W^X�Dmu��;&rp	�b��;m3���n��{���^�_m�} ����{w���t���̒�r��5M���:"�R��	�?�k)��Ȏ 6|��m��/_r�?��U�*^�Kl�f���,A\�h��;8�9��e��P��㬜6G�&���t�V����+	�sՖ���� ����1o�,���h�����cGLM�`,kSK2�٭c�ˑ7�`<��w[�lAU0V��,��#�
���1/1��0�L�Ah7[�T��Z�  O�d�I0�m"���v��Û�h�S��(�����OF(��i^m��+�T���{�beDH�����P�v �Ţ��5!�z����k�<�,<}��v�q��"1������ ��~�-wڇ/�`B�U�kt��أ�7�+6*�iY�������qў� �[���c՛� ��E��50�,�eh��S�S&�l^qiмH/"�ӭ�%X�Ԏ���G�%0��\ ]�Q:_��sub���7����m�2 [䈫1Ix��J�+���f�ɹN/�ʾlCU�+�ͯ%����D8zud��
kw�`$*jē�?7��a~׉!6Ȕ>9�a��3�6B���A	��TGca"s�����^w�=w�}0�)Ʀ��h�B��k�7x���F�}�l��1_j�e� K����L8QP�I'�_>���I�zm�E��aAK�������LzI}�ѳ�~��2Ճ0�ӒX�sx�%��l�_?R�k�V�ld�ۧ1�a����*�߸���y0���]���0��*1l�m�	��f��_:z�U("k��!�m���V&1��i7h�{E<䤈�������Џ&�%�ދ��ڡ"M�hg
a@��I&�w)�-�X������E�oV��`�µO�u�F�I���h�����!�L��~�L;��g����D���F���N7���ٟ��xe�ԕ;��,�E��+��GW�墆 �9��F���'5����83	7�u��4ҝ���6�`1~��/>}?TN�[3�K�E�h5{�Iۺ(v:k����#t���M��O5�K�Ջ��Y)mN�zK�\�1�����[J)T\����ʏ-���&��S�p�ﾇ�߮��8P4�����$}[���̵۠�z��:R5�#�8��y)'؄���CqZ��6��t�0a|�LQfaIj�KZ٢�O9�l��X���^;~��9��$�6����|�6e�F^�۳];pSJ��^�A *�?.)"�}#
���xs^7<����=e�D�#0 �K}Fo�O)J�7-�O{��W��=�PPVh�#�9E�E�s��.c_Z3��� �:pd)G�ߐ��憗�2�e�������T	�졑{�����uq��Ѳ�V�2(�'9�����c�?�/Tֺke*o�)9�b�Vh�2r���Pt;�Zcn��;�i�D>-�}%(^��࿦�pv>���?r���̫M5C��`���ҭEN���V����Q(0�QZ�}��.����_���Xi�&�
���K����]�
ow:$�9���x� ���mf�D��*rn�A)Yu���擝�o��僙�tո僠ro}���c�~b���;Y�؊s����\���G�iG�j�0� ����4�^pA�,����d{�|XFm����$w8�c[���Tk�@�"5�#���Ct7b��,^��k��Aـ�(��ɿ��<�͊�,�\�uGhWڛ\�B��|]�ʴ�V���Ŵu�O=98���nKe�����;�o�Fe���t�/�?S-�Ԗ�����L����)?0�A��ko�93��2���jj�8�T�;xA���,ժ1�	�� �X 3�YE�	���R_�NL��Et1$��.���(���o��T]��M���ܲc��B=���/͒�����@�=�w�h<�{��Vp�ct1���� b��\i6����Ҕb�Y"��I��� �;J��W�Z��>�?������#�B�������}�&|��#e0��=7/@��+����.{؈���jo�)�h���e���Bʤe	�L�8�{���I�(e����*�����nvjE>v4�N�������?g�{����� �:���=�0���6*��ل��&����]UK�{L�.�4;qF����U~6�S�KE���?��<�Q,�N:��@Ʋ]�wsNRm�q;��SB�N1��7�u!��n�����BM��]�	2��3����I5�7�<�L�P/�}q19(�T��^��ku�����@܊��2Q���;u9�K|��*tNe�����6�����]�Xz�������F�(V�Ln~�iDlN�t�Ǆ'��?�R$�]k;�pѝb -Ys�Q�Й�舍�V�Hj�N��		����>[\s)l�J������ݵ���+G$�X�	UEE6Z.�wu;a ���-�T�-��jW	1n>��p�z]6yf��^�(��E�J�����0<@���;��p�8�1XI�mB�||X�}�kt9~��n��d���΋�N�����7�^�&�fXVu`��Aᯪ}D3KIxQ���Ǻ�S �LH�;'�YH�6�033i⠡�l�3u��+��f��ʌ��4�8�#�z�U���vV9�}�QSj��Q���"�<nv��]��.�ɀ����GYιR��d����
�L�M	����j�'2���/AH���>h���s��ؙt_\<I�S�<�'��;��PC��c�z�볁QI<0J��>l��/�*��8S����b����H�s1mIA���B��%���z�%!���YB��I�yvjb�DLh��,�Аs������~g�O��&��ia(~���]�!*2�2v�g;3�/��gTG���Y�,��:�tp�F��������c�Tk�R�dcD:A�я֪}L������°Qc�X�"B��'YRɐ�$J�E���)��cR[���"';qq�� .�Bb��=6�Ł-���	�N&�B� `f�uM�X��Gy�e������&�kP��.�ǭ��1�	�s[�1��3��y&�l��0�_g�����f/�V3��+B�o��<���9��t�k��{V	p����u�ZQ!#���%v���#��q��l4���]������*����s�"�f��5
��tQ�T�2��s���\䅴�Q�4�~����.���f3��q���������&��Ӕ�k
���T�｡�qQ���)d�̆1�#&0gU��g���Ř��v��ɦ��oL�:�u+L��b��fR����9Fj)e�+J��Q�󲏪���,MhI��،x�kMl��U�G�o(H(�vYbx8��qb�򆼂\�oK�T� ���Z�"1������&U�d]6��JV�RW�m��i)�&��
7�VS�Q�R�]��+�8v��������`+q>�)4�ש�C��QL R�yu�!&)��Q�ip㪩�6)���|Śwĳ��3��(}h�
#�&� ~���N��Sسi���G��[��bO�i�h���q!f0�$v4T̞��!񈹿)♉{"��&_�Na�`�s��ec�<%��6���U" g�pSkF7�ѽ����R "}�� �U�������w�j_�?^2�x&�BN��Y^�>�(�D���9����z��)�>|�$�+PW��a�VnED�:�8���W_����J���B��djj������*ik#Sd�F�<��Y؉��) �L|c��i-vS[�V�ި���-��DS�𽽢�jK���b���b���ق��[S��%!�_10-�At�C�o7����w�w��gsm���6*|:n4��崌V�M"���������I+����&"�w��4%�c���sO��ĩW=7�ӶI42�� >sP�i�փ��EP�~�% 4�O�O$i���B�l�ه�k�"X����Ȝem�:q���R�ed���/����K8r��]��3�N�V��3ˎhR-��pL^�M��#�>��A�z-��'bu��H=�>�@;g�K��ZVG����6m7CO��q�+fPPo���������<{~u<o^(	`�ط���-�,Y����ǂ�og���YH&�(�Pz��^H,���¸@�*�n��$�>(!��j�+k='��ݱs�xp�9F�����Q��dl�C�0�X$l�ᢳ`cȡer���%B�<mu���Hok�����Á���N)��ɩ�ͶS�X�*e86ٜ�3�6��Q	k5����F;��9���)�G��Q��0�>A�m��zYJ�F���
g������5��ɖ`�v��t�3��1�R�E1���*H�Kgn�dy��g���"G�&��B�`�P���Œ�j�׹���ae�k~�d9��>���-�XN�$}Ũ�HƟ���Z�q/&/�2�A�Vݺ����A4��.Y��st\V\�(�,#,�xȂ:0�6���+�ӑ:7�ؤ�Mv�شRF"�3�R�7 �t��U_`<�&��|qi���&�}x&	�(1���/��|�̈́��Sё������b1]{GF�J�sT"tˍ��K��b��h=Q?eg'o�p��oT�'Y)L���=���uz��L%9WkzAoHڨ�H������q�1m�&������f���T�n�磎�Jr���e��Y���6G*�E@\x��"�Է�F���8ߜ��*��%/���_tТ�P�<VA<�(��+���Q��	]��&W9���w�.�C���h��`�/��{�Rt�{nW�ꊽ+�O&�G\���o�(z�T���E)��H�$�M���/>�R�Z��Ì�����or���9r���W<(L^B��e,�w�̋����LOZ(`�
/��Q���������a�
 5q �@ZDH���/<*B;ƙKH�g���flA���k؂3�B�q���a�T甞>���տ/K�J���I�>b��Axh�|���U������,_���k^�	m5�H��������t?N�Q�R��{ps`29��qC@Y��te� ���l�Pl^�m��:���K�j��4��#����w�{r���]��Ș�[�E���t38iCeE�\s�,)%n}���8����v]:�);��T�ٽ�ZX�mʸ���>U�����=U%�j�p)�*��k�^C_4�-QS�9�s9Z͍pW�
w���,��C�5]�N3�R��ߴ6���?;w<�?�v7
�=�o�����3�1a@��������S��3�%�c�Z��x��ًfh�B�'�w;B��Ҋ��������h��=�#��X�&y�U��2f��;��x���$�����Y�89���?�:�^6a��^yd��R�nq��*�i�"O����S�Ż^3SΝl{�K��7s����3�d���m����筌�8�.�Z\֖秾��Ҳ	���kv�U�����2J��'�p�g���.�9�)v�vA-�H�q]O����V՚�eY��W����zOb	rSLGu��'=�1���"PEE���m͵��,��O��BAw���K��1����G�A�!O�;L�q���k]�U�V�r�m��"��cq8pK�)�aJYeZ��3�u����X
 i��&#�s^��7	Dz۶��:��N\�+lDef\��ba��r޶��]��nk�69U-5��2�]�Z�*�o� �%�v*��5p,9W-1\��e�u"b�Έ��k���i8�T�Q[`������'~�+��rzsZ��E;HD?j/�	��׹�7�\�������lv��/a9i�JY�,����qB.������j���Y��N� �� �HS��>� �]�G�t� ���r�˞��C��x8�v�#;a"� ��h��i�e�%�O�z���n�g�Lt;�憑�,���Wՠ�H�\ :@���5}-�"�� _)VP3L�Le���Ә�tq¤�^����:͢ZJ5��ՇS� �s�Vr��,B�ﰮhWw�Lɵ�p���/}0��6�x��v��$����ĺ��nȚ.�C.�����_�$q^���^錢T�+ё5��K�J ��Q���Χ�C�+���9�z4���g��������8T��dM��J\��������'fo�G����c�q��q@�+���v��n����� �H%:�Ɠ�| �į���~"�d�P������Ĝ�r�����W�T����۫��o�1~y�"���&*h�M��4Y\2=��zv�gf�NS�rh��sL��Aj�dy(��X�F n���?ۤ��d�¼�P-�g+0���z$c7i51��m+��B{u�π��d��]OȈt-��k��o����y���=B�����A�u��՗)�SG\���"���qp��x����
�铲+3�ײ�Tc+n��/`<Y�����q�u0DGE�}���<p����PXĹ�a�j�'���5>hr�q8*�?ZO��;\A(�v}!�i�=�p���O�*5�rB�/������ڣ��M�����u����h7�ᨥ8>�PL!�AL���W����F	�:���&�����h��h��9�jV@'�#�8�A�/̋;*S|"<��}
 ��?M��X[��	y��'�>Z��?�X��?�$4W���8&~�G#0f�Wq8CB�Zg=�����n~i+�b�*=��,Q�ѱ�'���1����3]��Ao@�����8c^�)EK��s_�΄�V#$�،�Y�Y�j���_-�,���3?��S�ȝvg.S���wK���'r���v©� ߟrD����_��d�P_�n5
$�����v���)=�0�QS�vN>Y
M��%gK��e�_xF@ɽ��H�;���{[vs%�3�������Q _�Y�b���"gʋ�ǻbHZ�t��.|� ��4}?��+"�T�R�`˃
i+�K�Dp' �!�Hθo�3:�VL��ם�8�e@U���Y�]<s"O��A1Y��Ŵo�¯��`�����'��/m=�|ĵ�ͮ'�l�����vr ?�� -��1�H*�r\x_�c��y/+#�Ж�6Y׭\�طY��;����tk"�.��n��sh"��{8F��T�#�M��9�2Y��8����&[�	%j
���V��ة�:�����k��њ	k�X���4�1UX��e��r`���-y0� ���7U9 @��_���G�\��t�vBy�|ы`�nZ������qe�4VV���(�Q���v;K,z�V�I	�7��K/�
��r@�*�)��)���s�G�(tT�I1S;f�rW�fah�������eB��y��Z�CUb��O(�x/���Bi�bs��hYƾ�8���Z>�b/�ܘ�-�H�S�
݆����.Vo��XNW�	��6�?�/4�,�7 �5�����|������Uk���7,���
	��;��E�G���j�oĭ6w=$�຾@EJ�mѼ�nhYEĳ��|�)�v���c ����e�̬��Uϑ���"���t�F��<HdE�aw\9)J3{�nh(u���16hL1i+C�v��h�`�Z��0d�"���Q�T�S
Ĝݶ��_U�u��y�Sww��rU�A�ˇϕ��_J��L�lL����&MM5Ì���d�7�'Q��Y��j+}�L��O��(�%���Q?;G��f�Is��$+üJ|���P�D��E���t�?8:Ƚ�&���qͱ����:E6/DH�lix
H���k�o�X��gt�;z 6
@+ƻ����U����r�χk@V��|���ap���`�^8�N:�/�E�����}H/���sm���;$b�GM^*c���I�eIZ>������T�|a��z�k�	t�X _���K/-��Hl�:a�]v6iPT�|25�Pso�^	F>�*�̪�r��:�#��78��-�M�R�.D0yC��L�U^��v���oF~�!����b��$<l�f����0��W�k��M+�K�'���|�gh�\�&��W&�SI��~��z�/�����x����3�0=�L��#�Ar��k�P����:]:6t�!��ԑ�S71ǟ�n���d5��!�}r���;�"a�f��A%�˯�}�L1^`���^���.ߍ~U�m�4*N"��� ��`�����l{�S���[ǫ�,PU!��S�Ϊ��٢�;�rN���ى[��ެ8<fS��z&=�(��E�m��+�HG�Td�1X�q�_0�*dՠe��a�7�g����.�O�x����"*���Wy�2�	�ɖ��>�6�� y��.���&�%��F!��6t������W8;���Ŕe^7�P�T��r�#�p�/�y�����;u�b��x�L���8;#i��B�^�A�振�lq�{�V�^OZ:�J[���>�b�oǺ�UpV{@A�� B�I�k�ɞ3��H����=�j�{��#��=B�ηeU.��W-��tG�5�J؛ߞ��x�mԡ��X�Vu��Bv-��S-�pͥ�m��Gͱb�uY��PD�4��'�ɚ��DQ}E��W��O�J�"El�R��T��vk�(������p�̪��1�fJ�](�fI�O�@ ��ٞ=�@0��h���/w	ب	�bL?��^Z5�V�t�`��D�k>�6f�㑅̓�bR��+y��TVSq��!"���� �[�u0�mP�>^���FJe�(�C��wA��j�g�J|��k90'R��|�p9n���g#%-�Jw6ĉ	Ӡ����7s�,ѹx�Y?}g�v�Y��
*]O&'q	^�P���}r6w�j�L���F���n<I�FkÈ�r�Aߙ8�l��q��s��0�۔V��l/h5;��$�H����]���,�������
�iv�7mZ�sa�;�����a	�=�Ag9�@E���f/�܎�]���)���p��/V�g��fٖ�*#��R���*D���'<K	���=x��E��������[��B�Q=��;V���Z�2��|n�~�=�)[�Nw�I��3�F������2t�F��HΆ�v9`�D����[�$��K���D0�y7�k������S��
��O�p�͆^���e�6ݬ$~��2T�ίqb�T��naF��܈+&A���w|�R)g��M�1!kF� ����㔂�a�[Xտ����������0�)hh���t3U�ާ��S��8߲f��+�8|p{�¥n#�ٸ��ߒ�a�ێ"�m�R"U��Xq��V%�#(	�n�y^��S�(;`��d��`������0�-�g��r��a\�\�sm�j��x�)���G��]Y>�Z}*]t4{�W'�;�fz�V���{VP�T&\a�y�4���8�+�{n���W�L��G�c�Gs˹%��%7VQ�i$��jW�*^�ʗ�a.�8Py/x�*E����>�u�匳�q�1��|�P�����&
�<ͣ	w0,
�Y[A�y��ԣd:��ʃ�%�Ō�9jG���[Dۂ����Gs������*���L��~`?Ep5]�
�	���T��a;8 ����:�n�(�n�$�P������iU�e�U9�77�=�.��0�-�o`f�����Z'�-�}�+Z�������V-�\ʫ*�o�6	k��b� �i~)�i,�L�{2��u`�Ө�l�r7;��_u�����*�L]�#?tH���e�@�
W��g>�I�I��=F9~<=�'��-��s�1�py�ʵc~:{Kk�����y��l�D����L�2��D�rA�i�O>/܋ћn;��!��hv�b<VЪ�l}N`��"H�����p�:������ 	�2���8ZpqI�p���ˋ\�p)�]nK��u��P

%>�W��UQLm.����~Jwn�D��8���ed��w�͕"w���UbQ��S�p���['�d�W��"���w!5�C����>�F���fs|(e�9Z��LL_��ZGN��Z�B�0*�������@�qgQ(��/�uً[Ϟ�YI�/�Ku�����ޝ2���x�%�����)P����9�V�w��J�W�aˁ����k�<:t���8���/g+���8��^ީ�R��qz2�Uc���8��͡4��tf��`�h:|��)
��}�|�Ƃ������U�Lf�
��7�C�v�GK�L�^S���6��z�MCN�˷���:<���e)zW�I�}�/oE�L��&%X�q�I��5߼Ic<#B�B�\�~W�����=���2�O�����%�7�����&�N���Զ���<�ô�5!ܮ���UY�L-nT*�җ��@ߋ��R��b5Qo8�=����*f�C� �_/ é(���Ų�I^�+�q�	e�6��N��
,�(�HT���廦Q��^�VK����2�QE���]B���rH��@gz���ˮ^�����W�ML��~�������
��_t���$,�r�x��a�;��"[���;�4�����G:�	%w�?=�5b�S�1A6�l�v�8�#��2��l%�O��u�-�4F[�/0�=�>��o2��>j�T�)[�4�[19 �Z�٨�*�N�W|��X�&S�����b,3�-�/��ޫ��qXa�9�k�&�g�M:���VY����c�����M?5m`A�$��%;����K�09Q����~�y�tl�"HR
)�{6��a��,M��A2�޻�4���D�^���<p��hѥ��!���޸��A����W�Rn�d��RE�+����;�B���KE��IvC^Y�b��>��e-A�E��;x_x�4HR�R�13��bɼ~��p���ǟn����q&��hIG�>�}ul��GN��
�����!��jl�;!���y�%D�D�y�f`I.FB��D�fC7��f}����n%O�Ќ�$��M_���l���\����6f�W�����* =ZT��{��Lf�.>[�0���h	��h��e�q��񟞝��0*��-��0P?�d�Ϣ�k�a�k�Ŕ�v��Q��5"W��yJ`�l�s�R�i�੩M��ۉ�)3�Ͼ��Ġr����O&�1��(�W�U0eV�
�yjW�Aڿ[9M
o�GqW'!A�;0�J��~�'�B�*��ѧ~�e�_��F�N[MOb��Β�q~w$��"�m�/o���n���`����#*���[<�c1���v-ΰ��-2�����5��!���(qQC��Y���7�i��I���J��n�U]�v��p�l�R�������`B)�<0:Q�:`�AO����P�]�9��t���/{�t�A�P��-҆�[;j�(OR���%��u�7tF�9w0��+�؝pU�A�,����`U�]�s[�U$\�JÁ��R��	\Wn�OO�.��;a܈K��μ�����[ugy��z9��-E�U\]�)��Ҳ�P�lF{4Y��7��	�����N|>$z���2��>}�{����h�ԑ��䫑���������'5��@a�f<�����Tb$�c/�=b�>p	T8:�ֿ�����W�lR<V�~��-�K
�h�q��7��̫FL\��x}0n�V���/�Z(���7H�����ᶆ\_Mg�qG,�3{Λ��&F�����˗��6&il���z�B&_�3\���A��-�ڞf�G��a\ p�s�cJFY�@�DQ�i�8�M'��XK�,�p�OZ;~��s�4�QM�,��Ò���$4
A�W*â�߿{ۈ�G�5�����<��� ��$c��h"Y;:u8��8#GI�-�ɐ`~��l��]QߘJ��!�~L�x#8���T�p�wr��%���-,�.H]渊���8X㶧ߡ?�$�5/4��\�6��ܣ��}����i2y�T��}7~�-AѮ�w�ao!����ُ�0������0;G�a����E����Xӊ 1�bl|�j4��$RQХ�.�໭:�E9���ӽ�'�ð-����ϸY�$�(Bⱼ�'.=���OB�Q�����C��k�ڟ�G�~�(��4�V��0�Õ��L3(�R��jQMX�8�j�Џm��3���k���aM�6]3�W�p����D�k��a�j��D@�XŢ9w��O�u�P�Y�c��o�N��j����4� ���7�ƪ>Ӡ�����_1�d�"3��P��[�,�_��;�Az���)�~�]c���Mme�M����k|��S���c�Y��gK�$5X���|A�?��+��1��RLb�4���S�1�	vRRgNխ���~U��,[�.f�0Y`�$��T�=�x�T6�Ek�9�1�a�0n�B␵S���&,�_F��G�cI��s4tm�k�0k�����;���#P���ʭʙ��J6t��GUe�mv���a:~�q7�����=�5)Q�����^ȕ.�����a��Nʌ�)��̛�(V��J��v�v�d��Zavgy/@t��եZG�6#ކ����M8��ZfsQ3�M���ue�7�D���X��!�jr�^��JC�2J�య����^�ǚ�|��3�ro�TC��'���������I�������3�#��� ����\����Z��7����[z���fn�I���&���ށ{U��� ��rF�����Da�ݗ%�:���I�R���qX� `\��C�\I$��I�?�
�O�+��&�_֏���F`F��V� �GĶ����kˈd z=�l�V�y�w7^���G��[������~`C8K�LHBU~�^����팸�((v|t�n��F0W���Wx3��R�>9K�R:k�fbm��O���29� ���������|(�.5�;��ۺ�nd�L��~^�b�>�6X
��Ff(�K��6W��lY�
ٕ��Ma�9�QI����k8����n˼؆/~�Ky| ג�J���?kW"�)�@������r��p�����m=^��P�D��C��� ĭ� ���K�|��f��=�N��a13@����.� l���,9���5��Q��zP��.>-���ζҋ�N�i��U\9i��.1����]�t��B��<d���.��{CR?/�V�c�u�D����Z����l(l	#��Z�.�v�������vϣ�k��E����/�f!]�(��L�;���T�g|��K�/c���&�Z`7��m[����6W���n��hQQ(�"�9���@�a�#H����Ь2omaD۸L=��ܰ�6�����Apfg)���r���)����F��կ��8��]�:G��:@�M���-uj)-Ʀ=���L�9�7�v���^Ք����'?K�T������0��P?ҝ�-���q�,��"(����5���)KQ�N�ݧ�U�5����{? ��ށ38F'8-�Źs�a��(}�2
OC�:/�ն,��gpE�+(��xc��Y"������g�{�T��9�[J���Br���\� �*���6�̗�G.$�)����oZ��� xSz�{���(2܎�h���gX��4�Z?g�X�0u���*|��[�!WՔ�cFc~=3����y5**�oEc�
xz�'ˇ7'_ 3W��LB��"�V"Jᅋj�<,e����VeM�9RtG���X\��Ď���<Ȱ��<D�^�f:O�4�?s�ډ��K��_�"E-NC��	��#2���ܼ-�Mő`0��� :Z�F͒�qU�k+뙃�DH�����Ż���U�ք��5v�͌)Z�Ģ�̍�!|@��`���tJ��h]��ԡ��r�H�B�����w	�&}��\�J��bL���&��X��pd�^��x46YE���Qyň�:���$AX�*~~4N��tm=�غ]�۪
�|��9���|�R�c�]/��C���jC��L�Zr{t�N^���_ts8`ߣ"�$�������<!���B�2��\$2�Ѯ]s�:�Q2 �5x������TEz��3����R��6[�.��XY}D�l=�Az� �w��i�믢�+%������G/n(#w��t�;G�����7B��Ӈ��1�9/c�Tq�U/m�ľ�(ͅ�K.-fÖ��D�\��+�4�ϱ�9"��s���`��[�F��$��>D� �����~G��E����FK����b�;q�r\ˡ���R~��b8�T��F�R��uց�x19�k�N���G�!���Ca�38Q��k'өt)�`EYK1޸�*�hu��(��!��l�W��vk��\2�T���+N/6G���tB��|+�p�?z�S[j,�}��4�n+(��*r~o;4b���i����d��D'"���&�D}��)�i��X�;\%�R )�:�Ok�]��;Vo�pS
�#��x��L�FL�+���q���c��e��]f��I�]4�lf,���Y����(��`3S5�+�U7�4��,ZX����M�С���
_��{�)��9˦:	'0��� a}��2eD8k���Hx��h4Y0R>��<>u�<��/�D��`n@� ��b�~��|�b���(�������n��?]h�<���+���7mWb:�H��nWTsK���R�or�����?C۳��Nr(_��0H�F���`fT���anF�/__��S����U��sE���&���19�w�
��5qU�";��S/�;�&	��Ǿ��7hR��J�I�il���P�(ζȺGjx�����7��G�q�&A�
 8on�Q���d�Eu���\@��\�[�V���k?.ډv��O�AJ�Vlq�5�}�����&�Ã,Ì��H!��eB�D���D��UN Pڧi�ۏ��cw��Sו~��{NNw0�ݝ��47��M����Y!��
,(7��gR�!!�,=:aF0>=����}�@��㉔20pܹ���4)�Y�[�[�pQ��0fiwr�{�B�}:�J��M�eR�a}��b���+6t�WWvs	�v��7I2ָDص������>�;�Q��a>�;Q���'+!�ﲺv��u�0��}$�n'�PՖ��<7s����z��E�j��G�.z��l��)�R��K{��d�<��T�6\�t��<g�4]��� GD�|&����.�LV���p�����S�É�;:m;-=��Q�*TtT.^��u?��Y���	�G���c�>�^3��
h�Z�5�dy;�\�Er�5��>D�3T��BeѐP�*��`����,]�_C�k�7�OUs ����&��^ֺ�Gu\ ����S�3�I�	��0��s:�j��Ql�}d����Ign�]n�v�iL��_dl��REJ�v׾g�E��ښ(�p�j��2�-)��n=�E`U ?O�w���Z[h�m� j�.��l9��d�{�N�'t�C���_��o�S��y�%JDRՠ�xs$�Y���n����Yj�<GC٠��Ig0�����Yz�s���f �-�6���b��/�����L�*6��V"�
����1�e�2�D�^$a��M�u��;���.��&��;}�#�Fۭxzڍ"$~X<��ޔ|��������a �`_�6�鑓A�';=�β�4,:Y4p�A4���7Fo���.*���a��X]�O�tL��>Ux'˿��_���qx���U2:�1�[�I�MCђ��c���	�;��z}�V@"�����Uۿ)o�Q_U�l�{�X�(*`T೉:��Y��Hp����[$��/��+e
�2����Л��н��@�L�]]V�����M�*MO`Y$Ha���c�,y,[�����=�א���0�	�E��)q|�=��J��7;8�Tv���~�S���E�L�-a�4W��o��3lL�Q��+��ӂ�ٍ6 ��h��̬�♧��6�y���]��������;�N㪞
P���u�*:�)��d�tR��! ;3�K�� /$B��+�j�|�=��z��Td./�E�����k%ɮ�ؖ�ޜ��uf%�hb��=��,��+G'��t������M��b o��E�Q�}՞��n����aO"��\��H�71D_�E�H"^_��e�c��b��#�&Q}�3���|��F-'�����O昑�A�E���"�`|/� ���.����P��|�L������
:j�J]̶_� �k�C�2�����"�E��ۀFMhti� ȭ1�7�㖝��}� �wi�v�97%���i��U�Tiw7��`[��)�� ���nN��k�3i�:��ޥ��I���*<�&	]_�y��]�b�	E(��Zˀ��ڋ]u;�ӂiQ�\�*�H����T�X-�}�Z��8�[t�]C'�_`�
��e#�=���=q_�W���"�<���\[�N�PL��|'Hz����渥���+_S��3��Zz�g�t�gRh�V{��a�������b���"r�j��R��k��џ�Ѕщ�R����}�"c�t�y��1H(T���_81�$���x�<z}���iu�˻��Z+>�M�?����޸�J7�$qf�y&����]�i����Fx2�-��U5��ܝ����"�72ݛ�X�����4i����]&�H�n�G6�����n��+���I�YK?�*6�;u���Q��c`z�g�z�HӉ�
ܑ���$����|���KUk��i�<�
{n���ۆ�`��[&3��:�P����y]�$gX[�9�'�FRhygP�m�l�戳����H������߭���.Ywp�_�`<�Xs,�C±�{�Di虺N�b"��S#������k0Qe*D񿨍S+=�
C�����k����N�F⵶�h�ŞS����\ݧ�vUm�_�2����fg�Y�	�c,�+��Aէ̏oF�o�(L�$�Drm�?w	�aRh�]�y%٥������S_�J�#3]��@��/��R��w@Q욎q!��_���
�R˪��9S4�9���Ʈ������s�~p\��2��|\��kJlz%c�!�WFݜ����R�WO��Xn��C���YZ��$�M�31����ܞњ����v�q�P�h�bEg�� �V��� ��\r�!�h�N1�mA�r}��"��VD�A�~����z��\g�BR}�*���GK��3] ����g�����|�R�B0�z��.��T��9 �wva�!�tǔ|��\M=�E�2��9BOj%�i���o ,|�v	G�6�|x�i�C;0\�bh2��Ӳ����٠驴�nݻ�ƈO�B����[\�g���@p�Ɯ��>�YͶG����L?N"$�'�� 
,��00h󍉧�1��.�~�T�s`9[G�g!�.ơ�����ى	`�k�ơW�:�>�_�������`�o��g
��O��F9�"f���705��b��Qҗyq`-S�����{f����π�;>��A
ԓ�߃��L�N�,J����8�X��UV!��U,U�l��C	>�lXb����v?�k���K�����=r���_Rǚ�8W�g����J�����lj����WW"���"5R�7GSB<���D�	��Ip�O����D����Z��`�b(�$�pb�	A9}����:+�
���$W5#p;C3TZ�z�}7bU�ש�#����Ģ���d�މ�?_w�.ك_�Ü��V�A [��>ɧ��@>.�x�X+��^���竚e�cn�z���<�f����O?�'v���	ת U��t����T�&:X[t�0X�1l� �|�B�lH?感��S����m�+�T��H�U[��,\�?@��E�C���F��A`�l^ѿP�H���3���Zg���B�X /j3��e���	�s3���Ɠ��^�����o]c�0 ��E�� ҇�3����4�"�������S�����F�1𮥛�J��J��c�������۲����3Pr�KN@�����pH!*��{�a./}��{�id^d�{��7T�h���)��
(�e��J<t��(:�U��>��5C��i��*3���38�m�B̲���������ٟ]�6 V$S�pE.yG���K2�)>'T�>V��9a�e���!�ִW�k{y*U�V��;,���L�Y��o�~���@u�R'���MB ��.���Ֆ��N�+ a�H7gڞX��NZ���y��w�/���m��
��M�1n��yj�4�B;���� ��=�7>���i�A4){֦���+�'jp����N��?�(`@�-��Q��,��R�$1�+����y�P�a �/�Y����Ι��!D����ɖ��ـ�z_Z�<����v���2���e��`{�qY�@֐>qkU�zJ�������/���^���Gđ����
�9C#ofZ^gT�Q�A�(��f�P��>X��S�����/� ��'�M�������������>�Y��J��Z5����5��b�PQ����h����Y������M�8�� L����P��n����H�،�P�B/�3>�w��%��᚝�@y� 2��;
z�yJ{%�s�d�'��F�3B�V,!CN�hAA�,��������	���e$�ѤFDߎ�ҳU?M�Zr�s�ˬE�v�tt�����a�9U-*�o{���3��D׃� 1�^�����R�q����'�Γ����U\H�b��4����7b�0.=�[?R�TG��mHN�Uҭ U����dM�qW{1>|'<|��K/����,P�;'PN �A?CZ�!#�k"^���DIX�}�$�����m?W����|y!��f�x��:賂��_��D
��7�Z]�'X���Jue ��~�� �D)��ɲ�Y7�=��9!x���^l ���卨�Y��*(b�o����o�Px�+�G	��#���ɬY�ƹib��XQ��zΊ��Y ����8M��3�_���B��d�.��F$�-n�7
O��Sc/�fIz�D`��#���0=p	)q������W>�^ �͵��v�n(�E�2���ݚ1�į:���ßD�]G٦1��<B6�蠔֓�E���Y�
�,��-� Aӝ�E���'�"��Y[k���y�|R]-6��u��[@j�&C��l��M���Z ]��f?���������V,�Η�=!E���cU\���8���w�V����{"�³C�헍Ae4:j6?l�'���M# �� k~a��@���?�gg凌�}��צ(ym�&H�B����,������ ��Y�~�l�J)/� �=�G�̈́�a�E�N0SXY�fnE�½>�*�j�l���n�zfs�b ��<$�Q�+�������6��D�T�aMZR��K��Q^#Ca�^�Ou[�g����S���ä~?Z��C5�+��c5���H�B���жl��E�Pf���#�$$��*_����ZZx�<�G!�X	A��uqj���Ȝ���D����H���ܮ�MG�6�P^����7Yͦ3�ԟV��xĂw0��p@��9_�y�2�#���: j�4G�kqv�6���LB���>�e!�����.V�#�:�M��x�֢G���� 9\n����1�g�,((k�	�˕���F��p�w�8+ _"�K�9�,ܙs��@�M�(YqV:FJ�M�'ӕ�t� ����M!i��Pz
&;c5�s�ٍͮo���y��������納�O_�0&E[뫋o|�]�	�O�4 9��=QԱWw�B��#�gfZ�e�c�Ν���I��g̅�I-�u���Ě�QZK�*�S������y"����	(����M�^ȭF�8��f��Z�z���-vĪ�q�X�R}ć���)���}0L�����{��ghقT����=�M<V�w�f޴�r�y�WIx��)�z*��,��������W�Q-��8�ퟯ���a���>��<%?4~�O�_���S!GRh�p�yhf�fF�� h�����~R����M��Kc}Y^�ʐ+�uU�43��Vݮ��
�v�>��� u����	��qa�5��d���&4i�O�����t�
�� :�u���!��N)�����N� oր��CՕ�ۇ����P��U���=����(�g�BcT�S��,������;�����=�]�9L�1�w�_T��*�X��g�Hk9�ηI�jpW)z �
[˲�-l����^+6RD�ƙ�!�wB��p���� ���6\N�eΝ�Y�Էo\_��CM&ނ|�7�i?��x�B�h��ZPPu^�����yą�`�)b���C��*#(�jP� ��6U�Ϡ!�0�_$9΄^��ϥ�< ~��M�۰����� ~鍃��ZI1&�1d�ϫ��S �k�W�բkmx������"�۩���BFb,H��^��K(8�sg/l��ܽ�D8v���MLto�s��Ms�_7]�dN�i�㾟�P{�a�w�H�(^�Un"�R1��V��19�(�O���a؀�����i�6�� ���nW�&0vK'dP�k�~a��>�]ʎ���tP@�a��4�HčųF�����\��Z��G�z��ΙK�����G��sY�Q����[�_/�I�|������/�c���3�� Y���8����F���A�B��bvnP�$��x�ы��؂��}VdE�W��w�ä�W���(%T�b,��a g��1⿃}-�ޟ�mq�yo�y�Hۻ;�����Z�@�: �nF:8Q�Pɩe�t���8 d�\��cD2�qV���,s[7��0i��w�Ql��D�.��t<���� ApL���^W��nBU�]�E�;�^�{ !_�pH� ����J�����^�}z����!06��u��c�"��;�$X)�h��&�I3���e����H7�w4�u�[��`�g�A�6���c'���,�R}4��!���2�2�c�����4�k���p��.���
�B���f��"l��Z�f����\�O�N�!L�v#���!Kε�q��٥��yb�(����(a(&�#y�n�9�����_�S�V��5-Z`�^��t�F�$�@l����'���Qkrި����3p���9�̪sϹ�6v�����)]^��&�9��#§��Ɣc�	��*+�	���Wƭ�/�2��0���Ҧ[}��&��O��,�N�bHZ%��!��<�n�]�����yK��.��/��8l&-��O�iW��l�f�vYQZ�wl�@��3���Q��AI�ݟ%�/��
��,����K��A��n�X)��=R�l�^�#EV=�T�������9�_����U��lT���Jp2�
[Y���oA�τ���>�d��|����n��M�dD�&�B�(���Q�f�q���:���+�|���<��E�wi���2�`�:�>ڭ��]�59�#�U��34�)�V�5��5��Xt���1�X1�0�<��Ǵ��)��)pM�{@��
4"b�E����V��y�����> ��/��A�пx���5Ŏ�B|��)��)��V:@�;��#��+�O�_%������l�0�yP� �s���wF9����=~ %�a�Ƞh��`ɕ��)���6
$�͚�Md����ETQwg5��з�j|i!�`yp��b� �������K�F�Ss�!$s��˹�_��Zm���w\1�gzVM�1n$hs��]�e2Nތz�Er�8~مӴ�e��㗱j�gi���j�TN�=IR}���<��d�ϡU�n�Ec��u�G�K=��[��)�L�G�-*Ξp��nG�a7�f�e��t���hi�P"�TA�c��]�O�;�f��?��l1�:�ǫ�v��a��uW m]��t�X�WO�u.��i�,��� ���})ǜ,-�:^?�������Z�����j����K�sm�Vf����Ūw5���,�����vO�SQFrjs��U���ADLC>�Ņ�I�� H��<���e��@��F���0k������?�Fr���O�>�P=����ߦu��w�r�,�ʷX���MGQ�ҷ�_Z0���G=JO˓�V	B��l#�QE0,a��BƓ&��9���6��vZ&A�0���FթZ�'Jrj'.�8�F�pL�5վ��]g�ϰ�9���P��4r���ǉ����
D]�}_U��,��[�2Z$�˩��7�NraO�e�a��6*h�~�	2��EL��JK
�IެG��n�/w�y~V���9��"�����0�p��/_�\���p$�]�T�������_ukн�q�]I�l�l��/��[�50��3~4�5�Cer�CA�,���&ʈ��
r�j1b0�3��G]�[��A�os�CJ\�,�Nj�l����`��wu��KG�s�'i �U HW����I��ڐ����*�%��q ȇam��1V���qe׋θT�o�D,�c�x�X3z�!��K���:H���N�=$i���^�5f�ex���N������O�X�;(�ž���iY���N����u{�Z��&�`�2��R(3�q��Gr�D�N�o�cbp�*i��a�#�o�S�Hu�4�;v{�Ca8C?����}��t��~�:�K��K������ck9Je���:N�i�cߑ
�m����ұ��I� ���F4�9u�Ze�Lc�Ptm��k�M��$)A�NI��eT��ϒ�[��qFIC��M��o�3����	����`$�r`0J�9]ѱ�� ����B�����]h���U$��߶A��;��iԇ� ��p��2�}BQ�'B�S�NG^��|�w��x�e��E��~Kdk�Y����%�-�Ý�º���f�ł���
w���2�����D�옧ݣ��d�5��������˅B'6�a(�U���-'��B�vb����m����f����ύ���0������A咽�#�.�'�NՏ?�@)���L<wS��rl���P�OZ�(��� ��pl:�CE���`��
�e�M��k�9+��P�C��M
��j��U�+e�<��9���~ �ȷ^-���z����>˅���.9UK�}Ŷ2�X�|��[w~�2��Y��`��ޯ'	� [�v��lH�e|�
¾���"qF&(i��^?\�;q6�Ν
�,�!�F��Vn�-8^��x@:�a�x���j�k<�nLf��i��sE�p�/a�kޡސ1(dT��v� �n�����o�a	�������=��^�����7.��Q�����~���ne��G#����)u �
���GT��� �a�̕�jh�eJ?����{�V��P~!�6�W𳐀�}�5M���^����*&XW���|ʩ!�6J�����u�g��'�9��ҷ�I�u@í��V�p`#����������ې�n���p�!�*Cq��kw��Pu��N2�(�a�RK8�f��vq%[�u@~�Mص QW����˙��oe�ݰ�����$'�9>AD��Z���dT�f.j��4����4&�I�:��-B\�R0Q"��*�G��ā�2nD"TE
�z�&��LK�2�r|۷��Ťc7���N�l����I��,۩x=�W�Y�<eOX�c��t���&��W��'	�L�m��S��5ړ4(�*�0��g��7�u��h�}=S��2Ǌ �i�+��<�0���L�Ye3�rp�����]�1���Q�$�V�6�%߫+�GD^de�X)1UI��2��g{�)��۶���h�̶`}Et$˺���I�P
M���r�OQL(�3E�����sk�r���i?kq[�x��Ns�Gkm۔8�D� r�Y����T�Hl,��
�8߿iq1R	����m@X45�~��-�Iɢ��c��P~/?8��L���Bd��N���kG7U�-r���^$mPԼ��4��E�șR9�> �qr_��Qٕj�a���;Y�߃��]rV`25\�i�$��P_2C�t�?k�=Ӆ�������`��?	�_�B���w+��<m2�{�۠���]����A]?hv��3B�U)u�Z���?�,X������Z'��HMQ!���r���7@ni�*h�V�w�h���+�Lq�/�	�z��8!x��C�HT7 ʣ�14E�d+d �Ĕ��m���L~[i�<�v{} ��겟
Xw� �+Oc
i��.��tV��d:�8�B"l^:ݐ<�sS��q�x�����d�r��h�`��sw2����ۑ"#/��p�o7 ���	E{��A��M�֎ڏV��x�P�O��e6ҙ{��vc.õ7G���E@`��Ê�L-Gq{,��Q�/Z\3' O���j���] 2@U��A������jt�@<�}�.�
�6X�~�g̛����k���75�Q%T¯tp�`�|�ߐ)�-����N8��Mw�(ۀ�*� �;kmy\\u�rm�CI3n��jTvf����N�G#�@0��2č?ʁρ3_Cn	�fw��9���4�;>�R�s��o��9�)z3
�J����x�r�8?$4���\"��a�FG�����IDgd3!���ַ:ԋ -�{�j�KX���y��|���Q���a�/ʦ�mc��M�1��@3Qh�ᾅ����9�L�ݧԠ��K�a˕b��z������v��x��V���%�o�е�ڔ�o�N��ҧF����w\�U�,y���%������8Wt�<�3���E�{�#���bj<v/@h˖�I/b��<��rJW
�>�/���uT/�w��24�fkjF]g���ڟ��C��KT�����%� 9����ja�w��Ӛ�NF�(�o� KWpε�U*���J�TLt���	2Ѫ��E�����ᵉEU�!Q0Z�m�.����b���P�����oc����-e�ʷ7�OM-+9��4�HE$Y���$.բ(C���\��H�ZQaC��H�`�ߓ�@S�Vsh	�q�}�c2���Ñ�G�U�x��5����S���Fyg�6�B}���*�Ɇ���k����i�d��K�L����fqL5,Yq�Gq������R����s���I���xlg]g�4�ʑ���fA�^~\f<33I��MeA��+�ΊՊ�a�RǨ4�P�tZ��0
�u���ђ�3�#��f9Э0���	�Ɋ��<me��!�ӈ9�q���R��c��^����L[|��z�w�
�52GI _�#Gw�� [�4�F��#��,�EVʣuw\����>��6}Tb��K(��k�9e�@�!.�FeƇO}.]b��J���Cc���I`���q��IS����5`6J�����k:�?�x�>�so	4�q/����3F���}V.h)�	/�-N� n��+nhr/=%2c��Ѿ
p�O�@��%�.���{:�b�tI��4������Qd
�Q��=���`� ��t��~���v��}F�S�	Vw�h&�\r�D~��c�`O
7����h=��,Q�9�_捆��`�b�D���a4uy��1���I?L�#(��<�c���A�	�LF��Tdbԧd��#��O��D�RQw��j�sl�<N�{ ۨS1�W݊B���NP��0���i<p�wM8b�9�ğ,�j�Q���".�uoh��\G�a>D^8�հ��蜉������k4��l~��y>v���Q�F$+�"���'т��k{n�NU"͏C������PaC�N��1@�O8�aEri?X�e��kc��@o&�fO�l=���@�P�,��ߎ�x�����ću5�J��q����:�����dLo>w]����y����^����I�C���f������얽��2@�	������Μu8��鲞�2/*+����m�&'?KW�j��:�����Y�75}�S�z[�����\�G�m	�� B?{�E|Cj���,{c�w�x[暧P������nnW.�����,�s9q�b�=j�r����D�2��D��襐��`f�D�(�hΖ�9��<�!�w'I���]S��L8GL�`�qd� -��A8M	����!M�+]��^������b; ����}�ܓ<;ݭ������.��7c/jf���T�zo�'y !�Q��]�c�k���o1��Uݸ��)X�ٕ�g�rR����.��3m>!YP�W8m�3�)����%��K6��P2c����xq��F_�)�	`���\�η/���.}�2*V�KԐhks�m����.�U?�m��#ح���4��Iz�f𩾜c����=?Η(:����T�ya�I��,�7��Ԍ�sM �t�Z���t�3����!�B�2�ʘЅ�̆��K�]%]�J��]�����Mu̍_���m�k����s^2yr���d�Z(L$�)9n"ص4ƽ�^���a�~V��)�<%A��)���C!�R� -V:i�5;Vpz@ҝ�[ҠXT-Z� �u ��zL��7b�N�E�R�$@���W;��"X5�ڣ-ȭ��������`9����Ԣֻ�Y���f'��]��`��n���'Fu]r���w��q��Yp� f���wa`n`�5��q��ք�_��n��Xf�َ��y�8�*wQ4��+l����Q-d�Bk�U�k����Ðx}��3pV?�<R���V����|n�2@5�s䛅���C���zf���ޅ(6+�B� L]�RrS����r۸�PʬT����u��~�e����}�W��㤖��1�8�m0����1���04�T1�{�3�P�		wg|�:�8�Ά7?�@0 o%Ѓ#�.���`�2|bN��y%�zeŇ}Dq�����)�1(B��M��?��mW�G��_|J�j/���<u�����{���!�j�[ۥ� ��5iE�6Hc��!��.�4���`�tX��<O�x���V���i� �������F(=	��xf�n���~��Ƃ?�uA�~7K>��D����)@Q�9�BN�!i΄5>�3D�?r����q�T6��K���Xݪ0�ݤ�����J\���]�NV�G��U�VH7�u�:��o�ܿ:,[��9}[j�L�s_hP0|�A���?T��dpg{F��_L&���٤"fa"���7������gW�nZaBQ���w�]׃�z[w�	3��D�^�v��������kn�g·����q�"0C�O�j���?�Ik`�_��L�[ӉҿmW@ 	�N���Y�,�xk=s�c�$�
���6(q;��)2��[g`���o��-���+GyJ����������5�a~����f:��b�:Ѻ��&F��4{�8>���������%�O�ӣ�~���}���YW�%M]�GH���N���kq��O���S�R+M�}��}�܉��t����.�Ob���>��č+M���L���@5��t0㻡�
�{Y^�6���+��*{����W����n�V?�tҷ����)��(�&d3�D����5�i�2�DԂ��P��?J	������J����&��ث<'�f^��]v���窅t_��c?�x;r5���
L��Xm[�n�8c����������n��Z�TD}]'t�}��6�)w3�uS�0�է)�,���0hX&'k��	;����f>���Ԓr1�=��v�Pk}|��Kt?�НF�d�{�ہ���e�:F��.Զ�|�#��p9bzw<�xd5��	%��!c9=�6Y�k���3���X�����[`��p33�3�U����?)d3�O�������=�8ݡ��}=#N��˿��R'V�;u�"!�6�����y����(�*&3��9CB;|�4ܠ]��34�Ԇ�p_X�
i=�	�������k#I��{X����Y����d�v/������Cݦk�ܿ��fש_���1���͏B��%b?���6�(C�����bu��Ot�O@uO�R�Ӆ֝k�0D�rW�1F�����vx��/
�5\���~\�����b�*��N��Z�P�Ν��/&�<�wm6O��0�>�Ai �y��[�"����#��f��)�ӎ}+��X�&(a�p,2*�S�y�/Nm �
Ӂ���F����t��0�+m�&u��h�Ō�6֥K7X��{;`�֋�@�|X����u�\O�pm��қW�t4&D�P���C0�6��?}v��6��G�@q�Y��1%���;�@���W1-o���h3T夐������[m�'����.�z����G�v]Y�9�(P���p�<�ʒ��>Sj�<6����
������#���!,�N�z�r����}���@���y꼚��ц���~;�g�kLvV��Ov�i�^��Ǚ��zY��A!���bp����x�c;olz�`/���d:���� ������C6$�Pc�z��󝈣�N&����'t^��A`��r���=�~$�X>Ʋ5O��K�$Ns!�@�y���0m	�� v�W�*nӷ��Y�3>��Uظ'H}����P�`KfF~�8�{9r�F�f�+�e�,I2�.�SB��#Xn��$zE��EVS��̉6��8JM�T�H}tSE�PD�=6E]m+�٪�ۻ����$��av��wM�H�Qz��Z4�|��5�|��7��e{֓������%�����xW]�3A+`�q^��?-��SY��?��\>[��������6F_*�W�+�ز�%D3�#9D�c��Y;��d1a�S�6����rg}��F�˘��7o&�z��L,;]���p��czMWS�ͧU3/I�(��	��y��i^��l�}O#��0�y��d�JE&�ʷ�>�$�NB������ի���g��n ��V\^%�ש