��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�'�+2�HZl��̜� +a`ۤ �^P����*X�d��{�����.d�}���r3��_~�M���7[6�W�}�2��Z��w��Ww�PWCS�1���+�ܙ�Q�EN:5�#���w>yX�D�x��P{h�_O���ml,.�P�'�����*T1+��W��)K�YY�u���$�h�Y/ ��o�b:�W���e�T++�%�t�FX��iqu��,��t`����m�a��6�e�vx�+��P_G8;�eE$׏��:J٤���]	����2U	���z�q‎]���̄�_���CG}wc�IJs[�2e��01�̿�<�k�t�jՈա�r�F���{Mi��M��u�m�,LǄa*�����bVQ����Y��s�N�!ɺR�.{�P2��+��T���5,��߈w%�� �:�x� iW�`kȒ�t��vwCU��um�ֹv(L&�I[��U�Ap��{�T����'E3�܀�hʮ�d���Y�6�������}��ͩ�l����p��h�'�Ú�Wcn�=�X��sG��[�b@���.�7
i��9��f3I/ߕ���?�����~ߧ����\�.WW�,����H�퓈�z��`�Z4�d�P�0?����uc�P���30PPz�<6��<4�����S�����v-W��������1��ˡ�i�K�3��q!k�[��)���N�T+��6�)v��#7��#'B͎C�h1�v��������I���a(�	x�f]�t�R�-B	-o�.���i��������]~'_�����~�xܩ�j����0z`W1��g6��X@�nz�4d��r�P�Z��M���.�}n���=�Y�> �w^�A�J"P�@/�o�2DJ���&:��2��4؈�N�q�M�_�+*_�h��>�r����C�w9����%�Ƶ8T�V��"R��!'
	�(��?R���Xe�$�f{�Ԑ��0p*��Q���-c�~fW@Z\�����C���(#;�Ak�YF�=q�'n��*+�xb,� v+#����S�2o�H��t�0\��1z)٤O�mI��Ζb1��u�m��Y � iAng�Ys��Ȳ�b�SG�ґ�+�C�X��v� @R%8��b#;^����1z!�4��d;�!�c�������� �m8V:w�=ʭ�=�b�C�^�0^7Y����yY�~��Џ�I��+=`���,z�^TA߱�T�eCaK�!Y�<��Nl��/j���?Z��ҙ6�-o�����c�rK�0��Fxs�G�9��$f%�<�#/��Iv/�`�B�u���p�0ӽv�v�n:Y!���+C_�r�%�(���%�0�&�|1*@m��wq�K��u�_,�@����� W�����oe�9��=T�a腵}�])}A��'צU١e,�B/��W+���ϻ��3B���;.��zS�:��ф[���
%D��n��@+�ꬅ�F�H��6�����Q�?Ӟ�$(e|nZ���l��)Jm��sF{�)k�Mr�>rv8{.=1������[7����$��U2;���+`hnV��l
��ecG5a�h{�� �?��R�R�;�Wjr۝�Јq��+��/�����⸉b���<X��7�Y�#���{掀�C@���rͭr
Mn���h뾛	bs��rР�ܱM�&JN>��Oba��j+V���N��Al`�U>������Ҋ�ǁ���<q��߇�>���7͛u���.'i����s���Yus16�����b��E�H!r;����pw_K�A��������d-�U��3Dzeq�s'X�m�S����e���	=CĜ\zJꃆጃ���<��
��v1��4�
�y���2$��#���y2:J��Jb�?��6\��e�M1��Oz���O�u�K�@Uyr���ߘ����%��MY�c�7�mDtߛ]#C�w����\{Ӿ�3���t�|�f��� e�V�e�К�L��� ���Ʊp~��bk�8cN#]jv&�4e+��G��%X����բ�@�5c�[��_�B?w_0�LSp���ЅQ�X� `r.`9{\��؟��JŘ�`��w�,5�1h=P���T�_�5�^���{�Fr�9g�=[�[�x&�"�p[���om8rv6��5�J82
����o$�wWZ�o��D�����-=�;��'3�/@�:����� ��;�o�Я2���)~��yz~�pP��n�s'�����}O�O��MH��y��9���#��ϻ2�9<�N�U�?��&h���Y���.ɬ,$��!��P ��	Ռ���:����7	�8č8�^�^�N�f�Y͐������`�Xn��)8�Ex]+q�A��՛}��c�@��w�����i|w��@�wd�,~�TZPr���[y0��m���J�$���s��d������D�-&�$VTh��P͖�r�:C�-�;s(�J5C�8�N��ig
jE��Cqo�=����Ni������{�<���g��[O�"VR�簠�}�m�%��G!���0Z���N�z���;:b�C�"PT���蓭]m�K�EY{=k8���w�;?���8�T6w����'2��h P ����X�"�qQ,�GU�筘������Xf�K`�b��?�/d�M�_-D�ɽ��E�.��_�@$@ǉkm9'���_Tn7u����������z�z�Ze?��n7��X�(~�J�ua4]�8I�?bV,�S�U�^�&aʰ�57���i�2(1���7f'p�o>t��.��0ӌU�)�����:��Cg�'=�$��O�i�i�zVѢ��].��A�qt��s�9(3�p�#+?|��Qw�%����ȿ�aC����i����A7�$�-��+S���G�`+��P��؉ ���|��p��:a� �%1o���A���#�Ҋ�Q4Pk�+ɚ��?6�P��B�kڕ�r/�~��?����n���Y���HꐳX�Wtle�M%,'o��¼���3�u���ǽcĠ l�-�*�f���l�4)�V�!� ��W��R��˯a����X[�
>�ٴ�y�o�Ç�rf�YQ��)K���>�b��J�ÿ�O���YKw�_����ϵ�����R13Bx+m	��9�ya���,P�ӽ}�[�bt�4_�Z��p_��P����+G^�j�Zc�ß�@59l��AV=�n����z�r��%�UO3�r%�Ҹ�w�Ҵ�a���GQfT���27"�v�|���pg᯿��9#m�S/�l��Qz�E�[�t �4����.6�,Y��Q��Ra�����U����V]�;���un=��g�acF79�M��j-��:�!i�/Z��i3
���;������S���,G�����C�h�B���*����k���35i��<sp(,����i�0�1���r�?}OH��t�����_�5�W.������z��)q<���?F��=�Z@*��4�5�Iw9T�O����a�.���T+]Q��S�K�ԏ�%V�{��'��[�iv����j����Ħ�N4�E��K#��Q��Z�,a��Eԛ"��Sz"�C���K��*1��� 2J[?��P�g���L���$C���8!����4B��~dN�+V� �g�L�A3w�hoLM��X�.��&O(\�s`Ӊy����f�����~RI�O�G�ǾJ�����7�;����ߎvG�j�jf~4���F�
M^��D���m��*"�b�7���a�q��7�+�NWeTM��.��γCn���|3#���+��z��Ɋ���eh`/�F�0 �ѓ�F~�>N��$i+k��)���EX�=y�nknh����縉��g�8U�(N����)�@�Rn��A����1&T����H(tߕG_ja+xǤ�_Ļ�bt��{LS2��,�;0��|2���eF
�lΈ�p�'Us��l5��O����Ǟ��6��=�=��M����ꃻcPQc3H|~�{X�� �ƥ�(pձoX�߱�����a�=��-J�q�&v�E��7*`�^@Ҏ�r-
;��sS����[���$�	C���tVi��oz�a<��F_��֓�ɭGf�5���Cd�����?�/K<�q���C%�2?�.�����;���u52N�
��hcI~�����ju��i�������8ZK!�x����L1J�kU�(s���h�u��Ѭj����Х�����bO�1w�w0��eu�`R���<��%YXk���)�1���L9۶p'��K=m"oƦ�2�cgiV�{c-�\�,)Tf�U�:��H�Ь��d�	�V�j6M��C��8ފ��w2�;ҭ}h�_U�>���	U�Ю�-�Z�X�>����A��/�z�T�&�A�.a�Mh ��鼧��+3 �l}�� ��eK��\{�M��L���n����t�݄��H���7,�[�s�([�`8M�`��%n���&�h�a�0�o�8�2��3�����#>˾x��cb����)��\͑I|�P"H�_(S�yk������?��B�#�ےW���������a}����`'�;#�6yFץZ)��cyj�m�~;',�ca��R��MY�]��/��|}GИm���F�M�i����h�މ��^����]���esr�j�u�Wy�٫ćTǃh���יA��T��dǕpu8���00��JW�3�y�:f@7��a���ܴT7�~�+h���n�mn�
�CJ�F�k����eA5���no�4�,�'��+��T-�5�|�E�Z��K�*h����F.��j���O�,�1ZNI'�D��*��������Bd�c����,I ���
��I�ꟺ
/�L�k6X�س|����t�V��ܘ���6��;f��
@�vB����h/��MU>�Q�֫�}����of�g�Y�mZ�u�+&����4�1a$�G�3�A6^)9N��g��O�7��g��W���ʗ������-^9��Zf��S0cU)Ѻ��8��P��;H���I+$�Z)p�ͺ�����Z��;���=�:��:I�}B\^Ê�f�_ƽ�@�KR�#A 8�����u.����C���ϐrH1�[��� ��m4�)�!�n9�V��Mv�-��	��(��OMC�N1d%S�Q��U��o��D���*�;  ���{��!����^���N��GYbB�"�U��U�����=�jy���(;�o�➲(���������0�V�@��Z�:��0��a1˼�ڶ��c*�{��S%�W��_���YQG�;8���90���;�J�����-Z}�����ѾX3�A<��F"�<loL~�_?�d��,���_+j�՘��+��ʹ�&ftvԞz�_�Cd���UA�t���j*^lQ/��*L/���.�Srb��n�:OD��{+c�����!�/@�h�]	��Jӽ���'RJƦA�n�f��ytqQ�E��`'A���(g��W>au��$R�,��@��<}��%>�Mw�'����jآ�e�i��;h�kU�׀�]�?
�r�l�W\4�u���Z�:����>�����D�����]�8G�Mu���e+�y��1͵�Hx�,��
��d��i�OŴ����7�����n�:�E���.������2��(� i�qi"����_��Ω�V�`�42^A�-�Y.-/��Y��c�S��j��ԓX�˛���#m�9�q�Wj�旕�a&����?6�z\t�1��¸"�����&��^{d�\�JfbN���C/g���a�7S�y|(�����_�r{�^�+U=(�����9�L�ּٙ�c��Ƽի��@�
���^���,ÛE�w�����䝞�\#�	�`N����"%y�+���M�
!�-x՘�$E�Z,������D����3�	��i�+���w.d�7>c���u��؇�[��A�]�A8��"�8}�0}��&eT�}Xr4Z��`���(�9��*����c@�P<�Na�����H�U��P�1�/Ƨ+uK�/�ڼw]~@`�)$�� �0�M.F
9�GD&ɺ�w�τm�gO��NI;ω�=��/ X��h8�*�H*^
��P���x����(���>ޛ��:C[��+���E�y&��}��z���[���pwc����&74];���qh��LMu|�o�Y3D�xeu2ƫ�m�k!��ql8i|��D�HU��}��S����Н�]�JO����܃v㮶��~�����P�v? �)R�qUNQRM���6���|��g��Q�c�2(+�q�8��5�C��&�. ����2����	���+<|�\  $�r���9��2�����@��w���c�v�01��p%Kr�y�ξ	���u�?m�l��(_*\Zv�0��?ծ��t-��R���h=B���KrW6{_2��CxؠnR�����������~�x��������A`v�\[$cqs���Dlx��x���&5����OUN�m��\^~w(�S��-Û�&f�rI����ٓ�3�YL���̫�F�o�z�����L���ʌN����ۧ��f2}Ì	�����Udô"Ͻ	��e�~jf/1X�:)k����4p`UkΕ*�����R���}�٧�yPd�<Z��}��d}����(?3f��tN>�a�d�uޚ���5!l�D��/]�4� �$w&��9R������U!?M����6�&[.=fM&i20��kR�@�xg��=�Ó�p�h�#܂|C��u��ί�o�w���[���0��>�_�SL�kU���N��F.��?��gu�'+n�8��9�����P���vřs��"z���׶?IU��U�(��e��nڿy�ޗq5��X���(e$vtF�� PD��G��
#�v>�U�à��(���0I�_��a�n~Q�`�BJS�˲�>�	��h�]���*�_�t�[���}-(-V��8aq��u�5�x{V˥۷"�~����K�6��O5�s���!�kyI-�Fl�h8����q`�y~['�Įt��OuHh����7���S�����<��1.��Q@s��N���P��bm���O5���%�4���d��u}M���"o&+
@���a>��ɣ�~X��?�9�rE΢Ʃ{yd;�2˯��!苓Y��F�$�-sp)�@N$vU���R�0h�a-x�~߉���E�KX,�Υ[ި-%�GJ�����~�O�G��P]�0�Wm��|�3����_�#x:c�5�9���ׅ�o(�u�2���`swc�AT9��N�����a��yɰ�a=�`z���j��6H�@��c�,��u�T(v7"2�͊�ZNF��U��#l+S�S��	����8Li�9�2���\s�`oȭI6�r_��z���ql�	w��c����AIV"��A��Սc��%X��RG �����X��l������Zu��5�B'��~6s��=[���)p$�=���M91�X����Ѣ�a���jtH@��(��uNб��@�W�\�"�}����t���jC�s#_�5�w��7�VEOi,BIUL/�w&]��G�K��t]N�¹la���`�I�H�QHHÉ�=D�9���1�d�Eo�6�΁�M>��S:�"o���e�'~$b��_U4�9x$�G�\���;�����h���Yy��R*r�5��S�������V��G�ݎ�~�N`B�V5\��N�����(/�k�j�𨡥1��}�ԇ�;W02�Կ�y�o}e��?Z��Q��@�ɶdF��F�v��"R �W a0���![q>t�G�{-dW�:}TK��V���ҭ7��8]_׳��
/���a-����B�*d�����(f<X��[�E&h��H�$F�������R���,�0��08�������������ӗwfBVR��v�BК_ �iu��lA��UZM�>�lc�ki?�S�:)�7U��wɒ& ��{-�eq����^iG�*�".������0�����tL��{)w��@�����D��؉��b���>�;X@��%_q{��R �N ��;����@[���0��!还ICjnz4ġ0(1�S�(����z����k@��y��&������S�<{`������c�$��΢�Lv�G�ł�;��3���%���=*n�̀6l���p��9����"�q��6̺�o�dgl �{QǶ�=?�B����{ÿu5��4�d�h晇(>А�>��;�'�l ��:�:��_��ל#c�zmjH� Ъ���zO�ē[v�C����DJ�yN���!���/�z�N� ��7������� ����?L�-�z�F>ﹴ�R8�ęh&��X3��1��SXi���!���G�M��p�� ^�HnKZ��JL2�r�ߐʌ*�[gn��~p�F���T�.Z�1>k����宻��a֗��#z�1d�Zm,��+�O3�v�����`qu��[��_M��sAw��s;w�^�s��g ܯ���B��0��%E�0R�=W����"Y:=�*!�a�[�����jN{_��0��8`R���R�Rd���vsg��8��V��GG0.� c'�f�KP�4�a����$a�ϒ~��eF6T� ;�S��O���}�v���%���',��6��t���v'i���<R��J��2�2��y����h�ꗓ:Dՠ�u%5���������SG�iTP�>�?�N.c��5 ��J|��"�}��
����]�r����m�7N
�o�����"����n�u��.���O��1+Jy��Mc�?ݡ`��O����)=�n0�C�U@o�Ƈ:�7�㉈��漛EN�Y���|�Y�֔9d��$���|�|bKW���1}�#�Ƣ���Tl=#y�S�(3J��	�'���=������J�8i�-�ظl��Ρz%{6����d��=�$BIHwĺJ�NU��dޯD�X��bb�]��+'�~�h�5w���\&��(w��3 �>��v���*�Z�P�U/�yyt+��oq0���񂎮m�4�B�ͼ��Y���p�x�,Ɲ��wH�w�o&�Z��C�'����J /8r-m
5^��ʆ�_�S3�ŝ�m�!�π��L���c��jD�n�5�x�xI�'�����l�U��c�M�n�_��_�]�'�q����|�������:#3q|U�A�&�?�oM��Yϼ�~�s!Aώ�9�cP#wEo�Sn�f��zW�<S�u�+-;/�D2��a̰"Y�6��<���'��+˳7^�&�G�U=�KAU��P��D�D�<3Ut1�:��M3A��s�}�;|��l�����,�4�9;�f��}�y~�U�9T���a�C7�M�%	3���39X)uA�Sf�J֝0�Y*���饂��r� �y��5G�ظY�MȽ0��D�Qg�C,9j��	XToN��:*�kR?�v�ϔ�U��D-����~�q�傰�'Ot%8w��#Q،�<��n��:�6��c2f���ZBb�M�Y��B�Z�M���Y)�����wZ�G[[l��p���B��Jdt(�01�d+�8}`o�_��A��b_����ZR��?�b��=��'ep��a��"C{�_=/��k/��e� ��>y�8`��O<)�+~3���T���,��"�(��`V����魃9����v��oς/];����xoj6,����]~��tU�y��_l�޻gt��N{���od�����d��1Ј\�� �S-�H�G=�\���o��|fI=�j����4�-��9}2�����1sˏ
���ͧ������1>�NН��nf�c�QS�&��#���eކ�/zZ�k|�k�|^dgN��H��f�#\<�s�c I�w�Bm���L�ڽ��n%h#�ಔy׀�&!u�4w��������_��T;�?:y�"��,`*�1[,�'3����0Pz2��޵t�q1e��P�#�DZI �k�M�t��<5P��D]��G���`hs�JXc�������h���C��1��Ȟ@I�(�T��D2�����x��z+���uB�vN&�`���[��bp
�Ci���%��C({)�U�/�g��������ۈ�m�;�ҵ���D��]/����I*������u�H-�.*��h����)�%�p���l�+=害������iȢ�Xy�c�6Au�tV� ��Fu��$�q����'(L���諔�ʄ�+�b� V�/v� �(ԛ�fw��el�ZP
�b茮�\A��Hk.z5��˒�K*H����y���j�0�P��Q����$���^���l|��P�**av	d���V"6v�8�A-h�H��a:�Z�K�
�Y����h�������T��Y
�@��:����m��2}Nז���R��~��|�zqT�N�Պ�+9��P���<������3����g�2�3У�&�eQ��@�8	���D�ە^�����}����ƒ-��y�LmQQh�	��^݌}R�d{��1Q�fT���OTE0��/��E�\�m��^w�4l�m��W1ϡ�{��L��xl}�!
��7-�-�������.��F����N$���HJ�A���,�l���C�V��؀!��Zέ��6v������t��I1:e���J�S�{y��۴��`�g�J=N��HeP>C`�)a�d,/E
ͦ�Ȃ����3O�tc墆 �.���l�6��{��,`�w��܏.j��O�Hid�p7uqF�V��UK���k<L����[�&�˂�%�E��^�s��/��f+$�zJ�R��c!S�$N�Nm|��֩��kuq�k����@���s钨���׏�e��̫;��U�G[K���0�S��Ȫ��hCD*\ ����ڝ%褧	C5�0ݝ�Y{b�ȸ�i�)�Qa4 }�Jj���YV�b��o�+�GҜ�'���f����F2a��85t0��~"�R�f����gw��uTC�q.%�1�3�n�d��>����d�@�~
��w3x$(�SL�Pc�JX�:d��=���QEWyε�µ�+�{���.�tE]��]T��2��aZj���7V9�l��+K2��"	������3~��C0-P��mė�pU'�UY��rG�2�ۅ��;Igs\��%s���X�O��^����X��5�K��'�柊�2F6������空d¸���ˉ\���\��V�K��8�h���x�8�m�R��)��đ�s(QVd��n9����0��}���i�l�K�;�R<<��=<���=��%�e�����+z����� q\���C���Y/(�-�蜠t$đ	n����86�G�9k6c���Pɤ�޷Y�N2�1�Vm/3β{�����o��=$K�y��͆k�MW�~\����DU�򭫻ͧ%��5�)�Ġ[��k���r��قT��[�m��dU�d�3�Ν9��� x�u�:�,������*s�Uw̄m�b{!ҷ~�R��pSR
-��KĲ���x��%����VZ�Ζ����Ř����ʍ(������[��[�D?���X7�9�&�mŝ��/�|�¨Ka,GG��Q��H�M�3��5��tY���G�'����0Q���W�1c�����e�e���sIQ���C	�)�Q[���K�6@2��U��N��Ή���C�� H$ȍ� �t���vd����{��ҷsL�EB)�C�J�\G(��DTly����#I�e��r�()UYf���}H�bh�,���0ŏ�0��_6&��2���m��Ժx5{'��c�Mv���!h-C� �:$IB䠼����cF¶�i�nZÖ���]�tҠv�>5��$�.�q3����`�fl󪁪hH^*w��"�����&���D�C���|� �z��R�ոs�x��Ŀ$�> �,�_�I#�=]�y�A����(V"��	��D�n��v��z.���""T�S����m��;H����P��� ��4��/w!���AX��iQp�cIA0-��1��&}��r6m�4r�����'Y�|�	��� ������~�㑜$X�D�|�$9�3b�0���O�*������M�:STpO���%d!�om"\�i!��5�����*9 ����]W
�g%ul���F�����U�.6NN�{q֢v�U�M����1�"�k� �3d�M���0'	V��v�F��Qv/��Y%�V��,x$3ґ����Г/��L����7Ы��@�#�$P�f1h��҅P�bcz�h����B�mΝ�z�=�Dfr��zܣ{gz]8��V�k���k��/��(mؗ�
�'���5U�h��>8��"�;��۰�!Aw�o���R]]#���9�~���Λ,����x`GM��1COnd]���$��$�jͰ�A���こɠ��ɭ��Q�����`h�VD�I���n�=�Ͼ���=���k�;�a��60��t}�31�ư��S���D��DZ<�K�����-B���C:N~�_���I�/�8Ę1�뱯���:ζ�����U��u)Q�\H��z��}Az;2���&�@cu^&�f�����Ӱ�B	��E}��R��'R��V��T<�}�������Jt%B��J.�[�@LZ�t�����+�1NJ��,��
��$3����x}N��/-$�qS��&�rm�y>���2�x�-��$�#�&�}�{8;"�)�,6���_4�&�*���o�ψhx2�b$��Ƹb���`:+w)�W�x�X	�hh�˵����eY��t���+iFf���XҲc�5�6�y0P���e�Zpc	�8[��Fy����A^5Y����4׃�����7y8K��gR�d`�|��{YsAm?�֍�JwZ���YN�3^^�<�)_�Z�Z��z����aVl���N���!}�a4������]�����P<n�S�%�/��J`��'�޴6�Q��@io#Y�rPv�5���QŸs��=�&�f�T9d��H��=/��kx�<�K�Q��9�lKd���%�86�\>�Hv��7еg�k�.s�f���M��ڂ��G�ɔȧmŲ۾��J0��&� ^*�#n,���˹�c���'{�6�E,�/����1�=):.^�"��!_'����wԓh�t�sI�f�ֳ�n���>���m>������w��C���A�3拾SD3Mt�����ݸ�2�KcI�{Ccqd��/�
S����Ƞ��jMD(��J�jpd'��ٚ�\���t��P�����619�,8�H�H��۫�9������������z��f�\�c��R��2�48�5�s:c�n�<��贜���afs�Gt�[�`>g��I`J[GE�-�WY��<�ixw�/zpU�J���6U�zȭ�%���6�����,�
)�0��}pN�x'�=�9������\_�A{M��z�3�%���#�"�k� ��1��S�.�ӧ���q`�e(=i�9�KoX�T���
�����v[;c�=�X{�A��Ra7��I���E�f�A��U�2!	:mM�84�sٹ/�t��Mn0/��e�G���1�~mmf��Q:	��0����Ae;u�"���6������O�'�����
�����~�`�(�����G<4 N�W�/]�Ok"-|n���2�#���N4J��qxXZ���>�s��H��$@��'1����T�c����Y�}�K�h��Ӄ-w\�����(ٽF���W;F���e#r��cq3Wd�\<%�,���ck�Ȅ�Ĕ���"b`�����<z*�Ъ�.nK��3߿5�
���
�������{+�
Y�q=]c+����s��6�?��(�G9��=d\\��N
ښ�#Ɓ$.<�#�Kr�X�kÜ��U�579� 5`5	��7���(Au�y�U�g4��ק�q٘���ɯ#�l���胰�k�n����Q���Z[���2�b�^��A���W?ς�Qm�ω�!Zj���)=�o�Œ�RG�	)=xU� x���ʋ1q�G��Sְ������v	��,R���8�q\�q}j�W���)ނj(T�5�r(��u�E��|Hk��ֺ;da4 2�����>�0���>���� ��0d�׷�qs�<[�#9b�$����Ou`!�5��^:o��Q�Q�I�/�8"!����s�L�0Nܷ���թ(uD�Ȣ@�S[�c�A�mE&��#̜��ƟdR��U2k�?��E�	���Č����~}�Вd?X:���1GS���(�~�9�-$R��g�t[���7�=�܊y3��p��cI�f�����
d�X+l�>�|Ǔ� ����ԍ���c�5�I�vILeB�QE�\�\��J���E�rZ�.�FJ~~C�	D�{4�rOʸ��贈�C?�x�3�X8�`�	���h#Q��e.R��R�`�r]��^��ϛ\G��\}���vTZ��}\|]05kr�7}�r�ŉO�����K���<���S�Bq��uCӼ�/C���-�r�c��V`R���]�%!֣��۱�e%<H�7�����+\����z�Pq\�ΤH<�8Ջ��$���nͧ�M�����vPb��G��q�J�A�tn22v����ޯ'@����ؼ�H#;k�߬��8�C%%��U(ѮN�m�5@����d@:}�{�I�#5�<6k���D���o�Q�~���s�b$�Td�c>:A��Q��e�Sa�#�hq�\�rr����k��ջ����띭.HRɟ����M���.@�}M�BU�"�qs��:||��e�G�U��\O�ɍ��9��$h`E��
%��u-� u�{1�@��ph�;Z|��ݱؗEn�x�I��:+y��RnH[I�܌��<�P�s�=����ڻ���l�Igl[��������aɎR�xvR���7)]�+0Ԟ�w6舫,!<é�=_�L�'�@�=!�QH��XSD�T[Γ:�^-R_g�@Ͽ���!Wdw6��j�/A�j"HL�<��=��#$}��A8.�8=�~�[Z�C����6�u
1��[g�K�h�,��(���g�����v�MPd�Z���@��v�pz�y��G��.�<��A�*6Ŷ�-G�Ҿ(����4�gi1x�:��:�Г��Sixy�>��ļ��^���/8M��	ĲZ��b"��/W�|N� X�H�yԡ�P���o�}Y�VEU)�)��<��3\0d�l�8�Eu�$���؈�J���<j�G� �;�wR=U߆ǧyG+2�q��Y�}b���Y#��rn�q��@��0��m��R��P�g���>��F����V[�cЛ�qq���	Lo��jz��Y��ʺ��C#�%!	ʄ��x8���wTۖW�Z?�|5�POf��\��c�Q��p��tWz�F��]r6�0@�q�e�Hۥ��t�#D�L�:�ͩ8�ohR$�ާ�
/CH2
�.u�w~�B,� "��f�z��m�G5>2h�.�4��R �^���6�����ܧv����,�DX޶��N31�`�4�UBR�&(�� �uG�'��������ҜB}T��Zxb��ޞ��zz��1,��,�ya��*Tr����oP(LF���Y�1��6�grJ��,�nzْ�)��,�O������?U_+���(�l�F��v�+�=�ϻ���Jd���v���x���'�O�'ؒi.'/���Z{��Wc+'SCK����!��A�(��2�<�x� ���3��n��ΰ�U�W�@WO�X�P���q���Io2
`Լ�!�	�͝8;�7����hU�z�''F�-#�.j]�N�y-�4)��H�c��+L�u��O�;%�y٤L����&�ϵ�캲�)��Md�v]_�Xs�q5r  '��{�������iM=�R�����9�����t+ܬ���<Hc�Uq��Y��|��v��#���J����J���ؽ����r�L\S��Q�)�n�(��̵E����!i2vBjU+G����GsAi6��������p���E9`�*I�6y�s{&=��LL�@�V���% #�9�p7�Ё�.H�OÐ�@(��Z��|�)��6��t�e�<h��z�"�A���v�=Vpb��?oN�e�U�j�I���Kf���0-�;/;�S�9T%)����d�'����J��Q��ޫ��v�I*X8F5���67y�ĶV�qF_�f���Bn)�)w�������k��(u2 ��M�k?������*5��c^i�8uB �������Y���hpp��m�Rt�`�2�7.����o�&�����^��"�=��WG�M�pp����m8XBt���7T%%�V��bIH��4%I����뎯Mu)q���'�0mk�$]�@}r=�&C9y�c%gb��=�����Zt�����I����-��^�J"$�L���m/h�㝙�͠Q��
8�ׯ�0;��&7��%�-�`���\�4�as�9�2s��s�Ѫ�\��O�1X��Q7I�ksr�0,���e�k���%o��Y���V���uZ7���}GD�$_mři��}\��6�0���ӳG�����TU���Ѽ��P��6HJ�F�TQ}�d1Պi�m(�MHrZ�~�um1�ۯ�����E:�l��G�s[_��eP<�,Ɗ⸅��%�=ڌ¾hhQ)O�O�
��~�A��x~�bS��"��m�^�8��j��Y��T�L��7ݚ3-^�T��w�eӉ�G)Refk�xh
��'	�)gS�-(����Q�~�w&*,�R)�URr���)�U��,�9(X���&���os�H���<Qh�@d�|�p��.j<�U�3�^5�8$�c����!��D[_F���X���9�wi�/B�<�B�樯s��N)mzo�˴L�}���/;�H��l�]px���Ir�+!������3�U���-���ŵ��+L���c����9i�[e����VT��9vv�3�rU�C�xD���(�nt=��Ab�c�60�\�μ����t��֜I�X���V���1]�5�Ա��t�xsY�����)�F(�� ���n�	��XD��+U`��jN���VY�V�����ꗖ����ni�gvd��٬�ǺP��[E���h����՗1����,�ܕ1�����n���3�:��v�����[�f��	v�&�o�9�c�BU��f��-,=�������G��h�<�F�D��s��̀R6.������?��!�x����l��#t��|dQ��[�|��/����OYYb? ���T:M�8#<�+G7R��7or��î�7�
o�c"-���aa�o���)3ts a衇1�r�b~2.��S.K��X����$+<���������/�{D��}����g�"�(hh��3�sE77,�n�My v/�\'RmS� ��F���g�S��T�72��o=���~���	e0C�q������M0�5�CZ�V�� "ͳ<Dj�-w���U����A��*~L_��v�3+$pǮmA�Xޔ�7�>��n^�������m�g�~ɏ?x`�����g�����<=|�$��ſ$�0�E���,qR(����{�9��ז�z&'�ˉIh ����=[�d�Á3Մ�j���_}oΑE�>����h"t�t�]�dl?�)c;Q��
c�f�q;�V�נ���x���v�(^3�s����y�sʑ?�}vъ�`|�:9���%,��+��Q�Na{�ٛ1�L�ꏞ��-:�7E�V;�V��%�Y�|VMb�x� �� p$�M �"e��w��*��|��=J؍#EиZ���z�75�m�v���PT��K�ו��>A(���P��3V�w�g}����",���d�ymĜ��_\3�YZ�U�
]��[ũ��kTl���G;��/Ζ��L��{ܺ�_Yg��
����NWw�0����w���gْqk\`@F��6�/l�N����O�3⸪*�z�׀�����K��~��GMT;�H�ӌk�2�x]7B,MS!F�7 �7�b���k~�t�x)&NԶ#������sEY{�m8��3�A0��zb�b�I^>G�� �!
|��r����P�4�*����XǪ�%��)�V����}	+�qyz��������9<��ԗͣ�M����J$=��9+�$�Dɱ&*��������C�Lk�
���h�1I?�dd�d{��\�ܥ/�Vć���I�e���.`�B��R�Z�޳W�-_$L�J�H����Hj�s�XE`_�ξz�}�%e;����CV��*n�wG������vJ�ř��Mҭ�CQ���eP ���NFI� ��8ӁR@�>m��G�1�hͷ���6���p�;�����R`m��𭂖�EANrxJ�%���n�͍J\�n��fo�J�y	�`� {«�`�����h�E��wѫe5[<fh�@�)l[uY�UV�G��G��y�'���p�$��ʯX�W6�p�bel
�a�8�Ĳ?��[^|�g����G!F_� ��r}*g6�GW2_�I�a�攆O7��(qh@��+U�p3�tU�5gY�IZ��6��������;���Z
�����=��k����<A��=������'v�5E�Guz�^�m��ձ([uQ�'��Gqse�=t떯0����o��k]��($h*Ogj�~�P�s"�[��|�I��c@
k��{Wi%J�tm��i�����pj�'/�����0e(>���0E���n*��9��ua֮�w�sU���D ���EXF����k�p��$ǚ����������:D�}�WY�a��8\Ļ��������:V���O���8B��$���֨b2d�$}pNǂ�0��� ��IcZ�~��>�+�@R,�y%�v�.3�̬$�r�Q:�0��=�!�����.�`�����3��8��l� l�2��yl8>W�G7�z���Y>/�.����m�o��lZ���Nddr��Fgt�V�(CeZ);ߊ�i�ͿI��n�A���Ǧ��Z��!`��p�.��vWʳ�4��|���p3:�]�4����5�� ����[1�f|OcE��=y���&*�����R��)�֋�Dz�����DK�qg����: Y����D@�s��7����:�e�J3���j�l��a�,�ԕPɪ�"ُ�uϗ��`��ϖ
<qJ����l����C`�-5��9bI��-�NT�OT�`bN
]
�F���\�%�7�ު���uXd:�Z�� �qs��/:�p}ʼmæ��e�Q�m�c��NR�1�{�pF��N��f&��(�z��C�H���sIU�³�������
m���l�&m{�,���W����ǁ3�JZ��A{\���xA�&�L�R}!�p�pǅhwx^4�_m�dVoD�(��ғ5�Z�u`���G���"�3Y5����簫�^ Id���Ї��;_b�͎����G�˓�P��W-Mãw�>����aߢ�X�,l�zWo0a�8H���)s���҇:�Y����u�D�q�!fw�� �����2���G��@+ϝ@F��Ӫ���������t����_g�YaҞ�/o�������T-���Bv���Tg�`P\z�H(ZmW��y0��x�»Ľ
�UF5�Im�茹�oG���8�GoY�7�ko�uQ;A���2eH��טW J��m���,nXK)'�S0�s��U�h�*o�1̒6�dR,Z��{1U"�
>��M�I�I��k7"��Ax���z����/�|�a�5��ǐ	�dK�÷P�����_�%&���I�"��|�ʬ7���1{���x�����(ޥ�X`
��+�P5'i����k�Y�3I�:��KU�1K��ܶ˔��ΎH�Ƿ ߗW4
��FE�;#? ��3l�Ѣ^7ˤ�{����b5qQM�XL��۳�g��,�Ee@�[�w���hU;}~ O�T�1�u�bu�qAFf����V ��1_��C?Bؠm��M�����Q���Uw]��9�vga�S��mjH�ܬ�#.�\�9\w,5����AY�k��}f����wGHa�{��a&֐�rI��_�_kM��t����6�KԾT��˞�Vj�PN�hy
N.Yl�����޸Q�,ǔ�1J2!$����y��ܥ�1Mm��
�2�F�8f?���ٜ�*V^d�ӏ N�)��J��q�"����g�����zHi'&C=��_m`?(�j[�?������/����XNA	`��4�#���x2 Tm�>�Le��U%��<�G���+l{�s7E�K��I�m�G~h*N~e-{/�Oɂ<�W��nW�O����U���"�/r�q"e�1Y�$�E`�Rz5�KF!'����i��-]r�ϐ�9��=���ғ�8�$�����2e.3e\[f���Ʋ�z�@����~�~h9Q6�(��X�1\��s����]b�r^̄U4���HE-��80�xc�6�p��Ҳ����v��%�W�� u�`��i
g���۶�!�V�k��s/���mE�H 2`v`�Himt�u>��	�`/�&C�)<ټr8���P�Ǣ���L ���{ϒ����ya՜��~7���b~A�#Z/|-L�J�0�x�g��	�D�\���5/�t��_�*�R��D�g�Yb>�����!D,0y��P D���M�%or����ܖ�0f`c���İ@�x�c��P��Au�~5Fy�L�,�˄V2"],�DǦ�JE/ՠm��uհh����tmC����ص� %G_뭟H�H	<��Wu��W@v��r�2F ϶��M���:���E�5��t���Q����+�>q�wµ�����=�g�ɛCUG@pW�s5��,��LiN����3.4�c�V��`X5�娢�$�5"u��:[����^�����G���Ժ��@����w�e���
l���Rm� Q��`�E0���
����$�[��]��^�aZIaňA[a�" �E�ߊ��B%����l�y@Fj�cІ���H��[qZ|�����Jjx͸�6�c1���Q� ��ô2;ey���9�<��{l�r�P���cu-㝋 %�H ���\�N�|�T ��W
T_~gc΋��N�r��9$��b8�OW�|����^$����5�v�;85����	�sH(_�4>X�|��т�6��A����\5&�`�;��d�v+�֮G�5��F�������7. "D��kj��I�n���/
P� L�F9�&�)l1���KO�w(�R������pp]���[~x����v�t�M�"r�Y�MP��(��;&�ЮR���e>�Ep8��TDڧ�G�!��m ͟��PvC~*ׇN�f,�IӍ'6v-�0R�\~�u��	%��l���*gs�ϲ��v��,���v�k�M�7$���Oz��Ǟ��,"X�h|h"����J��.V8Ə#�����*�eSJ��׻�G{���7v�������p���FKp�t)�K��"�r�q7�I~p΢�zvz̻��=rW�@UjhI7tS�QpJ�S?`����� ف���}�.���/�7�K��f��NsE���iy{�F�I�.�M]��DH�Ȏy��[��l��hZt������:P��S^�Q�� r9��T��UsaR�)u���6�z!�4����xNG~�"_��YL�R%��?/�f��*�l�{��1mY.Y!��Es�a�n����Dip��c�L⧴���"�K?���r![�	)Mz�k�@���E��ܳ����܌dv���v����!��Ω�2Ag���WU���0GEh�7i�c-���K"u�9�Vc\�$��5�خH���T?vk�r�4.l�)	�/l2e-E�}ŉ��A�3	�r��=K[�s6����G&j]a��R3�Hڠ�o�����˪כu�ˮ����XF��9v.��^��0e�(?��%�f�l����3����4$A�y.���3�8Na\zl���L��L��5�сc]Z���G�|k���!G�t��nc\u��r#'FO�Fd������yzqRj�������/��:�����Ŵ�I����m $D�*�q���
����K�V�8S�la�����S�,���n0���\�~�5AE�`$��J&�f.P`Os�?�ln
y��
�3����ԟ.ϒ!l%�8������L��~V�@Z���v� ���dɿdy���^={v�7�����/�J���\MƐER�U�|�!������Q�G��~�ʮ�;ht#����@��6��ʾmD6E��Gh3��LRѨ�0�T*ߛ��X�H�6��S�|����3�B�;NF�o�y�.P��u��?8�G5c�0V��ؿpy�{@��j�'E��*�T������%�1"`Y$^��'���5w�{��q�>�¼9��Σ�4��,v��U&���`���T���_V�Я��飆�~��Ar��JFB1���g.l$�ŀ���N�j�HQ� ��:�~��+-5���"3r�ޒ� oN��(8V�� �gƌg|@��g�H��h�?�q"-��`���[�;;����iE¬���[/�w;ݼ��==����vnR:V-�!&�z!v��p H)��������
H�����$��7��#�?�&e?����ItM�6$S"��}��y�=������Ge�ui$ �֢2�f�7�S1n N�9�+G�Ed�o��e9�S�[�\U�KC��rdRw��C��vVIwv��a=+!Y��₉/ZV�6�Ru�9	W���~��>�7��B�7�z�`b�Y\��*���n�K��E���݉�X���e|fO3�1�a�	�[�;�!=�2�v��u;P�h̑��,��g��}�Up%F
1��l�:w"�U2)Ml������"ߟ��k[3(��������q�Ze��*tK�T�5o��wb�<�,c?(�"�ŵ������k
���t��ޣ<��`�u�ي'$���#+zW�1_������H����g�.jTO83E��w 30=�oH�������;Y5m�Pz�0�A#�?���_ˏt�^�8��h�԰�k����q���y�X	�Mj"zIp(���4���2�P��ZJ_e:��@U��R�2F���"+>5��޵w8	��d�y�O��{T�L�_¾�BKI���%�������D�O��M���3����98J�(!��!Gqe�1zb�aB��k���GQ�p� ����xr�#l����	�ɨ����>0t։7�{t�ϰ��E22zT`ݐ�I���n���vs��T|�@b8;�-�6��__e}&��#�19	k�]���[�H�qG�� ]������D�ۄl`+F�	Ҥ�y[��� ����y�Z3ԅ�F��S���{�	M)�j���:mT���^�h/'-� �bR�!ؾ�Of������x6�5�����ԩ�U��t�W���oS۵3�&���O�*��#y�1�]�`=����*`[i_c�N)�.�:�
�v��&��#S#C�xi(��=��)�0���\�����LX�?�]�m=ȶ�82�ܯ���7`��A5r�$9�J���^�NQ�^qo�⥟�
R�)8�����`\C���J���E�&C(�U�YY�¯�p�g����e5�RK��Q���P+���{��z�ATu���?��H��W�z��e]%t����|��/8��fOz�l=$U�"����Ц7x(�{�z�XǍ�T�N��A�ʼD���B��ƪ~)�Ks?����r�Xَ�Ms�C�������Ǽ``�]�Uk��<�({ V�I���@����K�eu�b�����20�<�(�y�����^{p�(t9_�L{0/3�K`��btE�tM�v�G���4;exi���5k���V�����*c"���C�ܓ�B٘k�S�!�5�&X�@DJ(
�垺(x]\2|�\��wY�-��?��~q$��u�یX��`�'./�JıHr���/ײ�R�,�q��{��5�_�l��n�9EI?��+)t����HN-��/�,��
J���+g����m���"��;���z��!��\��NĄeo|"T�%W�YF��
��]�:V%r�.�ٕ���Դ�C��l����,sL}����X/ò������������h��@����7Z0Jl�HSrVҼ�`��D�\M������9���p;՛h-[�d<?�NPB���WW�1�p��>�Ā�6���5IQ'
a[%&6x	z�~	o�$}�"��RJh���9�������D�qt�5(e.���w�G����d��-5�|���O��e{w�R½��p鯳3��li\0�WSdd�f��`�LIV��	3��F/<�R	��o�����E����:��A�L*���4�d������{��N�:�unl|��!n�V������c�Ңޗ��]�X�=.�X'T�.�(d*s�a��m.�g_e�9k�[�c~C��2� =���D4��?���C"�L���$�z_�4���6e�ǂԦ%�&��G[�4-��w��[B��z4�9Mr����Ѷ����Pǒ��Û���S%����W��-�F喞��W�`v�m�n��]{V0s;�Q`�TUr�Etq�_��cL%3#�%������a��g�u?v�{$�KL�X�\l��Jo�w�ƍ!��M63�2|T���kdJ+�Y_څ�h=^���b�/vsh/�pt'V����C{Ϛ����8X�MH��VU�D[ �))=�3@�0Z�gvZ�*"����1d����%����_�s���g���N�Ҫ�p���dD}��wU��;f�`T���b�@���I�c܉c��<��y������Uv�����@��-����Sm��oP U�#0��[c�5ک+�N��7���bP�8�QCҕuH���ib�GQ����+��KgU���b�m��*E�(��q�N�g�}ݧ�(FiGC�`�^�e7�|�bP 97I�qTw����4_bܩ%����6��Ǜ����^p˞N���i������t���o��e��8c2���:i��Mq.t{�_sK'ͩHe�/x�<E�)�랕�2O���'�_O"���B\���-�7�Fx@�}��{kK��t8�`���q�p����wqT�xN_T����91_��y�
3�v�sD��VӚD�F��ǰ������B�@�Dr�R��K�ׂ�&��zS��\љ�䂫:I�c0-�>�n }x��[lH?s��_>+��\ʳ�g
m!,l# T��w��SbG��=�~=��
U[;�H�uÀ!|�P��K�N�	���]9�"�Q$}&SH�٫%gF���jkn����5�Hw��H��GJ��pI!���Y9x�|���݋<����}'H���oZ�hAC������3cI:�*D�7]��d>�!(��NZ.B"N]�t�����\(���X0؛ co���&Q�k�gT��f�-Q�Xڐ�˦M;�@��h���Rb�9���3���w��X� iWЩ�-!�m�A3x�!�
t�L��lǁ��xb�
�8`p�%!�����ߥ�@�����k�[��5t��������*��6��g.�MsA(�|�$mZ�]�^����!V7�A�w������MV)����<n} �?Y�T����r65���cs@�э|�P�p�4ؿ򋸌�G(ٺ���iRS�֪�MPR]D�3x+�nq�>��q�]��0�	��
���� ���h��АZ�>���9����yQS�qp^�.������i �Cf���|rλoy.C<1��� ��e�R�6�5�Y�c0�$�X"�zV��:EQ���e���2ͼQDDcz(���t׋}�BS�
F�E����7�ݘg��e�ǩ#­�+�L�h2	��A�R9zh"`�mή%��M�<E����0D�T��"ƿ(�^֩�*�����d�f�0A�;��pu������@�@��;d�M[*�����Y���;�'����H����&�_�[b~�v�'��f ��z�3�R��X��7�����*���t,����O��g�`��5-g� �+g3���v�Ƿ�Z ��okb�����Q쎔���]*�vc�L2O�c�[ᳰ������
�>�#��!Xfc�\|�+Ԋ<�V�K#��G_3�"}Ϥ=ؒ���u�M�Gq����TG�a)mz�l�o�vf�����wР��{�!����D��	(�,�+�|��R�*]
ٛRğCQ¬|�6�XW���uw��}��]�szAEĂk�1�t�as�f�V�M@���oR�JL&8��GYl?e��x(*��R1��-c�s('��O����ڠo�l��� B�ZmW݊ځ̚ZW��o�F��w�Fxq��@k��P4�6ql�ia�S�b|M���z��A�c�(�сN���mo��e4?�s^<x������v<�s��8�H\���K�p�3Iwj滴t�P�yeN��'ֻ& �����G8˓�-ՠ/|\��2��.���S��Sc��xZ�tN5Kh��OC�<�1sdŖ�_{����3��UY���- j��Jv����w���f�{�Kj��5Z�A
VM\���̴%�g0b�iԷ{�+-8���Zgn����)��mMi��J�s���'�Ƌ�!Q&3*�Hz�x-�}�Ҽ|�tN�퉊��9���l����;�L�݉[{	��W�Ju
��;T�r�;%�Ǯ��+��_�<�ŭi��.��x�pE(�S�a%�Z<�%�<#�|�������SbZ�5jwM`����,�0���ۃ�}w�hht�>�:xn;Ӛ����}9Q�|+�'^�?�]�R�'+2�<����NNQ	%-��>�R^��ճ�qI���;��Z @c�%ȉ�8�vg�.u�a:V$qјg�T�a�����Y���hT,WT��\q.��_M�j,��6,2x.�f�����ap�6%ʈP}C#���=��,t��ƽMy@��6s�[3�K�M*��;�+?����K�Q� ��!�~�)��s��h[\���}�k<�I�Pt���@�\/��Uळ�$�0%���*���5��Ǭ�v��'��Z�g&����$��2�׈����`F����(�bw?c�Ω�!Ѩ����B��O!)�D����Z���c}��N\� �W���Ph�;����e�LR��ܦ�T�{����8��������*�;5���_V�>�M�,��0v����D��c�}�^F�̪��Gle���CD^��,[����	uK�wv_l��̱� r�g6�流n:�����N{����c�H��Ʌi�\�M�\[�Z���&�1�Vy�#<7z���b��O�y�S��ZJf}�n��f���ܮ"�*g�ӱI��;=_"0F;�9��v�	�;'�7qi��ȕ��ք���GLms���^G����"�k�U�8f���f8*r�d�'v�Ni;|������A��䬦��V^��#g���d��!��3�