��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E�����>_�.�*�(e�{��?�4���I�x�Z��iWڲ��~&X4��-k��l���h����[��J>�B��:6��Hn9+}���xUU�s眓TM��Vm.�#�/cm.J�߉��UDX�ةo�!ժ�]>���>|S��Z�L*�EM ]���JXmk��J[V0�A��Aǧk"�\�����L=���7x�jt��Qc>�Sv,Q;���h�(�kHt�Oʍyh3p�0�����t�"��͛;<��'�޲S	[�^�E
����;	*��q<�[�`��{��LTPW��ic@�Y�Rxb��hI���w�7O��n�f0�E�m!��l\��6>��_�Z�5m:5>���C�p��P)�<\�.�|�PC��d���3����f�4�p y|M����h4�Uw���\������@sF��h�D����)J5���ѢC�E ����0j[��~~�����ű�ō<>�X/b��y�x~�D��ƻa��u�ae�-�����R��ڷ��j���H�;�B�ߓo��%�'V��3�)j��2��&vs6�����vk/]/���p�jI�l� �cR�,���t܂�����U�y��"�ɟBh����;��^��]ڀ'Q�	�/�N՘c���`i��
��PLi�w�am:Y���\���<>���*1��!�2��U,W ��|	��u_�]��|�����'Kս�i�N�C���GD[�V�gN��׌S\c�3���e�&w����9����f��#)`�%6�"���GG��ذ���[閯 �}TXK��d���!���l�nu���E�v���u_>?�ԏe���i���� ���ō�:�`[7y�#8_��+�7H��7�S�֊�����l3���M��8��9��pi!(�]y������N9�G!��9�JK]�*&�A�KQ�O-�⨋<��� ��t(]'ْ�̎�6�mO	��g��>�L���zH$�(���󏏁ޜ��!f8 gN�0���w�℟['Ap ӆ�9��r/Qֺ�����s�d�3o�,��X- ��0���j�9��t��S���5�t��w�t�L�i��P��6�;E�Z������`_�6;�b��	g�u{��Ø��N��d��	��qK�k�Tꑈ�����5�i������+��K�^A{�8� �
�8{�(|���d�����G��Z�T��OC� ��R�|��@�>��g'�R� A��	T��&�V�����ׂ��`�&�T�Gmw~���M/���m;{wydoGd��7�ރ_�O��؇0�_���=��l�n2٬>��Ղ�Y�&O��SZrO�K�չ�[A�ña�oA��6i6�k�`���|�V����O�"Y��f|� W����
t�޿��׽c��C���;ƭ�����
�|B�[�dr1��w��g��]0&�-�.�|u	yC�â�g�6!��9Q���X��[D+�F����"�4&��?י�j�ٵ��IQhLQO�'q��h.�,����&jM��=d�@..Rg�_�&�� �=C�D�I�K2��鲛�sj-N�R����ܼ�;�\��b*RM��e`Ȏڤ�Ř�-Y��&,�b���k��mK]�/2E��?>��.�0��.�~H�4TZ�w�ҸS��m%������&L�x	�\$���v%�zԲ7r:��Э&�*�$ �[�#�4�S�������w3��w�.�u�{�������|�� ��&�[�
8�����5���o��W�	ٮ��&�uI�����]�?���J)��މYL��AFC�k�1N��Xi��sTR��2j���䮳*r�9�L��XO�b�,��ƕ��N#WX^��)�`�B�:�N?:��$VmӬ�� ���-M� �G��>Z�l;[��#1�r0�J;��D*�B���j糷Um��L�N�)V���n�`��nM�jL0�o Xxe��RU�F4X_��D�\YN ��d[z[���!��lm����V=)���TkԴ+��xY��V�I5�)P�>1+ڝ����x��I��� J��V"^��J�!��<B7i���AO��_Je�E@G�4����F7妘��Vc�<���ɞ���āQs�+p
IR��+���@��\l���u�i@`/��Z�ɋ-970q��N��t5��U)~�uN�P;��T��m4��B�zؽ��L6v��MG8��y^y@]KI�J�6C˴4ޒ��V����A#|�x
O{��V�͒�Eؕ�>�������\���ѫ,�'����8�;�V��	�8�'�����4��GӔxo.�G��0��t]���פY����U�X��I('Bӷ^_�z��xj�IO]A����b21.:'��:GdD����@��f����OK�"�X�j+0��k�Ziu��5��`*s{��(J|O��3u�>y7V���=4:x���)r�G�O兊��? ��GF��o�/9͞\�3B���B��;��X�5"%�INX�b&	9"�����<�~ �Hm2Q'�S�"<��w�ne�>�f"�6�xw�9�V���E���z� ���y5��,'���*�F�����h:�r���x4ߏ@���o���c�8w�W;��S���������T���i/"�m0�ľ�`��غvpP'�Ϲ���B�:�q�S�4���`&�/��&��x�u&B���NyC�D�x�Ln�����ž
���7@�t���?�v����H�g�	Ŕ]=�����w�5,�~�����-~TD�NEIG\��W�5���?2���s)�w!��0 ����CI�L��|&1�;o����Li���̳��ӷ���;�$�n�
i�g�O�zr�9$��TK7v  �����Ӹ0�J�C���t����A����t�E�EA��Y���q ޖu��;��e���_΢/G鳾x����^�x���C����ne�[�zO"U�[�i��Lt�l�}b�=����;�&)�ƀ[����M:H7a̫��tz��Qm�qb>����3/��;/��DZ9�6�X˒\� ��!HqC	I��nRT�d+�#��o����F�c�k �J�<��N�~c��{t����`�;��\�T�1�G> 4��������9�n��`�|�P�A.�
��=�`SUtry�9�i�*<=-89�]5����=O����y���f�}���/��X�K�L����+ ��犆�l�3�D~�7+����͗Ewdf�\���G��O,X�����$��J�É�@p�w��Ʒ\։h���{!YQ��V��Ֆ�D���Q�(�{qV��{����߂��r<�`T�^7?j��� h
��%�D���������;n6樂ð����Ծ����>�˕�4�Pg�ʰ�>J1Y�]���>[l}�+9\�s�6EQ:�XT3����m����*�:�}mdW*LtĜ��=&W��	r��{�Ϸ$I���O��2x2���+�T��/<ϸ���痛YqEU�a�����M�����޹��ۮp>��9�x���� �Ua߄EL�+��6�ވ�>�(GX�@*)���x������D���G���g��^2�rɫ�z�a�4Ph)Ƞz���h��=�[��@����I{:�@̯_d�*������j!���,�u���;��	'�n0KV$������6m��ZX���-�V�l�V�[r�v
l�DzOӃ`�)U\�G�{
O�mھ�=%�xfc��r%l�����n�{��N���d�ʠ	��� I��MeQR�1(X�yZ�:�aP��/��Q7�%��"F*���!+H�D14���7���J`FoAX�D�����^A�%��ߏ�Sz�t��2�t'�&��U��* D�6D��˔ˠ]c5��[06�m�@�Җ���HC�<FϷ'�(����M��D���vUC��1(>��A���bI j*����+B���'SI�_]�߲�6��_��\�
$oB��S�}��Wt�����w�rL�@L�������B��ЖH�Ҷ��7.׀ݷ�|t�5 tfS���(M*��ص�^(��ȉr����$=�u���)���'�e�RF�OBE��BUTYQ�A� uUS}l7�*g�FML������2�X��5�ֽt����b��i�m�Ԅ��֘ٳ�cb'�3r
�g�a76�)�8�=y����'���c�T���o�����^��5���n{��!��FA�<�Y/@&= yA!��4.�nF��}m�>��@���.ȴ�J�v&ܹ�j[ԃõf]>��N>MTm��k�;�,ao�d���ti�G�ȼ�l;]܍[�L/��V7B�_U7-� ��q���Xy�xBi�z�x��6��Cn���E�O�!���?�/1Pxm�������� ����Δ��m&aG�@�p�y���U~�$Ei�r�χ}/��FXap���N �;��6^��rPE���}&G	L�\�q��s���T7�f�8_l*�(=�>�8�B�8�3�X��C�0�K��#O���X���3�5��]+bc�QW����GF�?�-�a��H�.�����4����LGht�v-ɧC���L5IU����d�_��<���)�}g]�f��2{�DܿV~Ge~2���W�<�>��8�n{��w�"����W~ۀ��g�
<:O5~I��'Q�²������/�	��`�
p�����a����y�\|��i��ҍ�Pfd]��{d^���|u�Ō{��;��Oq�[�^y�n��$_��.$�4��_񆿇$�A��b�Q^��u��8?��!� 9@�v�t�伨:�)�&���5T~��!�Ml��F��[:�IQ@���Mđo#��	�Uj4�ݥ�&I��w��v&�e��?c��>�Z��:06f�|��-�q�>�{��Y��F�'y�܎���e�7|���Bv����R*�y"L0.A
��+ð������:�
�q�-�f9n���Ĕ `�m��O��&&�@��@�!a���+~�w�������y��G
Rhzb1���l�����ǝ������Y���p^AzQ�Ӎ=qd��7G�@�J�
O�(�*O��a����a�� S8�IIɟ�I@�-z�Z�߃4���f�#�/���:��'2rMfq�f\�z0�2ߵ����O�W�������b��;�Hz�f`�[O�3M��1��9��+x��e�^CY{Hri����h��z�Q:�N@�ӂc0�f�S'��4"瞶�L;-B*��z�%KL�7qv�0�NQ�E��Hc!�p,U+�O��g�t���?Z@��ߊ��'��.鏇�-��[O��bL ?��|j62Z��v���t�4oȻ#��ۮ5{������Zۨt �d��w��ӛ� a��\?�x��)w��<:{I�8�Y:��ˬWX��!��_p=6�d�+�K��'���hm۱lx���Y��r���g�y��K�U��B��3 ��ؗ�pьv������N�#�N��u�� 0b�d$a�Qk��e��n�����%��Y�[3P�aY�$)��J�ݖk�u3��v(C�h,,)�٪z��f0��欩�g���'��6<���ԛ��ڞ�P�IQ.,��X;�Qu�w#��H���`�����Jo⏁��]�ܰ�|Sc��!=��� �S9*�w4�����hP��w���;+U�|'�x�$j�Po����\8	����}��?%����8?���Le�hA n!ĕ���!�ep����i$��%�ҩ�� �G8�1uB ��O�A���:Z�w7B̐��g�|�P^`�m�6uI��:k�5�;�Q�-ĳS$��,�~�>�T���f �-Jh���kմ��?y��'�`��hy���[����v�͗߼���L=�q�̆�ɏ�֤s��<�S�V�KK�(�+h��bpdhڱ"`d^z:R��,0?���靽�Q���W�i�"�i���a�%�sf�b';5�81��Y���02�Fhޜ.Ȅٳ�fH�����&�����Z��8|F�*�{3�;\X~�c�<WUA����;_?
�a~i��y��?����hڕx�
���b�\	�ݡ�Nҟ�[u��7�tZ��pt�3~�sH�|QN=?[�`��&^�"k�Q�Wյ��|1��Bjk�p��j�e9{zӋ�#0�[��gc����U��ќM(�{�K ~�@�0wUy��.7wkThq{�'�-���A���cj|hڗ]9#�i+@g6�H��+G����k�{����tq�����؝�Ԗ�`l�58Җ\$�-������b53O� ˊ�#����M�jSVcJ�wj�ڊ(���"~!��W�����l*2Eшz)��S�߆��KK��'{�u|䳏7)�D
�P��\ӈ&�,�s[i}��+~�]�T��I��`��ޜ��!�zr󬉾p�(���[�&�@\���&��W���ye�Cl�x�_�-uA�$EƐ�恅�YQ��r� Ʋ,��O�DU�q�LR^`�-�k� �r����Ǎ�k�g DxQ���W%��Co��bޑ�,7a�L��q�d�����\���[_��<x����]P3;�m.�g�8�*�Ѡ/)� Uրj��O'�~����oJ	��ƷD�
A?j���{	9��lR3��	넑�{�P+�r�O
�)mj�0rI>�ٵ�8 �
$zۡ����Q۩8=v~U�ê�܅w�J���Kmm��qt$��5�^J�E�7"4����R�ĺ�枚�[n]م�%�����uKA���(����"�O�_��a tE��5��$�g���Sk����z�o�a[���^���߀!���~��d�#�v�-�?�M���UGV;��n�a����ZL:��7,��?�I��DN'P]�dw��ld��Z���,�/���n�U�o�ы��~�O�����LS�Bwx�:%?|��KRߒņ��;GL(��5w���5�݉��=�NÒ*��_��K�#���Nb���A �hT�m���S��Wc?�U��A���
+��*23���^ F����t<��%��3O�l��bi����`|ʋ#��8�\��ssY������ܞ���1���fi�)�gI�?����v>�x*AA���r�Do�鯿Ps�bU��)�����Ue«��S#�L��Վ�$rNHh��=�
�.�c)]u�{X�����(��l�w��a(k�Aᵽ�QC�y�ΩW)�dH�c���	;Q��U��=��α��Mg�<�9n(�������@t�L3I?/`�V���]'Q���EH<E�Έ�O��ě_��7��=�IV�/GW>����`�����-)b��
��<�#T�/�3���F��x�)��JO��1����	��n��=c!��|����+ڇ$�,�h��,�=Â��ٽx�� ~�Э^�-���.G��# Y�xy���ҍ3��.��|Kf��ބ̸~bl	�H�I��lq|n�Sn���u)��ϒ���X�9�	�i��@��}O!�0�_�S Nc��<�k�������&Td�UA*<|v{�p���=�.��Z����Z�f�c?�My�F%�Ɏ��:M9FK��K�?B�/��!�_x�E- �V6<qS}�3X�j��4CV��'��s�5�5��Ԇ�\?�*�|ig;5�LB�N�kU׋�dg���c�#��)��f��=��do���k���aE�S�MW\�,�g�W*~3�b2q���{(,1:�9;>3�%/����e5%T�"R�Y)�6����{���^JGا����sp!�u��<���7��]}��ۺ޷{UF�$��Jq�V�^�^4� �Qo�|�(^c��?��'*�U'	��*�1(���Z�%�0}�n�b�(�o\Վ/$��{6��-M}�?����mh�0s{%���sL�� �do��NJ����]}p�<`�Ǟт(�~YzEK��@,h���{�2!m��0���<L� ��lA�ܿK��.X�G�9u"��QI}b��0yU&ZoM�(o���maP�����.��d��|\���^ţK��Ч��!�9�}Xdq�����em�J�K�ӨEUH�oɕ��h�W2�m���D��6����]���w�^�}��79G���yh�,�C�B	ɾt:+�"#W���#���H�k_�R�J��0�bW�3];�&u��x}���-�m\��`T%_4D�="��5����;�����6�+Dx��qC��&^.�r� EL�އ�ʋ'�B���KXV%������\J�C(F�ꭡ@#a��se���w�݆�G�et���{���̻i�UXWE~��H���R-�P�Tw��w`����i�.}�����f+0���y!!c0�o�3'^����o�v�v��n5�}��퀬��Ķ	OӕLp�q�Z&&�p�+��^H1U�Uu��.��3Vu��*�� �%�����Gl��Ő�����p��7;[?mp}@!� ��f�S�Ķ�m#��+�|J'�vg�u�e�x�5�t�Ѥ��ضL54�"j��Db�n�ΰĨ����d;튋��� \<РɛL�G����������غ�����f��[ޮ|�p!�Q��̬C2���C	�;>�}%s=��4� *'���L9cE�N�e(-�=RxI(`�18Yn N�_i�O�{�{#bh���N�>��Y��:쁯���YS�l[�T�V9����]c��nҝ��O����7��,�eG��_����� ��fY�aڊ��TS�^'�V�����Y��J��oVm�L�)�ZC){�cR�'�cl���,��$��0�g1��7��i2ht{�����/�k*��u_)��O�e���������6���i�b�j�D�3o�v�³��H�]5*��#�����$`���ͮ��n���C�I�2�](���t4&��:_-�?ĥ�*E�j�BV>c=��.E���Lm�S��<,�
��?�+n�H�]9���$�B�ߗ��E֊g��q��V��b��%l?=�	��FG�O\����@,���%I���W�ք>�f5((n`��� ����\r�"�������<� �e�d�i��,$��}ځ/��Q�Z\C7b��C `B�Rum��-,D	ɹ��<\1��J�7�a0��|"q+���'9��ٶH�n�CP4ļ��qP�G�Vv'3M;�~�͆e�{r	��Wi�0�ލ�ΐ����ɩ�"�t����ԹwF�/�h�����=e�I �7/������xckH�q%D�N�� �K���%"A2�a���6ELy��d��
���U_�a�x�7��ܛجQ���C��W��x<���T�ŗ��Rټ��������@v�pv�~vZ�=@{΀�j��QU�O�O� �f0����Zz�?�w�=���;�S5�*u�RE��R��7a�Ω��gx^�\̈́p�M�5j,��"ʮ�ʹ�C(�6W��v3!���l�s����Ս���Rht|��N�(j㣨
���YL�Yh�O�]^\�yh͜33'p�ۙJ*��g$��}����}+��.M@�����y��}���Z�}R��,�S�n9[n��Fq7��tWv}�U�X�����N�����s^�k�n�q�k�ĸD�+gc��rܨ�,..B�`�����)i`>5Y&p����D[R�fz�l%x�}�C�pt=t&N[	[h�����*�J�W��zO�*3���^��mPQ�� ;|�����(zY��Ӷm���(DM��M��ï��2�`�L­� #���8Y2�5iv�1��MG��>�5Mtu�6���Ø��}F�A\c8�b���q����K`�ױ�����.�_�h�Z�?A�v���njH(Na��{�x�ޡ�OT䑎�^��
��������0��9��K7�I����T�v�GpdMM�5n��f��U�F�u��^�>0��V���a������A�I� ���.��|���z��I�g7��nv����_���1h�H�#$,C�\�#�V�mӇyY�a��B��D7��|� �=R��;��`@��:T������)���U��-��x��a"���ͅp�������� ���bwQ�77X���P���VbW���
�(1��N�L'�������K��:�W�SXrMd�Iw�kWh��g�7*���ёx�5a,�R�׵D�Q�F ��u��lZ���I	�w��P3&�Ff�(�|BǱ�X��(D'�	���2��([�Ӫ�m=��z�p��sJh��j�J��j�����	TT>�XP���\��48�r���G4��?;�����)�ӧ8*�K�bӹ�K���={���9�v?���6��؎A����ޤ�u�YF�:Yo<A�`�=���N�I��~���R╳��	0���GY�Ȣ�V�`}�ǎf�v��UjB�.ų��G�<���-��J��򩅼n������(h���g�yo~ �4��st�N���?�"`���z��ѳm��3�8A?F���&��1��SU^��.YL���8��������(>;䔇'�+�²6Q��P���kG�O��cvzУH ��C�]')5�_qc�S�	�B�"������4�+��E��1��n�����Wu,,"�})����f��Ei��
�,.��W�{8��fv����{�dԘq�k��>���f��K�݆5��b9���AYںS2p�a�[��e���%�*�ww���&iǼ�xG��I������:�Y�`��3gQz���>�/?�W�{�1ҩA~� ���+����y�G^'�/�k��e�g��08Y�?H���3�m�Xc̤���=4F���4��A��?�B�nVZ��`w��M��h�����j~*����},d�k)��<B����0����$����1���������ľ��啜	[�Wu��4p�ئ��X�����ϕ���Ů�4��浖>�*���� 1���K����Xz�k�ҟ$W����U��H̲����R��yR���V��C���
k�sЄd�G%�.�����G��q�.��0�q�X�lɿ cP�gaQ?oFh��d�+o�9���"�j�F��G��^�fL>�G��z�K�z�m�(��b����UY�ҳ��c���DVP��o<�o�uv����U��r�=�s��|����U�G5@@�F��S?�\��5R�A��38Ts�W>�����&^h�0���Mq�y�%������i���Nv���Z[� lp�K]̮��-��g�w!��!s 4����.pA
���]�$ �ꃐ�/4��<�^����,s�t�!�H�25t;0=�6	�V���T�"�|?o���������D�����@T�����/�OKۑ
.鯚�e~���IJ�3B.A�?\���a9�6tӵe�����a���YArm��YTN�U�%����穚���xsX[�|������h��{�����`��g���?Q)���q�{�g$q�n��x ^ut�58�zim��Z5H�1�չ,�[��%�S�.�*tv�Ȱ��L�~�dL;�tC�q��������n?��P�����~~���W����NQ�No~�lqФ���_�VL<.	����U���X���!8n��)U��^�C�o�
�ѐ�
:�;*$O'�°���$cz�*齛[��٢\:�uqr�DP�i�O����¿>W��/��ywE��X/ߙ��ܦ��k�{��kl�z-CU5;k+�&C��2���*N5-{���c0�)L*�ӫ5�W�7���Ŵ��B�F0�Č���e [
�B�����_pש����+��Ed��\�>�	��ndǿ�(j ���B���j���2����m����j���|i�:�=�ֶ_s�Q�ȚT�j�+Ww���NE;r���C���&񻰟UO��B�u��;���E��?��^J.�ά��~��f4��s$[�]�پ��焬�p�6�EN@6ܝ! /���ĽS��P)i·�5o�Z�c�h�4�=�% �k�BE��2�̒�Vޣ/��$�o3Iq�G#�J	!t'pOD=+��z�b�>��-"���#���e_J!�F#C-�R��	�ROї���6�%����G�B�긗�LM����4~nP<)z�+?i�r'���eX,Y��x�T:(��)��9�����G��m1ܣ���(�aW�@*�hֳ���V��_UЭ[��I6�Q@�@e�j���@xK�L��]�JD<��ӄp�v(���ϱq��^��� e	R�
����2K�E$���1�]��S�*.xF��h�z�Ya�ַ�
�D�?ڒ`5��Nm���a�M5K����j��1ڑ9U����2W3����v^�l�)T�X���nO�k
���V��tpl��*����}ơ��GTI�w����mj�������$�̣��K1&9��^�0����O��r�����T�&O5Ϊ����lD��5�k������7��m�b�l�Ɓҗ����s���܉�mƩ٘� ��K���k���˅�(i�VFl1���ů��q`���gU}EUi��J���3܈%.n6(�`�a�B<F�S�,t���T�#����+G몁�h��`j5,��`)� ��7W�(Ֆ�+X�INl1��U�*�R�m�>��@49�t̑F�1�<�|v�����ۖ̅D;�¸qb^K3<���$R�;w}:�er��0�@%��d��w[���H1�#եf=%Ҳ���'�wI%���v!'"����ly���W� '���j=[m����r6P�[��8��5���ͦ�0��
�|�/�ig�Y\^��"�Q�e�3'�l����œ$,���w_}�1$�j�s�k���jT��$dx^�Q����hK'64�u	�X�<�*����?mZ�����A���msW��k�Ԧ����j"��.�}�x�iW�S��_�S�f_��A��?y}�@���,�u����-�}*���
[4�K,��n�E&���.A��8�iH�|5��溥��n��Y|{�Ԕ��=�x��2El>�A���3�H�r��w���C{��z�ŉ�xr�RT:��r\JM��'&I+\�0�K#t�����fa�,2�^Y�Q̶g��b��2�?�hN���+���ygf���h:�8a�����t���ƽ�τ���FCQR#��4w��3|��7:���,�b����Z�n	2�Ka��;�qw_ءf���dyWh�I(��������o�z�.߾tcmq�6b#�)6	^�<0����J�Ee�V�k�b�&��{�'�54�����r�&�	d\T�q|��7����P��F�q�G�%�=M���E���T�,�� �Ybg}ٝ�b�bs���I�4����e�_���\`���;�[�M�	���h��tڦX�G�&�,�ݱ4�P]ᴻ6���H��h��UsUN��}��<+gp���w���}��N���fu��&WƢ�=��z���(`�]���-�s��*�ro��Ē����u�Og_{�z��!u ����T��u�_�l��F��(�C�`�2<T�� ���.�����|Y��z����~�$A���>U<��[tS���;�h�\�,�S>�_�ӌ�(�����f?����;"4��p��HN8����P�j��..���pgO�d�G��Ҟ�"��T�NA�W���]��V�_�cb�j��s�r�6aZ־���'Q ��3J�w�A���ְ�,�ho���
T}#(M'M����hU�7��eُ�ά�(Eq��!�"��R��0o%�)Զ9���~Ż34��vů���s�;���B�@�|�tk�=�Rbk5�G��#z��T���cB0t{kH�
���wq����׊���^C�"76�q]��Z��~B�bt>���F��bk��U�����b�<�Lݍ9�Zq���މ.���S��	2�"<R_�RI
�H�M�q.e�+y4[��M}ݙ��c��~�l<�&�^��}\�5�w�g����T�g|�J*��n�������Fn�@^_2���	�~��T�W�\��[���zƲ���������W��G;�UtgO3<�KU�b��3!f����Ap\��]F!jF`�s}�o��?8�}�3�(1c=ﯵZ���r�Y���|0�֍����X=�YF;\w���D���Er�S�LH9W
��1�.��\`�q�`ze����M�\���OYcg�m�s%�K�o[�b��V���q�#ɧ8�V��#{�RI�q��R��w4��6}����r��
][�҃�[�Qɝ�2����Lr5U�*�&���a���ux�(!r�[��Py0�냏 �c��v�
<FM���b<�;�`1��]�������<����S��6�s���\Y�������Oe0��C��/� �yJU�4�~ٗ�ט�c��v�Y��-W��X"�A����#tT߷k/�z�1���;��;�k3����HJd���8�<��T(fg�7�h�P�%��M���ʁ�����)��G槹gx�=����V�����
�/��g~T(�P���	�캛1��}��	i��������H�{�i������@Y��7�S�3���lp�����t�%�AFF��*�S�j\{�ǩ��*�>�gX�U�e������ �KS�,!�<G�^'VM3%LlQ��d'Qu�UϚ%&sP�*�[\�@��h�U/��e�Pm1B�bɐ��D1���o����1n��f�5�ٞt�I,<��U��裏w(�dm���*cX�&��
F��l�4y4�r\6�aa���~���g���({ܘ
�!T��>���a��zC>�_�¶��{�s
6��h����{atL��i�ޜ���*��˰�[owLv��%�c@�e�|]�l��<�#'�膜ם�>`��.���r?�jM�Ir>��uk�PL�9���E7zu�{�Ʃ�T$1��4�m˪���vah��D�	'0�EcGemj����pb��I�`�|/����vG����o��a,=d�NN�ۧ�������0 [�p~�c~�+_�M6�G
k�>�|�~K�˝��ŕ���n�=��ƀ���l���o8���tO�!�s��I;�A�5�������#���ĉc�43)������62q�]��NZDT��ݼ���mh��X�v�M栏:;fB��:��Df�V0H	���k�r��9=�\�?�V<�j�MM;F�!����-�j�hu���@E��	ԲRxM��v����g	��R>X �����n���۷��f���f3Z�w���Px�YJג�u}�%�w����u�+���ǚ��S��n�v�n1���F�4r[M�q���0����7@h�%���
���s0yz�T���+	���X����t8�X��կ7�\s���(K>�z���A5؊h7��iR�\�&	2����>�n�YN�}�n_;C�ʫP���������*%Q��u$�=;UNU�D��#�{�ک���?o� �zQ6p���8
Z|�Xy=��C;��]�(��c�s��[�5.��v��v��ָ[Q�~��Oi��^g����%:� e�í�	0����dK�5WF��ˆ�����/���m?���hH�cM�������X���K6�z�)��9���vcԊ�X����ǰ@��<�h=7�1��z쨞�D8�.�(.
�ef�kej\h.�	T�n�������Ł�P� ��7ߑ�#(:�םe�Q4$ź����̥���~�#�a��x�5�����o�/X1Hu�>��"���d	�s��u��Z�U?.�	�yd�~˙��(��$Ã)k�I��ih�Ϥ�3�*��%E�P3������J���U�&���1�SC��reBϣR�˲��M�]���A#�ɍF3����������/4	Gt�m�g�y�w�/��V�v�a}�s8Tq��X �мk��;�M�&\/˦	mk�8으����&��%��������%����X���ǩ����'n�4��q��$�R���,=8�7�A*��P����5~*`I���J|��֟�PZ�^����e$YJ�S&�C��r|,���g���-�B�E��{�%S	�\�	�X�R��� h�ʲ�C�lx�s�p�'�0=�F8��|���G�OoO�f/ӽ朳����-*Ճ����d�򚹾��t)���t�qx/�P*�t�1�f�K(WV9��8��$�Oz{�k�=��Y�P�X��ku�P��c�f`�(y
&'[��F+�Oi�;���Ku���p�9#L@9�U{H��jM�}.�?��*���c�L{�n`��-��b�8�;��8uI������0!\�����(���"դ��:@S	��zJ瓊�)�<9��3���]ci��u뮞��ʎ�J��%e��!B <3�)��w�Ē���i�M�:�)�E��=�>��"�|0�g.�d��?�2t��T}�w(��fq""8ʋqy���	Z�xEKF�������nܓgJ��66@�,����/Eg4�g{)�hE�iHL���M��@��P�%�6}i�Զ�d04�94"�W&ɨ��hzܮ<��l4^�%^�l� Ep�Qܩ�s�2m�����fE0m�ݳ�Z�l�^W�!/�5xk>Һ���Q�֪���u>\��W������^��~o�]�3�g\�	��!���'�(L���B?o�aY�hܪo�׬<&�����UA���uB�d_��@�e��6�Mֆ![�$�M��y�w0��͹F-�DF�vJ&�&�Т��G�_:�?��$#mz]�B��LU�a��-�b�����:�#}j,�t��ul9���0*[�z�)����s�Rm:R�UnGB�!v�UO�)�sj�<��&J��.>#83�����V5�mA'��t���P@�݆����](=ɠ*��uX�@��#�f���b �����G_�Ք��*e��S�*�N))�����E�6�K���lɜ�������#G\��8�[�r����u�4B#�$�.j�M|��99d*��^���3 �YД�ʍ�����~��py\ȋ�~2S��E1�+eo&P-�q�G�@c�%<��F�,�/r��������B���d��gy��w�GmA��~��.��NG�=z����B-U���W��4(�۰���$tK��e�q�k�ǂe�����iܯ3W8����c� h��~��)y׺�,�$x\��h	e�Pn�\�y�ca�
?0��;���8���pU.�ZĀjN\4��h������`��d�D���lc�'�������Np JW)��r62{������I��"��FΑ���8��͈uт��@��.4�߁�CZ��~��$�[�K��"z���fQ4y�Ub�Z���}��2��뢃5�*Rm^	0c��b�-P'GQ���l��y�G�p�"��S������V���G%�s� �TQ�v��d��_�h���*�2������Aj?�\���Qd�yzT���#����8�."���t�֮coui�(�@S��1�"+���L5l�[n\�.6,�I��
U�=����ls�Y;>��j��߄enu᱖Q�Y��W<�rKz?2{u�:d�����Wm�_@�������b�&D.�R��}�w��h/-�u}�Z���s>^��n�,�ס�!+������iA���-�=
"�:����觌�<�
J��&�հͬ�Iiw�ψ)���bP�B�k-ŜO�a������)7�6�EkC/oz�x}V��r�f���5V��Mn�e����ӻ��|���\O{���c(ܹ��}�	<E��Vg��_cވ�(QL�lf�}��^�5�I�ր��b������o3����?�z�Pq�"��Y����t�b��	�N'e
��� �RV�ռ�Ҫ�5c͗�X�:���P�N�3�BLj�S�a�T4P-ݘVHr�o�V��X�Ӄ�H�X�"ƴ܈]���F{� �E����t��[v T��i4�Q7JS��	��H�U[�L-��!�X� ���z�Y�jD0�>���洀V��F����-��Q*Zߪ����4Rf�A�Z�\����|��:����%$@FHJ\Hg`��*�]Wp%�u�Gk�+������N� ���#*�I�8����K���m1v��O���n��N���zدx<UH�A�����L��d"�n�M��~�)]�����c�ѽ���/8���Z�8-��2XM��)�?�>���y�Z�"4.�؊���<�o*�薀\΋�mt��{�/���sˇ�p�m�'��iV�jH$u�n�]�̀���iN�����®����?ҵ��ٍ�K��w�:	�	]|�_�.-'
?FPˎV�<�`y#�۝���l5g��M�u5B�w���G�=2*�a\E��R��$�+��YO9��"�)Eu��/�v����_x���P>�$���4�}�����;Pq%���Y�5Xb��F�E����vod��B˒�G]���l��j��c�𐴫��S��e\0��O�:��]|L���f��������҄z��풣�,�j��m�
8ޚ�h��1�%6��M��w0U뇹�͒1��$>۾��Y�:�B����ě��f���Q�߯�޸Ft�9j��7�q�$�O� Ye�A��j����У�%�m�"�C]Y����G[�<�5z `�l��2�8B|�����F���xRr�c�/�W~�/�f%�2�zvW=�B�ڡ��t�мư�A�em?�WJ���Һזp�	��o	10�z2#Z��x`)�*�S֋,�CU(y�&�Ypt���}���>�-#�̛�qPڤD����A��6�:l�\�BG<lL�U�&3|�� W����<l∅��B�u"o#����?��M�3=����{Tٺ�� l�!&HM��3L酕!ؼ�Ь/Gr���I��'���L��R��g.0�}7�y8t�=���񠤢x�D�L?�q�U3M���Ik|H�R�揢�tC���W��2��Y*7�op��^juJ�p��(���%��n�DZ����W��$�D�V�e���[���H0�r��#��K;�\��-��R5ΒD/���J*p���>��n۝�D'����v�l�ua�ޙ�����&Smj�D,v?�'�g���ʼ���.�'�A���{;�9�+�Z)+�F���R���)]�'_YK�9�e��z8-!��T�`!Od��X�<~;e`E2�nL�_S��+��;���v�Q�͎���S�N�e�����`� 'Z���J]9��0"a��_�{��i�;`�YP�x%�=ɵ׈�Lk�}�G�ROo��}E�(�kz�g�uF���eS������6������Q�?&��&�ˊ.b����E�2�������&Y�_M���z"kت�}��H�h�������=3�K>����(�v�9������˷�m�M�L���>�޳_,�Wk�~��NF�C�+�CD���������ETo�ÜY_ov��&��(�<r�l��Dk ���a.������� ���
m��r�U��d�R2�^MO	��E1�q\y�Y�h{y�	�7%�T��w�H����=�~�ZO�l ��-�7Dq�+�v�]}�А�ǉ���� I�25a�71 �?�
�������޳���T�R^����^�(�9��W�&<Gc((��4�j��Z&��A�GL�08��螸u5�o��N�	F�)zN��\lG
��	���;8�M�s���_vl~nw��&��h�($���x�x�[���UN�̧F��y�P�<��/����%��$�U���_^�(k�e�ʔ��S>�#�b"W�Q�fp�*�1�X�kU���8)A0Ȧ�E���Q��U0;��cඛ�Z�OZ��uC��I��y����ER�Z�z�o��<�A���;�<��ܼᏍ����f6�,B�����rJ�B3�~qIP|���fz�BNw3�\$��&�c<ݬ�Yoz��r"࿗&0���W<ti�C�x+��N?4�4:�(�\ ������Is�f�ԣ��ǖ�X�ꆞ�X��NO���^�1 �AA�@�l�4� Q�l0G�g����v���W�y��?k̈vӂ���i��B?NB�Z�=\��n	ch��S��[�����HD�s�F"��.#��*�tv�BN��/H�&u��d��D��3�tH�������W���P�Q
}�c���2Wj-
s
�'�L�����<���-�	�(>��U��- �|��t�������NP��J�a�O|��PC�Vb6���U���y6gw�%J\��LP�3�����	�I��i�X��KmC �c�-�+��)��?
���}�h���i9!��U�o�aSw�G���(�ĩ���ޢ��gE�܅�HL5s2G6�Y��HyO���k�Gx�vȮGs��)�;=k%��@LK$:p�]�XZ�$c�}4��|X1�W��_�����|;�`w�.�fӵ�� t*��Ͽ��ܛ*��r�tt`�"=��5�����s�rR�w����ۅ�[{��B��:�d��w3��� 1�r����J���� s��rP�k����&����Z~*�����	�����q�.P�0(-1���ݺ�b�f4x��?�P��=������P{vn��w=*]χ����&+�h�{Y�BH�}�&gF2ّQ��&����l���be):��f,f�q����R*L���A�Ӌq�c�9�vs��+�.�)�&h�0�.���#+�4��R�� �H�*�C�����
��Ԓ��Ӕ������˝<���X�'�ɺ�Q�F_Or"��f�0$����k��	\H������hZ�x5�d�h�5�57��.F[�~�e��� �Q���<�͈�ܦ������*4�݁�X�p��-i�QG	W���m��iJ1�ȖT�� }�ɿ*�[[�ߝr��D��3�f	?��s�#�_>5�7��]����R������+�BtYiV1�n7�˧�/�.�+�8�7���Y�H8�ȵ���d�7�@������� �s]�q�,4u'攠��>�v�=b#p�h�_>-�,e�7*�A�Yq`z�>ov�~��ӻ�:4u��6
bulv�-�V���%}��s ,Ӊy��m�qT�S҅���.{(4'M, ?-�3�c%��"S��iI��k'�/v���$��|���6̝O��캘Ӊ�a|�Y�l!��c�x�j
��
DGi&ߡK�i�k�y�(BaS��=Ql
o���5�;��&G�b�M��Q$�ڸD	�ɦ궐e5m&��S�,Js�q����q2����A��R�FŃ��z̏���N�Q��t&�����C��D�ڑ'��B9��47����Tw�-��o��� ����q�t{����ܾ8�\�}]AqŇ�H�B��P��~.D�	��Զ8���k��X���������q���2{�U{���������Y9^Sr��I��q�Gӣ#�ެ*�e��U��w6)��28[@�a���'��d�H�&t@��'���g\k�O�\��Q� �u6�7)P�փ�S��W�m�#�mû<  \�x��Kb������,G��lI���F�����/$�,}M1� �mr�c~�_�[o����6�)`�l`�]m�Ǳ������R����98K��v`��8W�:e���h�J.[K�P�HB5��D�k��$)����$i[@�"���:��i�)R��e����e��|L�����O��������ɽ��R'�A��Y���J�:���A���������߰A��Z$�z�Ye$��aQ���� f�ˉ�VW\:��qP~����'Ȇm-;���ک��:��\6�G֪��k�K��[~�e�/��jɨ��+��>_��g���������~᦭%�Ҫ�b�`��!�c�n���(�~o˵	�]�U��;�.��k"	�8z8j�v7W���3�i�j/UO#w���ߔPg����L�p�����+��И��mߓB~(B̡:gG�q��<�e��e�Z��y>�x��i�ue��>;�0��t�^1K
O�Cy��r֯
���{���:�6�'�D͢��V��a����,)�f�L�tW&XV	�@qH���59ra���6D�7A+����H��:#��`?T��A�l�1]<:|�]�)��j,�G4�tTx_����vz�I},KZbs�~�G0���/�u��R�sI�j,���W��qJT(���D+=��H�P�����.R�L�{@�8&R%0�t�d��@ U/����+���������C8���Y�P�&Q2���|n��@�͌m�E�k>��2�h��L%M�[���4z��*⾄<��o?��D,��1d˒��[�~���.�^���gҢ��Г7�E�J;8��X����K�=�� ��w]�`�[o���r%�#�AJ���B5|x�o�mJ�~��XV�����m[�K<,;����(�n���JǙϹ���2�4�S��
�+VoHR�6�Ȟ8G�,��,&J8v�*1����-���Q���0#L��:�-� �*a�W�aqerpz�g��Uas�mh$���u�hQZ��o��ȕrkCœz	��m�'"p�������ːͿ�?�E��Nq�C�g��I�����bRH����|ԉl�V�a�H1��b����ᘀ�$�;���s��'@Zm	=�V�oc��_S��Z�����,4S��a�H	t��叁6YuV��Gt�N�$Փ\���������O�x#T��!�iM��OG=Wgcp��+�a�ޢ ߤ�f�4,R~��t
�T�E�@��ad����o!.�\�|^H��P9h�r��~���a#�f���A��{�E��������-�-K"�k�|M�grⅸVpu�#r��8�r�e{�r�-� -�<�Qr�A?��Iv�gtx��8�V] �>s���Z?d�E2_�05�7�Z�
Z�ӡ�B��b�SXt{�+�lcUܕ(�EV��ʢ�E1x�d̸���kL
!Y�x%`�i�SЄw�Qp-��U�a68�mS��zi�~Ba;��@���{��anø(�q�}�{:�1��ڧ�x�m�2�1����#׃=��C�2���?�<z)'�o��'s5EUD�h�s!�A;op���[VH��2<��?,���N�wȌ�����)1�y�;AAw#1H�"�;{���#4�t�2=2����T���8�A@ ��U�8@]�謔���%q�&�9��ސ<[���)�.�R	 �/�h��F�Ǆ�17(0�����H�U�`�$�݊�ݱ��l�uV�U��g~%C�p����V򵺑�%�7����U�L5Mk�H��V�F��emGj�~���*UAk�.�-z!��2gExx��0	W�S�$ߘƺKyC	��n�rMLdcz�T��\J��w'�H��|�?��/�DRo2��#�Q�N���j�\��u�I`f���a�1����Ҽē�5u	N�������ء��Oj>C�p$�>��7���=�W��)�-�VUo)�D�Z#�o
N���stgS슴t�j�62���*#W����X�m��7HV����]���_�Z"��7��,�E�~�����wE_r�MZa�^p��B)zn�O���U��#!��BI��GgSS�p"�ߚ����:3��`��m�g���b&�`�-`�z5��8��c����6r��.�V������g�s6w[w;��E@o2�����F�n6��L!��Nؙ��n�O}��>F�U��~.i&�d����w1&��-��vo�NHIv�D���c`��6�E�_&�]z�\
Wb�@�VN��b��OC(���Ч.<)k]���q����7�#u;C(E?��C�cq��F�@x|:�	�� E@?�!�Wa�afȀ�c̯	��}XАI��߃;8�����z�Xa?����h�5P\y���S��7�a�UDDq��
+����ϰ.m�ʫIE���?�P!V�R���[7j0��c��Tɸ�&�X�}��|����� e���1$����S����b���'�Wh�S΁�d= CUG82wP o�O�(<�B��L�}(�#�=�C�Ոv#O�|N�z��#�Qt��v[s��A5� �9��sz�&UX�{S�*c��}��`���?��l���2;����2^�{�:�θ�X�=��;r��GtZmm:�l���NV�u���n�ݒ��D��yPZ��Խ*��w��:�Qor]]ʚ��lt�l����5�JL������o��S�&��y�m�\�Rc$�w���\	�츯�*R��xf�u�Qn��I��C��L���Ք�Xߓ��!�vr=��n_���u��o�+�W#u�l���\+�ZEf�C!l'0"8�w׫�Ҧ<&�����:k�BA��mg����|^2x��Y��J�rű0'�0/��`�'�Ζ�O}�O��m��� ��<"<����&9,�����D�Mj K�t����կ���A�u��Co��s�7HY�y�d%�� �$��L�7�9��\/��w�	=c3׬x���	��к�{�4yHEr�@��S�g+pA��\R�k��q��d�lD%i����vGl����� @�`Y�#�uP��,�	�]]��8�L�(Ql�ӽ
^W��f9�:*��
ɳj�?ϯ�8�� g�٬NH�:Ń[*�搾eq���M�Q��ͤ���l"6���׌�_*����4ss�1j�6�x!i�C��0�|�[��S��r������=BwX�T%� +:3�� 6�ٳ������kd�Z���B��g��Bd��3>7��+2_g�lf��i*��Aw�o�
}+mA>�0>3]w �]�a|{1�*K�H1�8���	u�Z3�5��)1^��nA6�Ş�)�ʻ.�#�ǥ�6«�s����~��� ��s�Zv�����||��~K�N�؟=����G�K�L�����#[p����LL��sk�Ae���'%����5�b�*[����p���|�}e�.Yp�R'�/wb �����0W�L[!;���mM5�᭸&�h�����x��K�1���;�-�W��wP�Q��X@��t��pzb�it�񪯼�$xY��7���Ec�3ޖv��)[Q���5���~J����&�E���J�
ymP���e���6.7=�����p�m��:8��F/p��z�]����A��� �9����=d�A��R	g�q#I��6�3�3����4���f��|�bu���6^VȄ·�R�����>F q �ȌV��J�4T$1bm���7CW�CUyC�hm[����"@��p�b�3W:�+���/�n��R'JNGO����ƪ�^JZ�	F��J��Bv{���*Ƞ�B}�U:�b]�wD	�Mh��Gm\s%���A���$b�;7��"N�5��#�T�#����I�N.�l܎��t9"t����� E��zԐ�_M7d����t��PF]�w�r}KӜN����Y���C^�C��y"HBQ�e�����΃K��"Tp�C��2�ҡ�����lj|`w/p��fj#��?��F�� k�������;f��573I#}úQ�@)�2?7�4�L�,\T��9EJZ��ݝP���3/�$��O��Uq�c���;`��/Z�tm��{4$�,�a#Ag��'�(B�X���{��f^�.�~��YW�)��n�@Nr�`oTv�V3kA{Gz��Q��2>s��q N�^5��Ƅ��|��Zg]\):�1�Z�0�C0�a.�e�d΍#J�:��hn�l�.����xc�?�S�E��ׇ�T�YO����o��v�[`�-�AT���=�=�z5��̚D
�kf�~���0�u���!���\�Yz"Hgl/t<�ADAl����4�@�N��3R��P��	7C�;*�`�S������Y��a�)��hI����[	�	����ҌS��-S�I��p���E�a^�P߶Ä!��R�ہ��ӊ�d#JR�ei�B<�0�c�>M��w`�!��_Z]IJ`tz--
���vr�q��"��K�Wv�j�:��+K�v�b~��aR?�lkn���|�T.#@�'�8��gN��^sףmp�8�Դ�����=iP(k3�r{Ͷ��v�S2����d�Z�ڳL�j>�v��&H��tY�p�K;�.�׵��S�8����F��`$� (����>���O9�+a��`p�I[Ǆ��n1���^@J8is�`�� �QQ��Q�e?�_}ۀ��-�����@��Y�L;�����f]S�d$�}���+�J�a6�¾����.E�3Z�`�L����d`u[t|��,ɷ[��UJ�YH��* t��BeS���4�w���<?��Q�}޿Qy��__+��=J@��ރ�e��m	O{j�`��i��=����h��S`��Wq��`�3X�F�î�@�S�*}�L��Z~c@J7�I���񖀹�W�8J�C2x��o?A��I%�I�TiD��4H12�j���+=�@rq݀)�ʜ�L�d�C�� ^��ZMf��G8�0Y<�sM䤁�.�J�}�)��xG��q��T˹�l�c�ς xn��0�I����l���NV&[�??}�W��Y���;�_�kQ,Q�ma<A����3;�lIvz8"�Ĝ-;(�py_�_ ń�����>O�$&�~�p��4�S�=���hM~≍�+EX�n!u/�v��{��8���n���Э����?�~1͂�y��8/�����8ى��	�Z%�}ҁt��wQ�Ґ/�Ut��sbim��~M�����kP�� ��R��BJ�γ��%!�/�젯�,�?ӗ�������nIl���h�t�/�]��p�j�������qJ�jE��N�x펛g]�P�^	M��)-K��}��{sv$��V�Y7��z���b� ]��z�@8>��������9����C��bb�Q�4$��e�Úz�Y(�T�#h�@����xUp�Փ����Й���_��+ν�nT}���v�a
�Y~��Z(
�0VF�{# �C����r��JY݄�*�o ��ؕNF9��D:�����C�pOb�a�4�b�XŇX��SR��FO�(�4	~{�Q����6[���~v�'�?N�$���bz�~U�τ��)������Y�I`c��l	F�˭�f�~�N�w+q<��J���0��W�y�7J��zg�WA~��p���D�>��˗��«�J;Gɽ�jg{ʘ��_�J�p����;��u��0ɠi\@��9h�x��~+t�;�+�1�uܩ.����(������>Dc�T���0�Fo���'�c�5��un8T��a�#{��d�z���2�'U2���6f�:���X3P�6�(��T��i�8gUj�o��BEMz��m�ӹG)����_xq񯏿�T��v: S���t8@Y�o�D�˩�)@'��DT�u�oC6�V$%�r�`�Ũ���Z�ѧJ�y���%�[�kT!��sh(�8!���� d�UL^�G�Աn�q)?q@�ͨ�!bq��V�cE|Vr�����a���VJ}t��lEb�Ul��F[��~� ��ò���&x3�x�0�WJ>�o�[�e1�.�7͗܃�*����:=�uΏ&Ɨ,1kð��.��E����_��3���Ň�n&��G{i򱛴��o}|�������)-��_�A.2�dq@�91��@�g͙ pr���fm�HY��~{��vb����g�%`D�B-���"�LA�:�߸e^�����fisw���3���{����c���C�8�6zbWD�/�d��m`*��[�pߛ�r�i��Ϭ>��g�8U�f��|��ߪ.LҿT|\V�*3a�žA�!z3.U�8˼����<p�/�;Z�l���ӑt��A�~��;	6s�X?]�`y�3�i��������Q�W�fGt1D���gE_�_��J���K:h���h#x��!�?9�נ�&o��̓k�J�[������U�������Y�p��*	�])����0���n�-�:YK�4E#��"\a���'�O�S���c3�,�sگ�`ֿ���/smM�.Cђ��~������Ά�ﭪ���%�G�R�#�^2��u�-�#1b�hQ������)�z��@�[�ɩ �|��"��k�B�?\�x,�nӊ4����0���DH����Ʊ�dϭ�j\]��v�^h