��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6b�$�p��=a�7�-�kd9I��x804,�f�� <Q}k�CD�4A8vN4�'�
�
j
����b��!e�q�l���ub3�ڄ�_�:��eF��U�0Gx����'o.�
�Hl����z�$��K8|�Ex��]�C%�1��h5���L9M�NG�t���7|��_ 2=���[�&H�N��fy�_
��� ���W	�ęG@�V����s��ZǾ��XG���Q#!���i����|@���v�pX6>��;�����V&���o����&���]�����w?q-E*��s41	d�W����b�h���S�r�y���4�����y�6�w-��醢q�fx7S�� P?$�`*���Z���Ӥ��ǚ�ߝ�v�}�Y?�O5#�����V8mn��"�4ׁdY��j���I�+ڥX.f�C�%���(� ܽr�\��=y�O��Da������s���� ��]��|׬3Yp���
 ���y��a��	�~r��f��.�[ω��&$��>Y�Cr���ٟ!F�3�Ĝ�zd�H�k@��`ɤ�3�x�}^S��2+��7�+��Ϟ��[O$��Y�;���AF�jV�G���)�,��e�):Т��Z�j�ǡ�Q?ke�$�=`Qm�!��P8i�vj��c%W���[T!���dpνBv�w�c�U����<ǣ�H�ao�$J�>Ir�dv\��$ߌ$�8zV u�g�$O-DKVv&���e��>p?�=�XH����5Ks�P.�Z�`���:��TL�?X/��c)ם*˰�<ƜR��X�"��p�kk����\�54Ue¥a��;��`Km�6H^��2�M�&�*��{Fߡ�JG*O���$�p���k�ޣ��Vk�X�b�c�G��QT �/'��ȴ���X,%���5�6�=���M��s;���D�Ǧ��S0���G�n��W�A�spa�frW��C>b]|�,��=6	Qi��G΅:v�r��E�PQ�g�Y[J�~B�-�*���ٱ̅��,�}�E����.�����X��8����[��q�:yt�7�Pxt5��9o=������0+Wby����U�y?��_h�o}��R�Q�������Q��ҋ��v+���$�3qvJ�v.����n���6y5
�Sw&lw�zz�`z��y��Q)�ZG.�����i����@�H^�O%�&�*�#�ɉ8���u\C��eǭ����yC��?k�덫Se/C��9GF�G�󆾐�L�:�3m"��xf�q����&�@���>zj�A�!.����Vnh�����X�-��.�|��"~D���s����Yۈ,;ULߢ%H8_����$g��T����Wȡc��u�>�ժ՜cp3����݈��ߎ�] ��K-λo
v�T�&d7VDY¡B�n�ݺ5�UM%zKx������m� �m���� Al�L�5S:4�Q��tS�Nf��R"C��R-�y�zj�sIޙ��Jy2��ā�C��ҏ�����x>��c�շ+݈��
PC��c�&Z/ǟ|b���������Em��O5���j`�z�j6"�N�h2h(r���Lb�*��nq��$!�rCT�Ask/�m�Ѳ&�%�䰝�e�3����|��"�_�������KC��A�qq{1kp�<�Atj��:[�T||*y�R�b���	����K�}����`�a������iƒ��8��zJ�	OxԾ�?�*�("wpv���B�g
�@�����`|�æ�F.b��@s\��C%şP\�c:|�x���<Բ�zPނߚx�p8���_��?��x�o�#�׷R(�3uc0Pf��s�rbag{P�w��ٟK��K�n�YA�{K��(��gV��ɿ�K	3��`����e���$��#�����e����$��e���S��m8�
����F�m�w�p�m,KŞ��2�W!'���@�B=<o�:g�F��D7?~D��做qGB1G\�n�{�l�ճ7�Lԫ�-c�T ��6�߀�d�N�/�A.��/��'����1&�^O����P̷ꗨQ��ZQ7%�x�K���]\wU>��t���-@?�Vr�L�`�aBC���2I�6���Z���'��@�zf��8yk�f��_��	 t`o��:g�*]��(;VJe�c4q	�3��`��ʍb�N�+H�{����O��{swٓ����,8ߔ�
�
OW쵈�w�݅��.,�:�4���t:�-�6�cm������-��6 9�U�®U]^ʥ׾�q��<[5�G����~5_�%�<ʺ�����Ǌ}�w��|���T�!�1d�E¨�,�Ԕ�@�/�/���E� 1�K<�\��0�!��Dv6���̈���4y�+s�R?��QE`�5
b�c�	��眔�>V^�F^]bPq6�8�]��h���kllS*���
�������_�f�&(�K2| ��=�9 �DǢ1�<8ذ�Y�}
�w.�*�W�o���0q���Ӎ�kO^���1}V�̾���7O3I
����`\�)Dsd��V�71��➕�CO���;[��E�ed}[�$)��Iu]���}Ƣ��SG�$�;Q� ˿f��A�8G��8�\�l�p��a���G]z�Bu��/s���\x�N�asL*M䘙Db=z3�Q�jpp]�>�4�ǒ�kS0������VT�-.��L��>���R'>V\�	v4��[c̓�� ��E�x��W�
��D��H�Ss]�y��3��E�����a�e>�&�i�SI��4�ᑝ��7���,`�	{��*���0@�+�W5o�r'���N�����6yA#sBl�v+T(�.����O�Q�[8���>���4�U���xS��L�A�"�&�2��Z�"}
/��(�l�����WFP�˔(z%���N��,���K"���K�FpԆ�N��xs�n��`��0�>߼@�={�v./�u��$b���k��ӵ�8�8�����|��yg��Ļԯ����?���a�m��?��h�S��TA����!kG0�P�79J���;�,�gM��v��?��-I+�i�������8*�>>� iOAe�kX����<���f.�蝜ML �>�M)��+�+�-�3p2,9��
7�5�Ac�I ��y��#|�e���Ӕ�`w��d�9�&#ͼ�FI�2[-�^Jx�����EW��`�*����Q�#���GEk��bg/@�<��,�h�$�4T��ϒ�!�ۆr���Z:.ޠ�ĭ8����@�����+/���i�~�?$Ui�#�5l!��<�Ñ��� }�9��G<O	���麟��y��=�yz~�k̅���X`d��i���j%ed�:��O�Ǥ&����FN|��v���*�
�L�dU5��s�US�L��D���A�/[7bH��riԄ6 }B��[��#0�ZK��) 'h���(�WZM"�E���~����>�*��nF`����7�������: ���t���Y04Δ��:mR��6���6lKG��D���4�D�����O�sM��RD�M�����fPc�2��=Q]��Q���Z�X�̭�@&LQ�S�0���|�z��'o���*��g�7�{]�//f[;q9�s]���(S	viJ�c^�wws��{��-�v!��\Z�|O��O:,p���3V0�mo��(��)���8�Iv�;Y�T��!A;�I�8��<	Fz�	�bӤ�8�[�d_(���8���Ɯ��u}'K��G��`�8��t*���4�(��Y�`t»�ç�RGRK�ص����<j�?�3 ��ÿ����K�/������\\s�;>:���o@�c-����"�pW�v_�m�$1G�sURt��ɯ_�G�4c|C"Ί��3���b[��>b��'ʠ��+0Ȇ:�I���w
"��[�.�[)�P����� +Љ�R�h5� 6x��59��^��7��2�Һ�XS��!�r�_I��i����"ܫc���(pSQ����\�:��2�4/qG�֩Ch����:T�fg)H���cBRڊr��3�=��r �>�������ڱyK���$���03r����C?h�F�br��A�}�]q%��t�s��y4�
&͑P.�8�"կ��i�y�j����>�/&U='��HQ�z7��2L!��ugI4��]��]��`NY�������ia�8*��#�����(et�L���FF���D
Ժ(W�P�<Xt�ur�HϴG���A{ޜa�#����^
S�o��e�J��"UT��ݫr��_�9���J�;w���,W�`�O�z$T%"�"m��ܧuQaS���^�xА�����!/��&:KVJ;���u���Zy�d0�P��PD�Bm-���O�߼P��a�>D>��{ �8T2#Kl9"i�G���
8��Ad����e`X���/��J=ŭo�'uvcg'�)�a�]���t�uB8�Y�B@����9i���'JQ+D׾�ՙN�6��;���"N�A⳯��/�)�.w�����zθ���a`k�G�0� woٕ�D��1ҳD��"H�;�R	"0jx˯�R��[e�x�1�;��i@�M�ΆY�}_}Ľ���!�P�kB�
#o�
����đ�����7B��;���nIz�H��r���a�RƼN�����J�e�a�bx���sF�W�pW�r�K�����#w/Y��=gѧ̺�w�0����A,���1�-�5a彾�~'x���}�"k�/j?�����&�����}ޓv#,C��9ǜ��J�@	~�V��8�r��^�{�L�d^����>�f���l=}�=�*�Z.ZBʹu��9]}�[�+&���� %�{<<�?f�,�&*�yzA
���( �DgQ^*zJp�x�1(tP�7ơ��n̓��Y:wu	O�TO�5�X�Ѐ����Owb�1z��ַ���딐e��*XOψ,�ie{1p�E���][�F���n<����O�QB�W=JQ��IJ����ϟi��߸Ϻ���+8�=ixFf�!\��5�q�SD͛4��w
2u���1����H�$juᙡ���L�p�"#��#�J�0�u�Uk���;?�h�2���^��2`OBkfD.|��x&�Oyu��&�֔�A�Ю��B|Ǫ�@��Y�=[�1�i��'m�e�4��?��T'b�\[;qb�x(db)LZ(��i� ������|����ԟt�kX|"D�?`�|���E^���(�xla��L�@��6�����q��7��WJk�֐�1h<��ս��4>|bs��n��� 'r6D1�T�G�BFR"d�Y+�V��|kTyN�Z␴���'f���Zk�m�O�,B��xl��Y�]L%v�|\ٍ���>A�r�s�0(���ёN�S$��*ҥ%���s���u��nx��P1�% ^^y�2GH�*b��W���y���ю>ms!H�+�N��9t*f��-B<Հ�a6ӱ�b�B�_:����'��������hZ2�/��Sx�0<P���9.���������ޛƞP6����Z�b���{����Q�6��ˑS�X8QS�;6��v������F5r�S٨7�[���<��4������ly�7{LE0t"�W��ۉ�AU��Vm4�p�4�V�1�� ��.�G̳���F)����;S�q���&��o�>������E5����f(�nG�~7�\G����QHB���q��$.�ZYP�{o--<�d�m=�Ӵ��͍��3L%�'�Uݱ0�<����X��g ��"�_~I�G=��q����.����2,E!��U�{��fF)�dHג[l���Dy帟ʈ�V��>{�U��Kz۪H�������<D�Lu[��@�)oP8���p��B}ц��6����iU`��4��޾�}�/��{ލF$F���.��JS�m^�Ҟ��m�~J$}вym�/�)�#�#��n�@.�=�ן@�d���*��(%�|x���'ߦ��J�s{sK8z����wd������[��1%��ۭZ��j�6F~�l�|p�pN�����~���
vZ�]%����7ZQV&�'SuQVo�=�L����s����괐��{oG��	1Pu2��!��E9�aO
�9���|N�Z�扅i��P=k�D�J(���C���q�
�\�� �E���=�}���Ѫ�r�^�!�������4aJ��n�a��=�/"�vhB3����1��m>���!�V��B���	�����7u5:�DXv���p��͋[Y@ioM)lM ����oa�d�급Y�TЈ�o�Wy����a8C%�A����W�L	���'^$�e%�#�*
��p���?2��	y�@�Z:�ǧ"-������8�ݵ��擷{? -$��]@P�ű�e��208�+���Ϧ�p�!p���zC3ݐ�<�\����y�?a��&Id�kҤ55P�o?AD�\g����AQ�Bc�A���,�$��.����
�Ͻ!�C�2�X��Wl�$�@'�E��j;�$�	`a�#7�s"a�d��O�KS�E�U_;����W��$@Ɔt) 衏b�β�Rb�G@ܩ[�@� �q��H��O��F·�"Kp{����]�a�f���������1P������`��B�ALH�"IT��&����,Li����q�NP�|��
#;�Ak�ĶN  �<F;��#�Ê�Ć���ψ�,���mo�;�� ��*�3C��R��ٰ��f����@ z���tB�Rt���^jG�VY�ҨO��[=�<�'J�#��ߊ�P�����UG-��n��r�wc���?�����uO�6�`�d�8�?�;�R|�y����绽� !�T#燗��rϓ_F���дN�e���V�a�����D��1�;�"��*B����R�X
�X�l5����)�peB�H�ݜC��3�Σ���?f����]א�#�7���J���vn%W�q4��|�`,#��jcdE�^Qz�X����?!{��C�����e�`uD�x\�����kY��V�$���ڣh$��D̛]R�)��N���������׆+1u�<�QS����^`���Ͷ7p�������eU�S����`��gf����=��J�j ���f띙��=^;-+�`�(_T}����J�g�<�5�3F�8�O{X�eA\�p����p�f�Yޝg�b%�c��Y�Nf^g���Xp4��m�V����Ώ�\�k�mE8�U#@�;F'4w�ҳ��2O�|�"�	��5�����l��|����4v@H]8��{����� Gb�â�2�uP�)G0[� 	��XHa�~��,]�����|��!Z�&�:J3�)�[�X����c�>2�'���ԓh�F��i�"(vqӀ��E[~u�"���1����h3�p�!G	��X�I�����q���:����3��ӣ�����j@�M���dw;eg��@�jH����q�������v3��+��~e�gpW��.Ĭq�Ca��|��[ca�Mp�ď��lXcj�;K�����o93�w��O�k"�!�YH&�٧�24��Mf���,!߉�"q��om�o��[����:�u��%�x1���c��p_�p�8W��كƸ,kx����zs��~��?���Pg m����F�¬�ys��k�:���CC�I��?�*�S�̽{~�U2Y���n*�/�Nϥ�,���J�rF>(���`�:���R}1fR:22��"�ړ7��3�`>90��SW6?�S;Ⱦ��d��1F�F�A6����������)�D(m�5���y|�`�l<�'�0�)����+��[�?R,+i8�*�%z��N	�c4���mA!�bK@�qQ�؃�A	��j���/���N5��gR1��^��7pb_�$�o�µ�����Q�%��T��=�?��lL�g8
����oa\;"vE��[h�ݔ#�5�n��Q�"�Ch�砡O������:�L$-�ƪW�a�v���$d����;�����핾L�Ȏ���yVC�<�AAv��?���9�a���GR��'<���2G���o��>��?����ڛȸ��ǃ��>�f�4�v���-JY��I D&;��{{`�>��tLT[��_=u���Z�(g����\�h���{�fJ��ƻ���cCϟ�τ+f��?�0Y��\L<�,�-x]����ِ���n�H�T���|C�b��w�N�m������:�)��SXD?�_[�$����<D�?�ဩ.�����5���	�>�,<&��@�G�)�<�Q�r�~�e���t�f�C0�+5���\i�B�GJH/Ṃm6�
�Y��|ގP��?͗�Q��YT@�ߙ#���%�S�CH)�C2��3u q�4yÖu��F)��3���`�料Ї�P��t��]��*�T�%�::o[v !���FE���
I2u��/�UG�������IS�~WI3@��S�s�}�l�o�1��.Yl%���0a��k�)sbe�<�Q},��]�Θ��JM�q%H�#FY�&���3�`=Ӵ��S��v��6+���Ӽ7Z�׹"`9-J�WތJ�H�9Sԙ��>E&n���EPRF���!��s 	��Fx�b";i�R�����m��<��|�����.ز�:��%B����В�ܝ��P:�5v���֯d+����J� 0�.�DgL`�Y2E�߭��DDb�]���	�*�,ZyP�wʚy��j	l��E�~�R�����Nz ձ�"z�����L8�9�R���&��K��xJw[C��`�{�>��pO~xC�7�S^;�bM'�h�/�[[�ќU�HqM��c���;+�j��|y�0}�؇���2�+m�mJ�h*���I3���x��s�D�F��AU�o �= }�o)��W�Yb�g��N)]��u���"��h���/p�����{[?] yYB-+� �����F��/�t�P�������8O��p��>m)�2o�ȥ�R9+L]�s[�E����%*�+�w�a��V�;���U[4��N���I��c�8�0_��Fu�E��{d�ț�#�����4����ɥA.��mBu,��������s�ߛ��!I�H��Z�s�� W���������I���Ƚ5�B�6��������%8��k���w�V"�HL��B��� >��/ǌv}��Ő��+�`�V��B7�V��=���2�d�(>�>��ӧ�KDL.���}��n�Ф�P�Tn������;�����6w���ٛ���f��*X�͊D��'�`Rأ|�Z c5�u]�"�\��t!,�{4���� ˁ)sd3����B�&����@\�2�RS2�����g*�7�/�T�p(�{`�a�����A����'��m�!��ǂ��G޺,_���AN$^�[�5:����D��8����Pɻ�ͩD�RHzm٨��ޥP�2�7�ƌ�ޕ�-�i��P����7���@��~��_�8�_Znj
In�Y�VE,W9�g^'8a���a��3[�WN<����F���#b\W&����s�&��q�xr���>��(~�ZH㷋�94Ĩ�]����_S��\8���-�V�J�x�}��4���'e�֏��)e��K��G���U�3Xy;���'�d�� �2���O�5�� ;Q�������P��_��	T�� %)UU�s�TW� #��Z�e�'�2�͉2Qq���;߼\ý�T�biazƘ@��~&3T �a|����s��3�M���n[�㉞����_���xԽ(o�r���1���7fU�(�f�&~�=����,ZR� A�T	 ��zx-�>U3��H�H��\�%T%fn�F���q�ة8L�3Fm�Y��T����:����	�3���� �N綮��t�S�v��foi\�[�'4�c�H��У��J���6}`���1���\�o4��֫JP%�^��,B��<��oSqA��B�?"F���;�
���^��OjXȚ��4%n�Py�XB��2o��[�����4��L{�d�D���"-5A�z�+�RV����q��~��.�'��n�݁���r��I$�B��H&E��i��<W���맩�j�')�j�\x7���S���ƃ� _Z������.�ȓ�k�(��o�b�H�ܖ��wP��_��;���f�ڰZ���1�[��_b%ȇ��ǑG\`Fp��'6�v~(�!���c�hR�㙀o��j���֯��](�#�ڃ���Q�uT ��^��eʣ\����HGb�c���糔nؼ������M�i�ƥ =�P�0��sf�=��� va�N�zӌ'Ϋj���Un�ӭ�2�X^� e��ϥz��I_6^�f�o&]z��B�';	�:^H���uƵ��أ�Ѳs�b��V�9D�i���w�h�*[��P�>:�H:�H�*VZ�Tk��>���O����I�ި��G!�4q��-�{i7x��}N��,){��Qٞ��l��R���35�i�c㉧��2 چ���#D>����R�3�skG��^F��Ƨ�4h-�S��z~�.3�|�(�g�¨ ��^;>�s}Vj�	X�/Wr6�[Q���9"�.pD� m�YtmlU����ZHl�?5~�H������>�B�\e���<��������q�8��
G�Z�dȇc[�	z�<��XmQ�G��n��P�w)+s3p�V���R����fS�J��
ZJ2�c�J�
>S]2�˛�]�J��2���w!b�ϼ�&vZ��ƼvY���5W�?�IJ�|^�<Eb��)˖.y�n~Thb���F4����yFm�����J�����!�?���f��.�u�$��i;3��T\ ��Y�>�P'�>�	�.$֔�f�JӫF� #��e�8����i���u�P��� d������:��;�eb�g�,Y���C�7	z�tr4�gq�b�{n�N��T�0�:zxh��Qa�b෨[�o�N�x��va�����!��5���c �A/V$�o
��\�/��G_4YSt��x��Eեa�(�G9���s�.Dw'�k(;#�?�7lzMV��x��%��t?���?�K.	��0"��y��I�O�7�QB�
=AE_�]pڙ�� fe�Q4�����WS����qBs\��pi�K����Kt��p�j�b��q�U�Af�	\��1�S>��>�n���f�	�M`3ҕ!u
?[�_%�1�Ի=<}A���)�H���Qy�3�U_J�ש�SG��z��'���`r1a�������* ��Q��̛p���b<$b�]��L%��}��D����ޙ�T���_��(�Al�x�bC^�q���A}�$oݾ�db�4��Y�I��M���5�+O�#Q�|Z�s^��5�[<��B�l���=A�x�-P�����6b|�Ù�[)7����M��'�1���9���d_3i�	���+a���~����6�`���͗�d�L�3�6t��~La��,�]1�N�;_&a,���^��������B-�� }�OI `׊)[F@�|�@��G��X��G� �U�_��/Z�$i���L��~��	����ă�D/��fY��F%y�dT*ׇH��X40��ed�{�@�� fP!�"}ncc�a�MxZ���L�`��&կ������v�����}����tcF륰7٨ā�4@�١_lp̦�i=��A����Z�vBV��J�#.uk��h��ݟ�7�J�m�f����m>�D�\�k�K���ä�����	g�uJ�K5�Ҽ���cN:s�ڢuع@��	4[B�*VG"J4�����RTd3@�X��K�GQD�pr^��`q���#����H���Ue�v"��n8;<�N������5����]I#��R\�䋔��mvK��o;$�:��H�����������я�|-	yw��}m�FzPW��ޏL(���ԙ���6Z��ZⵛoN`����uF����6�\������n6��Q(�H$cs���i?t`� ���y�)����
�}�@��fenZ ��.>d�If7�p��5SNO���㲮é{�8e�y���G7���3���p���ʞJ��L��5w���S߲�_�}��=�����r�HI�z8>�H�b���(]zб7��%�Q��>���1"&�����4���-q�a`	��\��Fi�V��M-j K:��Z��Ar"�.���������P~jt�%�V����'�gz����.?�i|/ <rr��#��h���:�!/X��hE<.�F�?�;K��Gչ�5�.�� uY�8S2�3_�2��SN�u�Μk1O�OׄSҧ
6EpҬKfW܌k�T*ږ0䲆-�>���2�v@� 
B�w��=tk'K��"�/7�4��gu���Bn0;�����6�WF�ѓ�ගp����,��A<� �oK��g�s�*N���*�&�	o����'Ih�;E|��ՅZ�����	�9'���'+���ʬM�a�/�tI��H��G�;�|#�\E7s��n�qƁ]��Y�~��<f��A�&h�;�H!�*�ډ�Y��<(zu-l��D2�y��93�������#�&Ac��64���:
�o��6t��b���/��"̸-m��>nu��`[�r
���a���t�S�P�w(4X�5l j�����U�D�u|ן++UkT>�.*D6-��/��^��C�0���T7�;��F\�0��5
�5}`�@E�ȞE^�~9Ty�@̆.��~N���ٜ%�P��t�߾�?S�B(�:&�����qgD��m$=o뵄��* ��Z`0� �����\��VqBcJ��h���[��\��:��sAd:��~\�1p�f�
C��j��&�w{�	�ao4�4�;yj��}��N*�s�g|$*�hW���;{P�!w�G�0�*�ҲP�̜�X���'s�N<�.��n����b��h5!/�|+N�	�$I�,۾������2�S���1��X{�Q5�v>�?SF59�e�?�B�	6�Th�z ��^��v��,s	'mSϵxi�A�U�6bF�:ܴ�ON�O�ڦ�A \�
����/��A���8 ��9�Z�[���]�����#��+&|�������FЬч���%<�Y��p� =�~Z`��+�^�d�9w���h��)<ԟ�䔂d_,�������(#���PG�d80��x;_3�/^��_���~Y��R����1�:��o����>\��ܣ��ayU�O�����N�C-`(#R��7I�QĲ��{��>�gv˲fQ0#LU��k6�.�9�
�1*�s@���\�~�f}�5��Y�?. ZLI����Ϭ���(�B*1��q�>a���E�\P���1�6�L�mf?����C*	��|�Y���i���"�P���E�,?1�;����!�����Z���qߢl�Ѥ���aUD:��x:��}K
W��*�oXWe	|���zg�ߠ�)�n�^_�{�)�N��3��d�ـu����kd3�ɼ��S������� '��D:��O�����$���Nٯ�H�(t��´��F�Щ���h�?�����\���n�V<_���4��	��@�Q���9M�7�KTC\��|���R�U�iߚS�>ԫa
�3���;����j�r��w���-��٫����=�(8=��*��VZ���i��el� `�2$H������\9�G�Q]x�DqK��j��i�B8R		��b!��;��Yy���d��Q���wg���bQ�,2O�P=������(�ޮx�._�A)���ݎ	a�S�-����5���l���1��n`�og����ǅ�m���{��N���տ�"�O�n���� <Z1��$c��M�c4���S���sZ�FҶn���^`63��(Q ��l��V��1b|��,�t���;�����n����Su[:��*���!���6���;@�h����/��+������KߙH������}��Tf
��O�^�N{�Gh
#�zh�ۏ����T�4�,?7���Xp�u�u�*ٗFP�ь�CH�ZJ�L9D��k�r�.�jF�r��q���Zbǋ�*��� �p��0t�و���㼏�BU�{�vM��q1���px����W|ReIKZ
T��9g9$�.j0�����\�nu�`�H��o�Ƚ��Q�)]������ՙ	�����N�B�a;.� UL.���_���۳��{'�΢| I����ϓ������y�}��c�����%����lCT�T
��<#A<c5�i қ��v��*��-O��{_�}B�{�Mf˓����Gu$~,�����7ζ�n���y3C��J��k�b���<!���c�}��Ai<�q�o�rD��'O}0���ԓ��g�9nZ@���F�7�?�ԅ]Q�tw��H} 9^��L���o�`��&
���!�c�8�H!SK�~P���7EB�r�2�ؼ".�;M��s�i'L���!�v�$��-�< Ỷ�EfxU���?�����v!ׅ��v��PF�!!!�Jz$�P��1�ަ�j�� �����\{4�g�b��4�� ?�um[w	�7����Y5dk)g��␾��7Kw"�PS�9U�]���<x#�!J�<���x��X����Oʐy��T'R�I��n㴊�������:� �Q��J���S�w��[�N̦E3\�7�t%٭{-�k�"�G��m��Xi^wo/�������������3X�v���c��κf�Lg8-�����AW�R��= -�������QT�v-ƒ��C.���!P�wVk��F�2$A0��8���l��/8��;{ʷ��(:�px��J|�G��s���ލ���mQ�h�S�+L���1fÉ�LFA�hb��: �Y1� �<��XC�6#�B��w�ɧ߲�@������8�tV���F��'�EI[L�k�Mp������6-��3�0�f ,&Ui�Kg'���]�{S��m{%Ø��ư���
��'f��paF(� �b���[z�B',�w{aQq�*��8��X/@$زCM%��p����!�H��*�����"QG�M�lq%L.���n�7��L�m=���>W,�\��Q�8��5U����E��æ�5�xc������c���MqK��[��j�N��X	����e�أ��(���Q�����N�c>�'��e�h�ͷ(Щ�ԡd]�y4�X7dps�q롆���,٫/��π���:���bg�B���aG{hP�W���	= }�nky�+�$��6m]�TZ����QDcԄ�q�Gu����k�_���O|@�O1m|�N������K�Ho4��N�)��5o}�`��f�T�z���W�'mvF���^�<x���.b�h���x�T�ק�
��Qf��b�W^���� ˽�׏�����,f��X�X��C�a�Z#Sf�=�Nqq��y�ր��rj�H�
>�@�C#�qT1��Bd���-Y,F<+p>&�:��Ȝ���Yfu<ft�P�xh��`O�,T%�  ���8�D����ݑ"�EH5�l�[3=���u��9��Z�b��z��Q���A� ��b �9#A��$��@X�g�Y�$�YK���=Nc���j;� /j2��y�a/`M��ۇg;�c��9�due7�p5]�n��0��O�B�sM��r�Џ#<��S����q��b�lG;�0����LO��������"h��~�4�2��12�Ԧe+���K���l�	/� �x}��|9��`Qto
]�H=m����H۰N=�Y���!L^-~�U[�WyQ��p����Fc��x�	�%O�@���9#(6&�(�?�������Gd���A���S�>�.�Iݎ!�#-0��<(O_�Л+>h;e���k���
��#�Zб-y	��u2�R#5Ƚ_g& ���wВ�M�U��j���}L�*԰n���t
�`jՋV0y!�߷�W1�l ����U�ʉ}/V�����������I��!���A�qsJ���߄bB$���Q9�a��S�-�Dޘi�)���Z����[/df@���D�k�$���͋�O����H��A7F�-��.�Q�;�o�-��9�9=��lߓ�|㐘�NѬ驤��a���I~�fU����*�s�S�B�3	���C�厑/gA&#��rz�c�ci�@z�n�iE�v:l#��"�r�=0��j�E�E��$�5�[<��H�_�!9��$��Z��8�$X��V���Q:�J��-_�b����Ճ�,n�r�4y� ��m�9쪊mg�~�\E��A�,R�=Qf�|��'��B�p�g
��\O&��`u��Z���S�ec�+�OX���3L&L�_A�� �0+����j�mg�)��z�0S!d���"�x�{$',��B� 7>�Z�ӈ�<��ٙZV%	~:����h�Ix݅�Q�1.l3��� (Di�`J��|�Đ'��ol�Ĳ:E+F�`�2�E��(d��?��H��t�0S5J)d��2'K���|�L��Ef
��/K�q�.���{Vn��7z�]X����L����g+	Hq����s/65N�nu�m�)�2�_8����6�X��ɬ�4��.�)�����P�?Byg���'��7g}vN�-�4cO�,��8�L�H�4hҸ��N�	OU�J�H��T��O/�]jE=�
ްL�Tճ<��`!-r$��o|^`y�������i+:�'�p*�B~$�q��P��w����WW*Y�ʢޖQ4��@-�Z��=5�A�՘N��>?�e�ʁ���G�B904��Ɖ`��|�k��C��&9�� Z�K�
�:¡�Euִ�^Fa� s�@��i�f�v('+rMYO�zq1�w8ͭ=�*p�6��7�c���Np[��Kjf�T?�[8�`��p�`�>�.Z�r�c.Ã�B�Ӗ�5Pz�4+d�A��چ�_$���a��G*�}�e�!�WC�QEѫK{Y�=�g�Aٷz�I�t�w$y�p݁:�@���+�%��y}R����3����%�N6���|%`(�1��Ӫ�s-��ӵˍm,��/$#���L�\q�ṁ1�^�IM�����/��F6�0.�ZŶ@�{9�K��� �\Z>s��@ `|{�"c���C`�i-(gO��+D!Fo�"�@��X1���h7F��3��ʎ�U��C�5��r�i�%�5�Y��Hհ��r׬�7kC����������
�m����� ��B����˦Y��:u��f��`c�W��1�>_x�̰�X�3C�Ft������'#�� ׯW.�H��v�H�S(�#��u�t�}�������ro�8������;���}����Tv/P�N��]v71�����Iз������.�ۍ��S��F���Z_��%����A���+����]U�09R�)�����]��;9�r���Vҭm�����m�n_��;�K����yԚ�	u�_C�YP�� [B��x�roSĖ���~7��e��Wnن$�
9˝L񛋺�b-r؀�/I�%���� ���B�L����a�F��q.��tp�&���ӟ�	�bN=���B� i�����a�!��N3x8������K!.n{���|��7��K[�+f�|����lZbCc��ȡo9�{�,�Lc���.�<)��6�?"�Ѧo�Skt����O��ON���:i��섏��HG�jE�Y���A[oҾh�11(��ń��Ī|�4T��q^�]t�s�'%-f�w�Y�w ?�*�����7�[����*�̭)�I�;@�
S�YB΋�.��+p	�M�j��lŕ�)#�����[N��E��pG*9U�O�L�h��ሻM���Cn�8����p�d��R�Ëڝ5p�ݫV��v| �Йk�z�a`v���C���^�����ĸQU3*Ԍ)���b�w>y�>"ٍv���l.�V��x��ӽ�a��0 �j6kU�ޕ�U:r� ��1q��������M�Ab�Be�D���rǩY%�
��y�W�D-�E����=h	?�_�b_������~%d]���V�2FR3�V�t����kW~��[Q ]�)��@d<�J�����y�k� *���5�4P�%V����q^����ʅ��Q�h��~��6�^\5[��@l �&5]*m�������Ѫ�O7�\�Zh�e:��KK�Di/����9��;���d�6��#<C�kb�$<+�?�Q��<���As=����Ʊ"��+l��� m��ڢ?�f��i�1z�]��a��*���S�L5]7-�PH|{��	�
]b�1x���d��,�ʏ���M;y���o�g4E�O�h+s��1�@a4n`z���H�:���+y�z��.�y��)�����Z���W�>��n�KCA!R�VQ��S>�+FJ���U����Qh_p�ӏs���ק�w���j�¡��ߢz���(���@Ǐ$�2��{��uBX �F���It4j�.��O (x<�ʧN��fiv�aD�&"�����Ƣ�9T�� �����s��w/�z$�YԊ=8Q>S���+ �nk��F�c�
N��:�kG��j������ۀ�Y��Toy���?��K�a� �����N�?��Q}�}�p�M�ۑ�/L훛t��광̏�RE�'�?��JnTCΏ`���D��y8�`�t����Э v�Y�Xl�a�{�}`�����U�����F���ߣ2���Lh�f f*���X�ND��<��8�:�O�-�ĺO�~m+ѱ p��N�!�m ��%�x�؞
�s�E|'�o�ԅϐ�;��:Q����7��JI��B ��_�?!�E�������!��a	VĽ �x, ���:L2�ܙR��2��S�Q�"ً��y����?�ہ�x�ʋ���_��͞����7���'Z��8��p��@oܞ�iچXR���Oь]��P*����
۶;R��C����0�L��W
yn�C�f�#Ik����`�y'|�G
Q	��vr����4�&гѺ�<��*@5|Rk�y��渣^�[��
�( �Ĺn�,���_�d{�o��YH� Vej�a���i��{��0v# �.?&P~`�Ϛ�T��J�{.d@aChx���Er�P{�` ���r(%�Si�W?V�
���V���w�D��������Dz{����.�2�~df�����l��|��M���P!���d�m
�N�%�Z�+)�	J�㬺��/�`��"ޞN�.���^�I�_JW_��e�Y@_sB�k��X��tm�e/�ܽf����z�쎭�)*\��w��ɂ7��>�"�S�!
e3���OK7�#g��,�� �y���~�;i�m�@��"0�_5A�]7<��;�P`�����S��>�edkoj+��ԋ�H2�9y咱e�,�F���I�y �V3ۂT@^<@UF�]��|�?L���)�R�bԭ1$���Ş�^"�$����H0�9�N��U,u6+�~��҈tHs��'1Ps�	����;����ӝi<�{LL��x��p5�ŝX�Lc��W�]B�5�����Q�G�i
v_���
t`C�9	�����ہNd˾?Oxٱ�����RO�p6��U������a<��&���œ�C��j��]��c+�����J��%$��M��Z��K�NT�P���=�D���Z�F��� �� d۪�������[��}��&3�[\�aK�}P��!�k`����0�ھ`}�2?�^�g־�y#r����r�Y��}~�|-,@,ξ��z��hFA�c��3]��u�^�ⷓ�HP'L���&����ܴ�������}��aV���+i��i�X���M$�ak�n�ב��_��Z,��$��U��;��,��M����d��/���5�WY�)h���=zd��x�� JÉ��G ��p�V������:^y��?pE��ʎ��%�d2����z�h�.||�RbCӈ��^�T����c"�0���9"_�?m��1h�pƎ�i�cu�h�*i�,Y�Z �_0�"Ы��1=9�5�0�l`�=��/d��[��ZΕ���>D��5�9��g*xA
%kq�u���y�)ԩ>0��\���v�������S�9�Z4_�8 �ʜ���b|`F���d�sN�#.J��"W	�����H�_{�����h��aO՗MX��e��ټ�a��'7��vkPI*b*ɿ�t<�ጙ�\���7��}#�P��ႃ�r�4��	�~�U?�8M�2c5�Y-@���og�3�w��':����}���4�'�앆����a���/L�Ė��I@�m4���;�&=��w��p�g�͡���	{����X�k�����6�ɔ�.s�X-��*CqG�v�1�Y�Ug�~�<�^�����&�[c`F%��~��-e�Sr�f�2��[Ȃ@S�0N�?<-�xh ��p���aXFw6?ל�7��HH>vx��35�f�=���@8.ҙ����q �0{y���$�W��f����2HJާ�dL sj@�f"�m$��m*��G�_��r:�ׄU�Q����ע9N��,���Ę��
oc�K�ALz6�LO�������
R���w��C�b���0s��B�!��t���x���K)����~��C�|��ɵw
0�N�[�v�Ƒ}�1qE@O�I�/P�5]�\��i��ÿ*�^����>���d��3]��w[�SM�I-b���)��b����}�f|�Q�p���t��G����47���;��W��]��H��Q�ƍ_E��š��Rz�
 ~Y���2��M!�v��6mk�f�f����/춨ó֗��U۴5G��e�-w�D]h��s�9N��Zs.Ry��.�1��O�\�~& �=�~�qǎ�-"è2�D ?�HS���,$?K�ҿ��� ˒�Gb���v�E�]-��J�I9�\����k�)mG.��Vs�0R����B/�ᛏ�	�*�2H�����ҹ�p��?�4u���p����z����|B��޾	���%��O��+4���:}����T�W\����;�b��+m�Rwy���M�ǟ5���>#��P��a���=�sׇ
q�.#K��Xn��nj��vk_�^��:�Gd�q
D���`��M$�)y�/��_��/��v�jNu�UIk���i��x��p�2�Ɏ�^7^O��p��h�-�iM*��"�5֪���h�@бbK�w����A��FHf�zsn�;�
����л��s�U$I�Q��'J��gҡ�X���7_��sJXQ�L扮E-S��	�Տu#/��#ozcp�%0!K9��#��*;���]j^K�L�,�"��hB5B�B��BU�e�Q�)T�^�s���{:(���p��	a�P�o9���1�4��IgQtE�o5����9���������J��c� }�]�oNu�9�M�(����jF��lX����+4z����K@��cC�~"�V���	s�0�@�����g��J�N�z�v�"[��G�"_�A�Y���D���cĮ�q�d��ʝ\��)��X!�w\��c�C*�Xh�B�<��������zi�'��\��ݤ[��{w8[G�y7" �[���\����E�@���wE�"P�C;�69�V��]0������ ~A-���v��<�} 3��d�k01���=x2��A�I�!��"'�5��F�����1:%��"�S�78NmYI֪�<��X���m�m6y�YdU-�Sª�n�Z�i|2Z4�cDߌ:-�EAS/q�8G	�P�L�����[)LĨ�R��?w���a}���FO5vVG�9�Fd�\����a2�r����V%T�Ǖ��6�v!���b�`*:�k�k�XV	��5Ҙfۋ3ȺxpFh�kSw<YCB�F�X�3�pNN68:����J��\�Z�V?\����P{�C�ӇS^�Z�l������Ɉ�[�������:�,g �tN���𙆯V�o�uYݕ1�E��zza��m�_���DJ"��o��"QR�Fe����H�ړ���<�����B=�
���� /D 9�&	 ���_Ȫ���HP
Prsn�n�e�$����;�@��d��-"�1&�i�I7��f��FL���e2����-▵ �2toJD�;s
7�U�E0zhTi{"dӑ��o`�(����� lp�>��`a�r��?TV���e9Bsj�u [(�5�d�p�$���[\u�����wB���Q*�N9���!$ֽ�e��Jv;x�ͅڍ<�ѻ<)b��}���r -Z�֓]!v�!.���3*?p��^� ]48S�l��2Єk(�
dI�X��v���w��Lo�Hw�����þ{���v�uk��L�W���=M-�6,���$Iݷ�������x��/���~�}(��e�S��r��'1&���O6�Yo�A�����o{Z~=��m�dF�QSX��_�/������f�]r7/��.
@��jJ���S���)�`]oI�xa�>���d�zr� �bi}�M�u5�n��nR��ϙ��@^��Q���)514)9��P#S��M�Q�������B�v��K*x�DrQ����a�h7G�w}6%�!����f��¤ۆ�;�M0����S;�V���]��Py��n�G^�*)�V�9w5?k�$�(�[�������?�6ش7�3�6ʾ�Z�wF�*��?�?T�'�$:��2����U�Q��C�w8�NP�āD�u�/��>��v�s![z�
�ĵ2������q�d��<`J�lg�!-7r�O�J߆[�k���q��y#:<��Z�QN:����|ܞ�5�!ݦƗ�Gߨ�i������ͧ&]uo��q�Q!t�Z�3b�B�S��%��]��̊@u}�}'M���8���MAzL/�;�2`�U���裳֘� �n)A�`e����u+'��*�8�d}�{�g(Fh�?�5'����$Rg�2k�-�����M_�!�9�F�\VM	Y�9(xx���B��cH�X)y�F�5���85.���UVjK��:�0�&��:�/U��F,��^,[��Y%�Q[�'��6�ݯ3#��>�T���n������Xx��|��ҷ9�� 9�]>:<�/�L��?��#%���0#��T-Ĭ�U�p���I^Ȟ6KĖQk;p�͠�`]��?x��Gc'��3b���c�p�m���y�K5���ѕ|��[¥�6\S��oJ*�" a���x</-���s�c�b^��/)M�2�����EX��}�e��=�Ԙې��v՘1�7���F���祖�o�wx<>9z̋�-��~Gm7����� ]/Bj��4(��0
t��n�8I�=��I�4�/\cQ��z�>�0�2�V��S3���U���sY�-�(�&���,��[?E�kS�c�V0ٞ���2�Ȼ�?��F8q˅	�
��'w5��`]q��qK�?%\ �@�[�����Ȯo�J��=���5��G������#�Y�k:�m����[P�v|�Y����_$:D�l<�u\��V��:|����'�n�>6��1iy8�"/�(7�'bF �iwM�NY��~�kf�X.�yb��oJ����f=�F�Jh������+�v�<#����n���h��"R蓛�,�$�4)�m~u�K�TŊ�E���x-w�S��՞�Ă�����Ϟn݆	�~�s����Vb�.�O7f�>Q��2�}�.�}�S�Fa���zz�k���\���r1MI����X���b���\,����h�k���@H�34O�L�Jtz����@�\a+��)�y���ݎ4�Ѥ������sW���r�;�M��iir�~�_�򾯶�qA�<OLy�2��u�w����<uv"ѻ�����/��K ā�>��a��2�3���O�G�܈���|`$�c�up)�oFk�]T������]�>���jkZ�Cf���O2r/����g����L鮐r�ڎ��؜��?���	e#�q�:�ctiX�����^�� p���mO��;\v���D�΍����D�6����{�Uk�e�s�p#Z) "��ǥg�#o*�Ղ��=���dʦs� �L*��վ*a7���;��o� �]keN��Gy|1v ��z�5έt�h�ܢJ4yxv@�����tVb��T)���v�.�f���Cy�l3�{X�􇱟�Q�Rւ�
�!�>n���$�:,�pɗ��#*��0�AH�40w���HA�'��#y���!
����� W����]|�sd3z���/\�v��So�%}��sh�ΛF���B���M�+a��u-"�1{�����O��x �w����Rb�
��G!���@���&f�h`�2�գ[�*��g�(�v�����ܦ+�4(��ĭ��d�Ր�_FE�����n+�>�~o,�R2��Z&�����8V��O�f��������3"����=m�`Vːd���h��m�_a	s.s��\\v�p Eqn���R<�/Cdi�o���vG13��Y���>/�*��^�th�^8}���\�$�I���l���vhʈJ�9�&��"R�{�s�V0Q>ICY�;�+�l�!��5xܣ*�H's07��yXRBi���(��S�0�@+ij���GQ8o]�ze�
�p��R�&�@�l��an����?���[݆hWrU;�����igM��&=���j|�4��%>Cn�l���-2+l&w�W�iMv��g�%�+�n���
˺H�%�G���*����Y��e����ķ��%� $^���h��ଧL����1 �_cU���pPkpc�v�*`2*G=w�X��
�?�4pp��È�� b��ez�����C�4};2����ܻ��m�RF���ڒ�����x�!Ub�3�"D� �:���抒ϴ�-)<����Vk����G@¢D���e2N���y����}�@�2Iє�{F���@ <Gˬ#@V����u��A��*<���UM���N�e���f���� |��Q`>?���7/XS�'����f�[M��4��Xk��Y7D!��:�ʡ�~I.��[V�<WE���Yg�B���2ȸ)>wjE����NHV� ڼD�vj�L�`���x�h�7Bʂ-��ao&3w(�4{�n�Ywww�n����_8�>3��[��t#LU^�3G;[��I������ �N'��V�������_[���~�?���{־+��±XT}s�ɶ��MдQtH� �
E��B�OU�>0E��z"Tdx��,D�%4F�x�
�_�:���e����ֈ,�h�-b�y`o�mK 6Q��T��[�+�O{1�v�]6��u�Z����}R�e�G����m�X���r��*ͻ��G��$���.�vc3�YA~��д�n�k)�/���F:���vӈv�&���{Hž3����'j1�J�i�h~h�Q"��z!�d�S^"u�yX��!�$f6��Q��C%N�]�VR{;Fl�� p�dK���iv�E���Ұᴱ8�N�~�P[�Ws��"=%ʢ�W���� .hYZ'�?]���f��s����b�vܭD�ъ�U{ew͔��ۖ�`��PuS�{?�ߝ��	�Djȅ�����[�+Tڲqe�Ek�~�Ga�A\�k���n	@Ր��͘+�)�Slpf�?[��6��c���i} <���pN��n�l��H�CKFps������[�� �����nL�a��]�k?����,l�ǿ�B��/$/��<�擹l�����<����$$�.���Ȧ<(�(͉�aص���L$@H���<�9	�&f4r�|��x? ����VA!�*��ٶL�ک�(Ĩ��O�V5w2��e�o���Z��&���wp���.�ʂ������;r��Lnvk��+��j�FL&]�O3uH��B.T1�V�j�i#[Ӳ����y՘֪��lZ���#-����
i%� Y���I[��\�����j����#y|^�C�!��Xl�h6��_�6 *a.;����da�$��x
M�?ɿ��ѨF��D���y��d�?���(�U��c�+_ą@�,��A�n�rI _�����٥~��!Hd����̓!1�ѐ��=��(WG�dҘ2�Ǹ@(ɦm'o��+\���8�|�G	��+�p��K�:vز
jȵOu{��=���!�����&����k1�V��uU�aj̠� ;UC6W
�k!�PW�[N~_V��Ok+r.�,i\[ĞZ���h��M:3�3�GcZ�ٖhB(a0Ҿ#P�0�E3�:Ռ��K����hX�0�g�JB����\̷�_t�a#}�eI�كKݒI,ԍ���X��������K͙
���!R� ��uaX��C�Lm�_ؾů�7C8PƷ>C�WL���y�6��3�Fާ�s6		$��u7�-!�2;[k��b����!!
�pm!�!J�#�]&=bj��6V-���G� n�R�e:�5~�㉣��E�C#�ՙ�9o������V0����6� 8���e�_ؼ�Y :��6@u�7{�n�����3J�)���3J�O��'������֫u��/U<�`RT*=�3�'l�������	�w�{_�ۗ��%z�-F��n4'���j��ś=�N7��`d���$�h�9�DurX�s�|�ل����)��/`AN��%"�[Z����������Ѷ櫅+s�{����ͼ�H�?8}lcy��6Z�-iU���Q�ET]Qi���9 .<;�(����{ZC��1�
�?��)K����t�� �=!���$R���/j���*[P�l�=����nE�rY��Td�k���˔�P1Al�:ͻoR����>��Ii8��X���R�1ÉY?MTpeF�֒4���>��n�5s��$(�|�[^I#/,<S�\�Z�^&σHN��So&b���86P��f%�l��X�G ��h��2�$��#�YRf�[!�h%�b��̄�׀�B�O�[���$y
���a�� n�"4�01z��}C��x�����]9#q��ig]�t�R��]۝��~���;�{П9���F����������a),�MY�Z;�6WWȜIRS-�aڡt��ӗ���}g��Y��3_
� YU�G`�U��/�:6#$�D��R���6ybI��]G�,��A�'yCk�m�3^��;g�K�Bh��,�O~�c/ͫ�k�G�
q$.�C���i�-�X`���e�/T(d�� A�����$�$2�`�gY�3RQ���;e�uD�i���u�Y�p ���[�Ӈ��Q"�r.�h$R��J]�C���0Ml�
��f���	w���yU>*��]��+�$�h��}<C���G�^��2�����B�j�O��UW{��ֳ�s���&Ŭ�ś�b
�m8,|�IK��|P������ݤ�y�E��)l��z�{����!iRF���eԳ�p�&������Dm��R|�#�]%����-	u.M���w�;wa3�浍��V��b
V����Gsa�G������'��<%�[�s������-��E6���*d�g��ºOΓI��N
Qx��Z[P��5�P�4���e��!���/Ւ��e��%N�f(Z��k�������Np��+��������NE�{�޼�NW�y��a��џ$��EI�'W7���؄Pv�S�j��D)��lgܧk�}�G�fY�I}��H��`���ɨ� �-��м0��x�Ԭ�przE� ��spy�9���0�yTKb;������V�t�vN�i�$�N�s���#PG4-$?ؖ=�c�#�;�@��+�hU��kr�a���oL	ع�*���a�v��S{J)J�IXwɋ�@�e��~]Oo}��W��vU�׭���%�>��6�JJ����:멻�AZ�h���{������x��(*<����5[-x�q[KASѰ�?�=�ܣ}(��$\��]=5wЁٶ�bI�}�����^j�k ԯ�r(�fn�u�@��z�0E2Q@�6�pJ��	�����~ow���֭�� ��fפc�b��s�5�O��$�n̥#���V8���`�x������ݾ�|�Ɗ����1g��%�>�~��b��A��`�g$p��=�g�8N7񧔄����)�3R1��)��4xF���w��B8��&���n9*k�٫ ݩpXn�����R~�d�.� ��x��5 9�
u�4"�I�s���u�b��.�OQ���cz
����`���_�U��UR��L�m�r�Ek��k�v��H1y���(,�~nK�sAǕ?�;-x�=��!����	���V��]��X}�hjR+���LL[C�4�N���9�_�;�⩰\�Ծ0��#�|	=&z}�S�ծ��kq�MU�^�D�6�q�ښ��#�L8;�	χ����O�[d�	��{ŻĈ�tYv�Գq_B�rU����s�W)�	�29rh��� 
�2J�[�ت��w���K����b8���-��&��&�,o��x��}\�t؟�����qzDk�	U"3qU��p�^a{�hUL�4b����1�.��!���d�kN��w@f������=�YS����KS`ét�RN��P�v��)���G�y*�H�Ьf#�]2&���k#w����Ux�?_��K�-OX���)����R�ꪔ@��ob[��'%��|�s��埾ʄ[�g0A)_�V�����S�K�MCdn;�aTY��[�v��ފ�޳v�I�9�f�Q1j^�:!jRaˆ
��1�u1}�v{8���n*�.Ԙ	�ig@�jHFԻ��0P�WI�3<�/�UC�$��%��G+�� ��8����5t������ܬ~-��=��5�|Ȇ�m��dC���:� v|>�qe ��sl�I~�<�H���5tM�h믴^ �.d���d)��B����Y��Pt���uP����4�Jl�����<�c�fldVo��?�U��A��`���<��ȕ������b;?�G����r���F���Q��_��n#2-�z<Yx�u�y���@'�v�o�暬��<�,�h,��U����w��&R�c�cc{�_`r���E�&�t�����,�F���?�}���(W�t�%je䤫w�pR�,b��%����1(	/��?��C�Kw;���J�#e�.dN`�x1��Na��m�6�O�u�zј<�-����F� ��s�(��q�O�`.k�;osW����z��^�������/1�����;�LR �WAG��9U���d�K�Y:�A���:qW�\z#�2��Rna��hW�7�|:(��E��A���|�����.�/���XP��tW��~h��W��!'g�o�,�i�A��|��"=�)��<gz����DG����d #��2ǥ�}�>��fO������c��_�ݵ>���n�=]�Zb�aEoU͸������~^�x-�=��'d������"߱p֎������)]��\�n��{���l��۟��k^�c`/�'O��z Q<��/L�E0W\�P��Y�\@�l�Ұ�҂�\�ߴ�d��WZ�~ ��5��%_��>l$�9���T�Z�z�j���O<�E�[����vV�o�L��O�)��3QH�^�)Q���Ýь3���T��|�~g�Y����h��Xw.I��$�چ�����ulZ �n��ni�fC13"|n�pyY}���Ppz��Z��2}n��Y��$�F�W�^H���V;�@1Cڿh�����ш򾷋=����ȗ2�'���y"��o�ϫ���u{2�g�hmI���^d¥U���u*f(EH�pR�-�Oׅ�]p�\JN"ݒ"&R|���	&����'x��]}N]�><X��T������~m��a_�$�l5	��o��a��qz�]��ɱ�c���:��[��:����s��*� ���	[��y����6�k� ��л���~9	����b8�2���5�A�ߘ���G /v"���V*��J��POmݩ�=���[Ew&���)N�ō�n_@6���-mq��|�F�܁p�u�2�2cj�.��K��V������{#2�߬��K����.6� ���B��.]'����e��Li���n-yj.�]���I�(��x z�'�'�SGQ�,��:�'�P[��h�(�����o���\9�7(?־�ge;��p�C;�o�赻�h�eq�?���,q2�u�Φ=�v,�^�
(���w�6�-9���e��"i����J�ݻJ���O�sz�:&�ԘĽ:tNZn�"�q!^b��ˢ?I�0�kb�C��6�@Wp��g'�Zs�z�w���pq�	>�<���!�ʷ�������Qz4� ^��:8W�M,�f�0!>���ʲqo��5Ϯ�*1��h&*BT�(��p�|0N���(-��M?Qg5�����5bR`�j��.�LY���y!��T��L��ٲ�̟���\�����,W�J�W%p���J��՗$�ӈ͵e�f���Z�[f���@�xN�V��5��( �(��uQ-�ks�9����n�O߹p�'�!�~�WL�� (�T��\z�6,�����@�O�g��==.q�1�U�X�pVO�7�}xT�9{Y5��G��ۍ5g2��7��
��ߘ����k��&�E�*	�|f���D&�Yo��2���?��'��l�s�6�<�)�F�Ӗ~Cf��x�j��~"�<Jw���s��io/B�&�U�M�Y,��q�H~���'�(n6f�-������h��"�2{AK��{N�@p6i0#" ���mc��'ll�F(s�ˋ��]ڥ���7zG�������k��~��+&���2�B�����`i�-�#o�c��~
L`�r�H��
��3Б����
�:�"�[�,Q�_`׍�����RY��9�
z���f=�(SL�1 J���g�[����w��y��@~|`P};�ZWPW(J��0q�Z6?ꆥr��)m�ܶ����o�F��p�{ΧK�51H#�f�آ(�Z9�J.�`60wJ]��gnܳ�ar�A�U� w���CMk�sC�_�
��Ϛ�x�<����C�_ظ�;�%;χӦ.NP��Dh��p��i�y5@<�S�=/d���hջfd@�s6�6Լ/�_�'�W���B�Yy��e���x^/6Uv��\Q.�͵{_�����k,&;�o�T����y�~�q�)��g6o�[c���(�ЏrS�c&��4Cw{� 3Ì���ڔ�-ɦmS�I�y������^��ڮ��ҷ2C�OO%������Lz~<��xZ�@����r&�R��S��	���V�� ��)���W��0R���@84�F��|�� ڳg���x������������!D��v}�b��� .����w�D5tߴ�[�,·O)�hS��5��}�e-)S���Yl>r�OG���A��PKX�`�����bp��`*?�U2�|G	t������߉�&��+�ٝ���������_��-d&Q4�p��}�K��_��*�+��Hǌdߨ�kL.O�yF*�F{S�v�C5+ͪ�f>7C�����+�E)�)�#wt��C�T7bV�1q���ҟѪ��.e�!6~�$����! �>
�I��^(��\^��:�J�YIm�����������&,������u��9����Я2y��+�ل�͐d2��;7N�լ4�;B�kԜ%T�J��{+p��a:�����v�s�r�s�?��H9��qd�a�M��}��:�)�ǜ�����}�]�:��u��)�@��f�*AFH���8��\ܒ����# �r�X�gq�Bqى�P�}��^��0E[�G�:Z�O�M�n����oh��L ��ۙ���/�(*�Z�+�C]m%��fY���,>�Y���I$�#�2��ע�-.�D6J��ݖ&s��p?OgI�9�
 /�5�L9��w����Xh,D�7��[�`���j"�D�����HWSlgv�(��p��5ԛ����E��et�Un�}Z�)��w"�k|��>��Ys"�U/���ݍ.?�Sj�(d��^�g�{u�U��`��s�P��A����v��&�B֛'h��s��
��m[ ��OS:�</��
F��h���Z�9�S�;n:�Q�`��CLJ��\�Y����GR-��1}'y@�a�	a��q��Ę� P�y����l��N�h"�|'՞��6��OjP:\�m��Օ�e�6��UC��ci�Z��c�*���������綠�
Ļs��ձl>�cH;7^֚#��1O�=G	5+�F�[�$��<�N�}.ׂ i�����;1.;A�^�%��-�N��9��_ @CW�H�׶�@�Uɯ���ȡ��|:f�&`��&����"����3�nk/C��1��u�qb�i3{�p��Wҧ椁���	�ӌ8m����
�������0�iu$`����tN:���@��!�r��b}~���:�R��Q��K�J�o]��Ɍ�v�/\/���2ѹ���:ip��y���BV�oT�~��������J�*��Y�-'���"�5�,a�o��,��� �����RYOe��_�C ��&�mQ{~�@lN���	R��`�R�Ȑ����&�O?�!�x�R26�C0�DV���B�9�� �#��̀|1�XaM�kA�������9l]��2$+���sێ�C�80��q�(���&���i�)�e�/G\s�����Oe�+�@?3�_��;�)٧S�ݻ3Di`v��'yc�3PHş$e���v�f(�&�+����҄�ǉ��Ć]�'Rp������6ĭ����d�;�&?yR�v@}(u�cP�Nl]+S�?�W����y$$���`� =�،��ӓ����i$"�ur�<?�I�JL�BZ)A�r}^�Έ���[$/�S�V���Z��0����`� ���1����v�5:M�SYu�É9�%�Fz�� -�A��ˡ�¾g�6l�cx�	*��.%u�+jǳ���7�>���@�[�!R��L� ��0�PE��4�(�4c"������d3ʡ)r��o�nL�z����
d�.E�{�6X���-���ָ�޽i#ʍg��|�Q(�0�lbWnOp��A�5m��p��m�g�p��2�w�s�Ö(5X8��NR����\#A���/,��1}d�81���68�]>��C��+��.Th��z?��������ύGj��Ƹ&����n rDk>���f%f��a��k<Q�����!��Gs&��M9�I���OvO϶A���A��	a�ڂ�*��PƟ8#c�3 N#6ه� ����e��|�э�YA<����w�C��e�8���{�ͼw�e8��ŕ�|Te��H�F�$ꤘ�*��C#}B���c�e�K���ͨ��/;��u�{����AsZ
��C(u�������u5�FH��F:S�z�e@��<������7g��0j 0&zp(=�|�8\2��q��ʒ��M�#;C���d�ƞq,3X�f8�����<[���._�M��o�N���K�9��%���p�98�����?��#��j�s�><����k����{��1ݟߙ�a|�� �*X%H�P���͙�F=�����J-�y�'��c�A�����tT(AU����@J�z`�,O�L^�J5���{0D�xA�S�K����ע,tk�=p�n�m�Յ���j�L �-a�➅�	c����ʩ֪@�K2�NyB�7/Ue6�FNl��������֥6\�h�����&>u�?.��+�oi�,��z���V������Y����	��"'��9��*w�~e%�!׺���º*�čj@m���+��<�nNO�tSb�`pB�D2yL|�o���ֽW|W�յ��O��d�kh�x��Y�(���ۂ�k[����2]EtmW��,g����u�X�3惟QBͷ��=N�s�Ճ�Ozp���J�x��t>|�j���᱘T��p9��Y�'~q�� A����J�6�"ʞ���2�J��k�[z�g�T��s�˛:w�iVc�s����y�!��p'�r� �)l� �t�gV|��|�xﴏ����B����}0�_H���Q��#��b3�C�=��5�L�ڊu�	��h���B�B�j[9T�#cT��U�5_>�V$Ӊ ��J��ݷ3̘o8��R�2S�ع�^�����'Ck��b��b�@�A�?���7LMe�t��4G.Gh9��R{���� ��ʛz�w�Y�t�dG���h4���VG�M�ܪK�I��	�]D4�uϵ�
����z;�,��@P�aJ�^b!^�>��΢�<�5��?F�Q����Q�\�<�ٖ�eN-���A��76���;�Ϡ��6���zs9.�(��m�7D!�rt7�=���]g�|ߔ��q�q�����Э]�n��8�s����s{����'�.9�	���(�#�m�o/u�1u�f�сA'k������vi�'O�����`f�1��W�7h���ք�X�^��-tI���!�חX���*���и��ƞ���0�85W@� l,��QK{��̃Ռ����b��(27�AְZ������ɐ��c��AY��y|�-�D��!wb���rq����M��_F?�d*����空E9���yd5�I'?[�����7z�:�N��b��qh��+%c���RJ��H�r>DE)ޒ}�� H!����%��X�d,��+�^��,&�j(�4�	i��&殺��$��zV�)�Q ��8$U��9��@��r����?�4�����3��҃^�͹ �J�Y����p�&0��������|���0(Q�
rS�;lrsa�3[�@_�8���,;�����s߀:{�|w��^���:�iNY}��fV��߹s�bp)���%_LG� 9�I���c���U�-�j����� -�I�ĹJ�bk�R�6 �õQ�:b�-Ga�&��=���f-4|�0,�Q��:�p�4G���*IES��<E�#�z�8��4ѩJ�<�5h�%��M�ԔO���^%��� H�3��/&\z�:d߇4}O�
��#�崭+m��~��9��^�̼[.�n�Ė�48s�� ���>P��nH��bo=�)[����:�N�M|���n��?��ad��#o'<e($�C~�Q˿n��ū��
�mc�D���P�m�P�#����,����Aچz�`qZ�R]X���DMs�σ�.A�9�O.?b��O`f0@SL�,�1��|�5bg��u���#����+��G<]p�xp�6�d%���9f��	fp���^a��B"�Gx8��EG<<�{�e������9��B�����>83W+_����U�+ëo�MGm(i��X��1��!�ib��{,^��?�FD��y"Q�;{8���Fֵ֓�R�G�O����;�+�|Q��$��zi?D���|��6��y�1�<�[j�< ����Ny޹����������4Ɋ�����ZS"z��p��K-&��"����;�r⛺}�2B�{`GI��y̓�*s4ƞ�bXQ� 6�
�j�g�%�9�6�LD�h�a���[(pj$$nT��+蘠�$1�O�v��k�>���A�`�s�=��c��%�ƔL�θ�_6S�C2�fD�6�gN�Z̓���>��/�>�� n�J�c]�ן5Pջ.��)S�E��u����:�*кC���S��&n}W�'�����lCZ
�H��=���d#�����^�I��HL�	j)GU�@Yj�K� �9����;�!~%�+dF�QW�UŅ/قm��-�7n�S�[�0<ZZ෱�U�b��hG#�Xu���@�{���VU�L���8:[`�iP<�ϗ�=�]A EL^�>?:h���/]� ܠ�f���E���"��t���E�^�j[1k<ϻB����w!ldD?8J�����c���Bs�5�>��8�z���?�i��z�%=|���͉�B���r�Ù����m�j�~�U�@�4���E���c�Q���k�S(EWU�--~�l�R���W�T�/��mx��^��BKɊ�g��42}����(h�?��vI*
�U�)8���*n�����wM��e�^��R�k��Q��4���p���?%�	qJ������G��D`d�J�p��y6[|�8�� Sk�h��ag��.�l~D$7 W��Y�7|Z5����)�PUͣվO� �bvt)��j����F���_��"Vk�6^�w�+Q�L��{VI��`MwxQ>K����%o�Us��!����k����ycڶ��f�>���ը�!?he�g��#[}�,\%Dq���X���N`8��Ԧ:���)·<�2'r�H�-�a�C7"^$�Ѱ��O�r^F<�Ko,>Q������D��D�y���f]�\q.O�؇�>~չۉ�v6��e�B!��5�4�ϊ����<��5��	W9�B|N��5m_s"�+��%��p�
7KK��3+}�4?A�0�0�q3֝������F3����9�=SH�L
S^����re�jxS%<�Fa�\7����.dk5~g�Y�8���N6i������Tڃ����l&ҝL턌�] �ܫ41z�Y��D�jh��%L�*M��KN����Qa��Lx��s\�s���6F��_%�;6��.��m�������q^ij��c�[W{�C�&��(��mvyz�����(}Ge�)�t��KRe̲:��2�!�֗�1U]Ym>�}��=K<l�k,�D��P-�]�2�n������9$@S�yQ�t�vU���g�疒���1]�ںF���Z��:�����ӝ�;�>d��&#�/�JI,�����pB7�,��N��]m� 核�V�h��o����=7ʬ�.<弡�2�<�G�H+���<a3A�����TjV�[5���%f���~ �q��U���m	z/�7
'���L 1�����'h%���H���< U���0�g��_#���}����9ۆ�ާ�i�k�-�s�l;�kbQv<��5Tw�I��c��4�L�`q� �Ba��C9G��� R�@���銗׍�hyhf��10�-u	TM\V�ƕm�<(��뿎YF,H�$a:�$�gĪ9���tf�.G�I�~0�Z�^S�$����t�t^�����w#!�N�ֻ�N0�IRX�kN��3�	;mlV, k���P���p��"�pPɅ�o�²��]��w�����%dE�>lba�O{xjQIzo
������.ŉ��*T:�ms��e��������-��m��R���9y|$"R�����ӈy�r��\���T��
�g��w��s%���`��nNO��ʕ�Y�ׇ#��NЀ�ٞ�pča'��uϐ���Jh���c��Ԇ���(��M�5gu��%24�`��@������sҺٱ�҂��\�ą��a�P�V�4�O9���v��L-���dL����g5Qy��˄%^j��F�'�(	�̣�(���;��������u�j�"{���ñu;-ix(k[׶i{hE�A��TD}tZ`o������g����Aӛ�ۣo����cD�W�Sb8�0�>\��EN��s�:�Tm��њ�հ�	q�<9�e*N	=��	��[�v|�@FZk�J?����i5P9�K�qo��������}k5�Жx��UY��l�_>+<���J	h�WѤ�'���*z�/p�
���y9���9�4u��&	�Ŧ^��l6˒X�嵎�T���6����.	��b��g��e���=EcX�`�V�[��<�7�NKɐ���cs�ڊl�/(=sܬx�`��Yb�B���зj)��Pz��>u��% �ej
9�0Q�E�]�h��Έ�xE������̋�>��a����,�u��ȃ�O��Q*iQ�R5�K)��;��x^p!��"�+v��@
�ͱ��nOA\	W��$+��T{C��-r1d������w�64{���.t�Ƴ�<��` �Ye��NQ3"��?i���J�����mKd��1d��	n�L�iR���Nxw��@p��x�w��>�P��n��1g��z�A��6��7�wMTC�@�ԩ@��Ggxt7��Dt�����������{S$�/4���3��*��t�A�l���R�A���B1hކ�L�؎��㲺h�#4'�J&�_�%����gn�����QX�	{��FRK���-gI�!��$�Ũ�Eja1�������$Ҧ�Ҷ���]��Mo"��kCDE�bo�{�~0�G��ȁ�n`>�R�[���)�}��ᣀ(��~�������\��.��G�`�P�� TOSU��1�M�<�x�y?Ok{'�����
��A_X�&&�R�z��5�vJ �bX����z��OI��N��tK�K���oV�	y�v{#=1 �J��ه�蒸�J��@캦�2���X�G�z /%2�j;�����NH��%���$�nG��ŉZ��'��ytW�q�I��`w�ز��s�{�W����Ѹ�N�2� 'KY]�y&6Ŀ�qm�@�u8J����r��+���K벤zi�/N����z\S�__�]ۆ��(� ��;�3�ʞ�=�B%����W����`��`S�-S�&�=#��gf?nj��~�i�'��Q�"�I�U�p�E,����~��j�a��Z�.���b�r�,�QJ��O$ȗ�E�j� w`�Yn%s���  ���� h���8b����:V#��\�C��@4�.�񳜘��u�ek[�6����#�v��[����'��)��]���M�C8y�C�1�5����YIA�n���D�����x
m�{W���K��$���^��aw�/�\�����ɫX4���M�n�����Ф-���˙�^�o�ܡ����nb�MQ�� ��K,�<���6S���!.{%��1������3��U�%8�n������ã(6�0�ʪ��1iO�xf��52��+�mR`z�*�� �	�_S=��H=m5��k(؇�cس��NL]g*�+W�t�����Ej��[I�h⽞ߌ�V��&�j�ʲP���@Wc�Wͷ�d�
(�P�F7��E�>a�v!	�N3dZ�)�;o>Q�@���js�rC��5���-&�r�h�aZ�qWב����y��è����P������!GQą؍��ȓ����WW��Y���>23\�D؝�����	�x������zI��9@д���&Xv��J*�܏\W*��Ə7_X���WL���yd]%����ksʩT	�MM�h��Y~�Wb0s�,�!�o&�\<��=�ܛ ���=��)�E/Bǩ�X��{�8�d��ň=�vܣn��~�G�,�����g�.D��I��?��I6�zg?��[�����?���=8;�c�K���Y:3�7şw6�w߬��/�h�rf"���xz�-֐t[��w}Lg?��L�M���m[F�d����&�j�N����r�< 'J���PF��=�#���A�Z�C��'�G�r�nf<7�aw>j�P��Br9���^���ʏ��!�����S)���w֙�h�I�o�:���p`4��U��ɇؿ�f�f6`F+���]Z��b��n�@�DVi�
�l��b#��f��S�>+�I������k��U��a�Pn�$ ;nt�@ K<���A2r��(���z\Z�E�߸�Y�D���
|}��<�V�kӧα�%0f�MZ��:���-]�;X���.E!�4��kJ��U�\�p��f� �
?,��X���8����jѾ6�<�����`}���bFVㄦ�ՌU���Y�*!ؾW=,����x��f���'�1������:*��({��4���7n����U-%�ɫp{�3�߷3���W�~&υ{&{*��S�K,4+2Ċ/�ܥz���:�e��F��<�>Ԏ;�T�SR�9���Iu��W��$	S�-j.�b0I׾Ļ��~z��I��It�ض�D�g�2&�7e-λ	5YA�k��xO�dQQˇm���8m��&���W�3�̈́C8�q����z?=>"|��[j��h74t�ks�|�yv)���� �>}�Ǡ��s��W�X���!t�ry�o��!긽>����$�|7r�:j��v6��2~F�k�~�'? ��s��U��iO���#�OF~E�̫`)��*M�Ȑ:([��\wa�?[�D����R�&��w���$��^8����vC�p��XH��/���p+c��f�����]8��c��-�il�d�7�D�b�H���l���k~5���W��`r!���~�e������}�ԝ� ժ�wgc�L]�_6�M �xj�i(e;�~MY�vД�*�gfe���&���q�?�R�_�on4��1X���V:�J�(	�e�
����NS$�#�%N,g15��O�D���}ڕ�]E���9��T�������<���&�~�m�U��GF0/�g�7K4y$"�M�4��(�]�䉕�Kܮ�ޢ�}���А+X�U#�v��A��~�V��c��vK�ac;�>���W���F=c{Yڙd���;�e��R�L��ikZ�	��?�bEcC�W��c��
ޒu:	#j%
q?�����-�����F��;�<����
��%ȍ]�r�(�>��-H�-�O�K�}�!M�O��'mj�s ��R�u�stM�*va�N�1���D�R�Z�0�U��������J��d��ۙ�I�3�+����!W�bm�*�]n��{���v)�HڋmNN�{��;v~	�G�
�]qy9:��p�U�A=���m��I�C��a�t�H���Q�[��\gb�28�<�9�_�w?����	�|�/�a�r��Ү��°����I4�ѫ_���[.&R�խb�e����Q������PM�y�;��!\������b+H��2�d+䷚ĵ!���eD�xב�68�w&�Z]`%a�z�Ӟ�N�j3}�7�I�ú�]q{>�_]����UW�����me�7�"��,jY�h?#�0W=Ta�,ۦFȇ�;��C�$�o%CW�9���S�f�7�y�z{	@��)�Xι�,*�xW��u�A-��И|������t��Q�,� �u�����5��o�t� ԍW��u�!h�̳vë�����P5���H$U�(�i�y)3�1��Y��a�����:Eథ�-�����5
�L�7*��"s32&2�lY�/��Eݜ�q���pXIh��ح��*�PCȳ�t�'��.S�VrG�y�w���#�e���4dp�@C����C��H�r����O��M��L��A$#e�|�w�[t�u	����go���%�l�&6(D�m��n0���K`�ˋpbD�ߪ4J��c��Uď�0iPD��خ��=9O�Ox01��x�n�W���sPZ���g�뾮�t�-MVD�DMW�N�4^=��8��L�r	w���^vꁖ�!��9뢠@<�k��_��h���(�]7�+�`�u�9}�v	�[3ɞ���g���q�Ji:��H8&�n�ңi�mB�C6�x2���h$J�0�r�q�{Cz�����q�&j���J�D�r�_X��2�?	
��%���7q�a<��q[��KZKɈ�z���o�)��]�jU��"	L��@i��7�0d�1�U6}!�X`	L��?�In0k�y�	*u�KG��;��pN�Q�#�z�<�x`�Ц�0Lu����Z�%0��zH&��f�����<dk/ܬc�;�/��(�9���F��RN�~أԟ��ŭ����v@�t?p釣�cCI6�K+��������e��0��x�$�C ��G��	ܴ�`]��4u�Z"Z=&��Q�撫l��Cp�48��LUP5�)A�'D�S"�
Qv�zE���!nC�� ��%E��َ�f� K��[fa����
���国ď���Ya����L<j�����r��n�Ay������;�0$����0@9�bQ��1�+o����^҆C��Z��,�\t��;�ϻ���P9��9?�8w�����m���瑳JW�� �7�� u��>*:���!z���ՙ����Ӡ�%�C��ܲ��i��kԱ�nΥr�=���O��� ��v!��T�hGU�p���-���s��"+����^tPG�q�V�:d���p4Yʋޅ��|���1�^��J}��󥣮��s�	p0I�g6��kq���q���wW=Uhti�s��Wl�g)� s}�:����՛�^��l �8?������V�3פ9:��mYWF�1�󞚟iG��u���	�z��p䀛&65��6O)�.*��Ñ[gL��0o`^]�FB;��
��s�x��`���-I=5�~��Z���^в"m�cȐ��T�X��b�ޡZ�)��>�w�%���e���W��զ��ۉ��� �7�8H�' ���{�R�[�A�!�x��L��W��ɱ�r��-]��͋!�J��L�+��d���B�Ǳg��L]�����k����"��	6.�����d1������:��5`�/eh0��ğU��z@I��:"[�"��6�]i���N"�"괒����F#��+DP�@������s��5�my�gd�ZǓk�R��K�lhy��L���i��g�&S�"X!E5�����L.�_���4�3\Ep�1�@�� ��R=�j*����C��2R��(��x�Ͱ?�_�/�4��MȌ���6�y�Oڪvk�Yb�_	+o %��i>��dt�I�+��4�*��uv���0�|;t�1�F��
x��^��HP8eK���H�R##�"CGo�<(�%*���=	�v�J7kq;@]-��/��c�����|���>�~�k�M5%p&*�_�7���2�2kL����5ۍ��_�<�J�*P�@J0����1G�x��[za�fFS����hJ뢟RW��\�=���r�T֤�=��-?u��O]�� l�,��>��<6��ZR$c_;��c�o950��u�s� m�j�*#e��J���:q�v����V�n�O{�'|A�R�'>�lL���@S� B��v?�)�s�Q��w�c�VmhTX����
��r�/X	W�k�����&m���A�yH)�����p
?�E�N6�6�D#�.����P�.�@���k6Bb>����14��%5ǇR���)_fL��T�:v')��H��h�	�1���}��B΁�p;�Y���efҶ��D���=��P�MI���Z+��pH�C�&��[�d��bí�u�D��*?74X��IT��r3����W8D�'k�%�G�o��kC/.1묠��V쀢�����[�E
��8�]rCup̖˄9�Ҍ���ir�)�(��:����z2C��9c�SR��+�������b�2� �u����jN�(�#��S�����]�^�;��˖��<48�sm<���]S���!4@���T�E� v���r����V`�;(��m�"�E�2)�9G?�gWRG*��0�촟�����B}�u�:��P �h��3��G��{sh�`�^�\���/�eA� �r�u�X�> �iY?6_�N��z�h�͖�V}6M�D$��e�!�ݝ֒!���G����X��Q��4�n�yΤ~E!�@�iի��O���ׇ��u�%��SYђ[�Bv&��<�1�-0%*Usd 8we��7���ْ���;0�+�8��cS�O��m�������� D*vi���es��m9XN��q���W
XL8
;����׍3t�!�EVLb<�'�Q�L�I�x�$�]�q��@��u�K\�P��$����'���(�l�Ʌ�������v�{?A��o���Ǩ��:���껑����$���X �$�a=M��8����ݴl�:߼\J^T�t�����V�8�0�C�z���d/��%�f�5p	֧���R���f���a\e�J̭�W�N���S��m��4�e�VW�a٪<�Tc�z�y��H��_5.�5J԰���$l�����:&�RDŃ�,��Wf��>G�{�˅�fQ�n`;Gʗ��QSP�1���H���ctFC.��7k/���*��}�<|<˗c8#�֠3�P#�Cŕ0:p�"˭���B�D�{�m�ۏהq:��M;m�iH���nL�yL!�QlN|���K�Nk�Vüg�C��r����*�b�x�(!g�o�	ep5 �@�HC��GTM�T������W��zK�!�>�^)^9���j�10�8 ;��-��1���?�X�%������1�|zk�G���!>�T%߱x�o���<0� l�-j��T����s�ȹߡ�f�;��N�
�0�����~��Pt"	-�M����G��{2�:���x���eo�����f���=�"P���=���^��E�'NR�)�ڕ���|��C�c�U�#�v<�߾��nK/D�W4�*�)ᛙϱ�|X<+ggU�A��C�9�=lD1�i+X��%!c��}xC"��ц@h<��)�P%n��#���$
���X�E%��b��q!�r�T�Kse<l5b�j��:%a8�gS�]	bp���y�V����Z(ō�6|[?7����yL��bs��y#�E�\�S��t��ڬB� 	���{Ut�g�T/�����) ���꘿ʶGA�"��H��ns=�4��[e{��w�	4�sd����~_�eB]	؉��<H:����|�9x'��(�DHfh��wͧ����l`N��I� Z���o�l]h�T�|H)��ڸט2������/�FP����A���>[�_�[��/tӗ��L�Z��\�2'п�����J�#��E��=��"����%*�|�<Nْ�]5��v�XhP*5�z�[�3g^�,�ϱ;��4�~.��Tr���~ z�޶#�#�ܬy��X� ���~	���ǈ�r�V���,[��k�kf#HzC�so|B��
��PYj��6� G�{^�0��x�X���O����w��G��T�<�_���#dzyO���Y_}}��=��>��F ǲ�mO��o���8ɲkg+I�3�[\��Vvk���t/NA�=/f9����jdG��G��_|޶�XW݂
�Eu�-��
�?i��t�&�������	� �r�~ދ(�oR�iO_$M�q�r�?*]�<m����ԝ���9�n�
�7��2��5�z�0bl����M�\E9=��
D����[����T�O'H���:Q��L���8պg]�@<%�:�:g�;�
.���]>�.�A���K
�w� R�C.�`g�3	�4����p\�fV�Y��P�<r7ѿ���D�F~��\&�^�^<�UWȕ�wi����3��uXj��s�(���l�'�DM�D����n7��G�cS~��?��KT���q����INBA�My�1��#��7(W�{��ף�5
+9���ӭ �*���	 n������l�"6�,۳މl�<i]���?��ͫz�C���jL/�F7r-ٸ���ٸU��F}������G�������il���]$Cu���R�ʹ|��GT�b#��t�@�������/V�*$s���?�O�����1Dڸ
t������+a��6I��=���C��䮮�$����3N�����j�q��;u��6�i[bV'�Ӳ/t��ZG=�p:����H��*�i�rE�baL�Fy���{�!��	J����� �8;�����t#M�cz-v�����{��Q�%j����/v��������z#]��|AT��(ʁ���2}pޞ�5Vl��.T�:��Wk�6�&U�O��7����$�r'��\?�E/��c�WΘ[������҈7'�
�*���{E�� ��ڢ�h���m*+՝���`z�%I�� ��U�u�Cz�kQ�ᣤ������Iz�:����Bܜ2�&^w���:���W䄨k�����u�n�y��gg���@���!&�t_���)<��7�[�j$�Z� �j�{��I|V�&�H�it�℁�E���>�B���ƞc�@�κ�P�K�\�Cܘy�YN����2�����C�� ����'o�4N��K�v�=�s�J�x35����챛	��"+A07�X������M#ON�uG
�xN�����ʛ=��,4���N;�.�Z{�Z.����@K3�:�.a���i��<]q�#*Y��$p}籜��o}o�Y��K�v >$�y��=�i�穴���麀z�]P����I�MI�Y���:N/����?�oc�&_��� �{��z��RB�>+�"q+}��,���D:ߝ�$���da�\���q7yŋD��;߬��뢆)6½�#d��>�"Q��M�u��6Y�ύ�4�'����:�(Z�</*b
��6�pp��1`Λ%�´l��h��z0p�)�W�A��R�ꥪ�����8W��B{b�-�q?rF���
B�����g�W��z����(�2og���{P���
�c�ms	�L]�x(��i�3�\�����s�ÿp���C�M8��̭��=n�yv��4<�����h���/�Ƀ�G�f5��^�ARNV^�"]&�ˣvf,���6I��ׯ��[�`�(`��P^Τ�{FZ_��+4�@���7R�#t��ߌ���*i����e��v*�?+�tx��WV��Y=α�&cfË�]�l:O��^\z��C��g��r�6K�[��a�J�q3X���ejƏ�CW畞����!w[�2-�6��*��;!���:;�C#N[����Y�>icU�VF��Z��27+���hف���R@-k���ݵ"oƜ��FH��T/�v\�a��wqp�aw��l�,&<K��\��m�.7��,��2 �T�w����%Xz� L~�D��fO/S_o���!�@��C���p�!��	|z�O�<������g��2�d�Ȇx��	�_Nj�C�	i��9��W������:��_0�O��j�6�[��tZP\�o���:�0o���m��y��W�nuʖѐxV���� L� S�~�������'�ge�a-(s�5,�)������ae�Tr�e�h�Ŭ����1F�o�ewk����`Ar��F�r�BB�[}9:�~Yӭ��1�1�q&.�4:�,�CdQ&����������m�]��=��[�a4J��&��˭�
�vZ��3��vq�7�Gr	c&��w��Í��lDs�������;�T#�e-���-�T�|��ߐUu�L�MTW�5/�J`��9��)��1�FBFQ�~[���&���-�p���G��glt��+�t�puUo�Ѣ��$x��>���ԭ��_�s�!�wd�>Eݮ����A�+�p�\sG�{����?�0��d�)e	���d�=,e���p�X6��������x��"��Zuq���I���]lc�%�ʜoZ3nq(5?]h��ǣP�|'�gպ���Y�����Hn������@�r�������kA.�ht���+���1ס�Ho�#���+�Q�6왔(7]����o��{^2�������K԰:�w��fK�H����%�J���,�k�︰w�k��Pj�(����mG�����G�`?��>�{�s�_�뵐�BTDw2��w��W��2Y�so��Oֳۘ�
~�'�T���E���j�b�(ҀW����q�t�	��A߱^T��'��_�_�����ߢ�|{^����h�d����f��)^bz��Y���2E���r�P	����~�ˈay��q'P�[׺qf�
��Y3�*�^�&�ū�a��EBa�Hm���o��mē����1Ⱥ��P�3��� _�V`_���G ��Pۓ�hF+��i����N੖�D@
c^E���{qt��u�̹R�n�����¼���z����H��w@[	���R�T�7���A���B���a�]i�S_�9o�I����\sX��F�1��AL7��!�G��X��3(~�r��pja6b�Mv���rXr}��<D�	���/�YHWi�mb<}>5wW�d�`�h�Ä��g9{�1J���9u�J�KE���<N���>AB/��i�c�ݞ��N$����^��+���'f�fJ�ŗ��;�_͆+�җ�:rR. c.j�M~��-�J<��a��`�8���#���{2��� �x�)\���O�	��V��2��2�i9��УJu'.V'���J)+���Jh����LP����7uo°5S�=6l;t^t�+	��i�*N�<oA�����T�tN�G�Ĳ��*>s8�0���\�{~)А�j���Lt���Z������������,*Q<G9�j�Rq�x���� ���K�h䓽���OI��S���G`bm��#��W�G�sD?����4yR��;.;Ae�x��V�gU��$Adɣh��K��A�9��kW8�� ���_ޙ*o�<u�y��Pn�-��Ab��~����1�|)�.%g)�*Z���8e������Ӳһ�"	�#2|~��DK���С��&�*������g9�x$�����7�)��������$�C��A�e$�Q>��1�,O݅T3��ZX=��RT{�z� DX|$��Us�ltE�g^��[��0rk�x��k���_b��,/Cp�X�DËvl�M#D���웸,M�Hi��K�ܣl,�(��["��E��`�M!�P8ɸaȭ�\�C4���f
$�Ge���3�\�!\����a>x��p/\�"_���8�_©��{t��h�~���L�G%�c�gi:�l�A��������x���� �h؊}2Q���8j��B}Q����A�5��A���ݬǚ��zގ]-��9��nc����&�3>���=�%+`����Nd�s Ҷ�WwH�
��:��B)+Mt�[,�	<C��1���,�R!�W���&�=��z*�:�<�F�^�W�]�vk�_��@b	�&��q�.�@���P�v�K�w"�5Q���/x�rb�fj0Щ����Nn�* /bQj	C�E�
;��c�\de�>S�uO�Q[��x4����%)�da.8y����!�֔���T��/֫\Uq�0�:�6��"�ᵔ���7ڂ�$�j�3FJ�)gzϴ#���� J}Q���Ʃ(���J�GQ��#�#���}U��4�K�z�z���!@_k���#J�5��=���{Y��=��S�������>��G�F��k[��5.�e��kWO�o勋�����(��Dm6�=ی�?K�"�y��H����������g[��zO�嘆8��_͔�<���|���pti2Rܣ{(R!^&`x���~�96�B4���Ê���=��1�z��B�
�lr0��Gg����^K�؏�h1�:7�+E�󗷴{����:4��?[$F	���Ŝ���w0C���u�<Z��UeV�f^*3��Ա�|�;�v� �yk����QPz���fM��9�,����b��p|��<VIQ���ۛ61ͱ��j�`�-�bncl�*$k5�� fT��i7���s_���n�dDؘC�6哺_A���2�=A˪�˪n�y�q��6" ���������1��t�٘�eB{N�~
Yo���P��G��!�����wE*�摟�`��>W闀�I��d�^��۵v˫����Q��1��8~֧��/��#�_)~��l�'�ۋiesFk�'��U�z��� N������;j�m����ֲ�ҰdL~.�Ȋ�i����Hz�d~*N��v�CQ�d0(_����|�>R�OFp'�fH����g��儫D�&+���������f*���K��5,n�>Q���|���u4�"6������6���sl"2*���
p�1�?��(�qE�n�+��4pČ�*��=n��b	^OTT�tJ"�2[�!oVc���	�@�Oͷ<�_�c�OQ�pJ�C� ����Bb0��Wm�!C}^"l�0N����ڜ���z�5��L�����K�`3g��������D6u��9M����b�ӟ�m���5�uy�P��_�E���%q��������*��v�/��%�5k��H���1y�8AoTU,�Sٶ�A�\t�z�I��j�1Y�,S�&��-����z��Ao� [�B�0�d��ٲ[q�G�"ΆG�E�<��(=�]FPٱBJ�uSc#�� ��w�#!����$���óts��1���KO��j).�t[ߜ�D��K\��uc�����PA"�\�/��}����X&` r����L~�u�E���.lCo���6�\�=/�g�m��EKk�����)���U ��o�Ő:��2�,jG�� ,g�� ��6����v��`��"�Y����x�[B2#��{Cz�!�h�Ĳ3���9ֿ|/D 	#�!ʳ�a�=}U����k��F�Z��[BZ�d�uR�	���Um�	E��4<_�jt)%�Q�E���'_=�˓s���΃�Q��1s�D6�t����-R�Z���B�g�+�烪1��r����5_mr�3�8���uk�u�;=���w�T2X ����;�pv��Թ��^��O�v�"ˊ"&������l�!�Sn����a��"�\/�<!(9��{���ۻ>��S����jR[�|�@S�rWjs3mMuV���(�U
�LCF,nͳ.�e�A����2����\f�VY� �����w7�o�4��.�j87�Lf��������VFb梄�xRc_A�R�Z����Y>]�HG�$+sg�֕��i��t��ǔ.8�f�u[���٧)R�rD���$D���KD+�X�8��f���W�NF@��V�1�[8/��0��O�c({\�u,=�Bb!��:��S�K4)�fgٮa�JD��" FF�A����4��I/^�/�:�O;�b��7>��Z�����J��aF��/��9C��s"ZBa�g.�Й���Y��#�Es�$lwp-F!�J�enU*���##��Shn�el}�M�a�B������j�Nj$~UC`��E	>2��\�Sakϣ��젖g��p4��^;��^ý�sn�.;f�F}d/� �Ӝ4����]E`'D�I�(S��q���	�eR�p1`��ZȮv�<kM��c�2�����	�R_ ��jM�bS���/`X�fG�*N����a|�֌L�'��[]�r�E-�LP"/�)��5
�}YsC�_F3�F�7V ����{��a���U�T��. +Z��AۂA���oWs��ԖR윛U�'��$l]�}�vo���Z7/�N
"eW�dJ jn�y����6�ò��_��l�7E{(;a����J����YZo`ۓ�:Ofxn5�+{�/3�+7Q������̇����B
���ϽD��·/{�)ӷ��6��aZ��X��ݏVm|�����ڧ��E2�g&?�p�VR�KcYod�
�C��¨8 ��hZx6j�a��Ḱ=����a�a����5�;����x���j\��x�=E�<��;�`w,?O1�(�wQfHb�%�$U�#о�5�?2�e0�wj!uʂ{��w�#8%��5��nM��dnl�T�t9���w�F68��K$z��fW}`��4�9+�Nh-a4���cNC��)��iۅal�w�0��.�G����B��jS���rU��8xQ�t)��p$��g�XH�)%�Ku�n#�p�ЮUU9,X�/�v�v�[����`���e�Px�1�2B�^�.�IZw3�"�뎢(aܱͮ	H�j�b���M��!4�?g��׸l�l��璦>�ߢX%��8�rg)	7�x���S*3	|���������f�
�,z�\����2�����q/��&�LVz���`-g�Ð�s�
,D���c��<��i�p𙈰n4���B��^�|�#h�=�E�� H9[
�(��[b�ƙ��y���ؚ�`V�/¬3,6�o�=!���_Q��Z��xm��]�G8묆�?���P�|��ߚ�"ތHjA3ib9�>F�
��e�=T�H�7?�A�	ZXf��$�ID?Dm��%�9aF�����E�������U�
�)W���><L��	��� *��>�� l�q��#>�f^��Q��1�W؞LQ	/J����h��3�Q�m�6X�'�G�O���*�!E)��p؉!����[�I�Ԫ��1I���|F�ZQ�r�@>�e�����S��~ꟍn������a)H��HTG]�v�%���kB�eu�tL�����xi"���Y��A�����3�]�n�󕫹�\V�esg�~*��j�,��
��M6)�uC��0�S�~8_2eo,��m!�/ƶ��q
�f}l31�}T&�h�6�h���f'�$��5���UP�� u��?�3����Z�Ls��Ok��}[�{�1��ث��w�dM Um���4��G���#s;P��=������"���5�d"�]�<Rb��X�jIk��7T'�<@Hg�/�Ɔ�qrv�����3-xÚBȢ[�h�	�pyI#�Ԅ�n.}��t�sYlʱ_�z&������G+����k�����b9&���W��ӗ�����;_@�������:V(�N�c��p���ι���\�n���U�ut斓1�<�>k�_-6،_�Yx���:Mj�'��܌w�
�5�W�im��R.i7
V�)W�k@b��:7X�>���G�ۍh��|%��)#љ8Nl�e���y#`��Y/���d՘r@w/���u�
U�b[(��Wx�qF�?vȟ�h��������\�p��O�*��5�N�uJۙw�P���6�/sf/���E�]�p��P9)l�0��ǵ;�z�}�;a�f<U�փG�!hM&��3��}X
�G�#�%֯m^�w��:e��`��P4�i��`�)��y�J��m�+���%���a�ՓʖyV.��C"�?��G̈-�J�F�?s��~'yl������DP�s� p�`���a�\�.b�,y�?�`WM�P�YD���s_[�t��NȻ�|�by��+�>ض	t��a�q��fcg���4s����U��po�pH�7�T�SSy��Ӷ���LT+j��m�E�Q�ܸ�MWG�\I.ZF=D�4�����<ѠX�Or�J�Y�����~�=�ySf�d�f�uE>B��~�������&C	�@�a~M��Uؑ����p�E������$����:(ͪ.{W_�i~S6���G�z+xG�
�=6���wҚp���۶���d�8�U���gy!��.�əw:pֹ�пa�U'To��#���u�
�����yD�YCXw��Y8׉�OOڬ��I�|y���*\BXl��~������O+R�0v5��hGrEG�o� e��w��N(s�ON�4�p�y^������G,����I܌���#6i���e8�Y!�����M�.;{��-�sq�Zϛ�l$�,x���!���8�մCVD�������߲`�X��~5c����%�dlllC��X���X0a�H9_�d�b٭fbhmq�?b_��A{�VA���r�Q��DjCO*3���Zǻ=���&{��k׶�t���m�^����-�1�9�����I��6�0;�7z��	Z� ��n.���I�<R[�ں�����V'*q*��/�"-�p�b	��T9Y��2�>�A��Rni�s�-IyS/���(.3ɖ JQ�<��l�fJP�b�*�W����T	t��NP�FRs��5��n�/��tۀw��ێ��Ul���\OD,�g/o�|�@m���ڴ���G�2RO�HJx.<�W����|�z��`�8ڿ(W�gF�Q��p��C���(�I�gޕOd-E.l�N�映i��U$�ߴ�|l"�:!&[*��cp���d���a��)g�\SJ�ŀ��>��S[5�* ���� V9?S��)�����%�@�D�h����� �
Z�.*�DJ�����+��G{��6�^B��B��퍿�c1�$H�=��sH��-��c��p|�Ua��B�yv���m�y|̵�����j�ۛ��.�׮��������.hk^]҉�J�����=3�/:3��� ��	�~�I.���y��}��f���hq>4F^a��c�z1'2\r��XA����L���Wy�`e	E�lR��tS6�tDƩsYی�7h��X2�/��Y��^��gʝ�[�ƫ�i�x�m_�N��@tЃfb�f�v`%��j�Q�h����4��7��]��:�����vdG�QK���Hn����_��(&T1�:3ejV21�2�D����Zi�M�Ym~��in�n�)�G��R�o��� I�d.����}��B��:��/��P�\Xbv��L�)�����3i@v�'�b`���:�F�G[@'`���U�s�O���5��J�͞f�RYo����������أ���4��v�緩��ş�o���e��.�ʇ�hZ������t|�f���Г�h�m��s�s��K��:��P�2	 ��z�V�Q5���HV��=���.���@�.���s�$�һȽ�G����8�:fz~�c(lu��J�wK���ۜ{ ���0��{�W��y���J$�#4��¸�G����/*�t���5Wz��d�8b͹'j��F{��r�vA<w��xh�2G�Z��G�{��"�)J�$W��t���2�i�@�%���������iDI��0�d֗�.]�fJ�,p�b�_��\;V�u;��`Y��q:��� ��[� ��l���G�q038� 
�~tz����i�m���1�cڐ�^l�{XA�j9�f.�����2.��,[���}�21����b�r�ګ��{��v|�i�W���t{
}d�ɨn�$�5ub��ɶȇ���+bb&�V4�u|��j�t�DJX7�6٤���7�����@5�cY�	��斯�l�<������!�I�(�^�S�τ���m�B�'xZ)wF.s#'�8�x�n����&m~^��|[4����÷8Α�fҶ=��}T�������l"�e�,:�eQ�VNFsR2biD��h��+�v_��������74Hd[$轣Ғ�5�'e�\Xz��SB�B��M�J	x6��F}�m*2�
B�_ZHY�`W�������WЙ�z��Ռ�UN#~��UO�����Ke��m��3����,_<f��C`Q�S,r�l����c#S%s�P@S�G�+����+F��� �%��^�d�1�X�c>55F���X�;b]�f�k7��8A{���j�X�p�V�{jX&��?wנ0x�6I��?�yw{��x4�����Y�BP�$�_`��x�m5>XX��FЙ=䭀�@ëK��p,�%!Cw�]�횉�%ew6�,l��m�JȤ��,�x�K^��_����%����lS��`�� s�����IiO�J�7*L3�:H�uָ�[A��R].�Cs���J�bB{�4�a�#!>�6�Acâ��ْ�cϥn.I�moR�?��cr��!z�7���.��b�����d�W'�f7q�!ڋ���H��~o���jqi2�Քi_w��(i�\��cLY��5�N���NXU����%K��x������		k"�WY�(��d0��Ff�rȯ��2�$(˺.�"(���(�S��bE�H��gd K�?�;�p���g�p���W���1��z���'��^_u��+��3yډ�O7*�@�z"58.i�w���\��P�=ό��1��8���u��ˆ� �I�b4N�jL�ehӸ�*
~���-Ze'7·z/�DȵP�Y���"���%�"�3X�]E s���,�n��>~Ύ��T�WA���)8Iw%d݀�ϱ}x+{>����0|s9��!����{� ���X��:x����VF��;��L�!�B�uj4i�y�e����:m�>�kTM�Mv/��/�q4���=����H���6�QK�x5c�_X���#*��"��(��?OW\?Z�#����d�8뺖���zjZy��D� U+��1�4	�q
��F��Y]/��j�)�����"��0��
�y����hDC!pR�V�_f(�'��l�.��%������N��蝭�.���j�Ǣ��<;m"���D�?�-��3�GS�����.l-֦�'�L/����|�żC�r2[��Rf�N�� ��Yq�dOl.΄{���d���I�����&�.��hl��RJjmI���_�e5 ��:0���'Q�H�F��~N�o��*�I4�Z�U��O��a/;��5L��!H�F�֝8;*�/Z���Kh��l�ݸVg��d����u�M����Z&A_�/)2�0@�#���b�(ҏ�_Ǆ�#���0,�ši}�+!�q	�iK�g���l�'w�M�ͪ��d�o�;�d�U#�}��n�̑'Sp4�]K�������;TFh���%]�I/�,�2eWJ�תp�h�:5V�6����glE	i�LJ#{g��P��po7z�I%�[A�ux�3�/ ��-��~,5��1-&m��>#�n�s�!�ň�{�p��Kg׷܉����(<�ʪ,rܡ�V=��G|��A���x/���l�Yz��l�J_��gN����ccrp���G����R��a�u��[W������ۼ�a>{k�)���������@��$�X.�V�J�����5~�7&��n���A��3�<�vi�vY��3`K0�}�#�~>.-q�"\fJ����?��l�Ɨ��\��=gUjy�ُ�y��m9���j���9\�Bs0�I�n�#pY�BkH���ԉ�-}c^�e�V���M�"E1�����⁹j���+���b�W��� ph���*il�8��W���	�
�Ŭw��X��!Y������Z���3�"�e��¿��`EEs��1/   �i.:���hB�YpG):��K���.�u%��c��n��#{�~����1�R�r�����E��N�/is/�bD�� М���v���$��L>	���`+[�Kr�E�A�ut�r�Ĉ]րy��<�S�h���7e��K���=r~"��#���d�h<M�3��"���Rh@�3�����l������z.g@��S��[N�x�c�$,rU~Z�q�s`H�$#��w�ɵ��{�x��|�1�$�@f�T2��l��[�k�Y s���3�Y���w ��ߛ���2�nFQ?�z�)��冷2���}�
�C����K�Y
Sπ�I��f�a��\���������	-\PC�Љ׶���<8��rV�T�o�y�4�"5�Z!�j"�GEj,�ˬ�.��b,�FS_K�@��c ^�%)��,B��z����6d�/��c��Z��<�S��hQyʅ/A�*2�V%�0��k�|���a���nǖ(<宎��KL���MF%e3:ha�̱z���h��k)�~�`X��$���f�r�3��y(d�х�{x�	��ft�ؤ/�ѦF:RG;G>z֓G4C�S�q���y�����q�����R!R��`�:�O�e��6I;!��+^��轔5���)�C|E;�@gP���a)��>i�]b�T��I��HX{�#5+�z�wՅ����5����K��b�kÚ�]��y�$z89q�J�����\���k�����ag�ڼ�)�w�~:1��W���ik��}j���eD��N9��	#��/�ԥ�s\smC"̭����A��f
S��-��T̆UuuQ��3����ǆcڨ��R�P����[�L���R��۴ҝ�4C��?sƻ�b$)�}$�h��<��Z*Jw��!�b"��6�r%U*�k��K��a��Ƣ���sNݽ�ZUՖ�����Ӥ��a��~��������m�^u��Oؓ�=a�s��~����u�,�s���:ۛĘvE_����{e��#jڎ7~󌪩�d���V��=^U��D�c�EV�'�P��@ڧZ�H<��b��z�o�c����o[ΧPnja�܄$>(nx/tv��CvT�7�mȏ����|A�R�nj�� �4�����u��=sS�S,�K�*6����5;�NJ�����p9'�g��ɚ?���\���^^@u���Hn	DIZ�6����� �TE���;Ԭ$p{:��n���r����G/��R��?w���&*t~�se�26�Q�Ŝ����L�f}���ߕA��El��HcW��@
Zʲ�\M�Ey�bї.��*D�t�9j�21������1�O�=�r����ϹG�"+�x�cW]�D����g�[��½�E��� ���p�A�$)1�֩"�nfޗ��Dϴ(f�#�Jky�<F�߈]T⌊я��t���c!b m���ӽ"B��:&���:͸�+�h5e�E2��j�6�iE��
٣�����(q��O��0�P�xO���rٮ��ATi����b�n�S�<��>���Ί�7#�F���#:�O!��`���@��g�o��R(q���l����0��_�/�Wf؂��^�d�P~�K��D~����5�;��NT W�5��R�k���8�3�Z���v�CT�ۈx#(���ཽ����۔C- �[|�4a�}޻�zb"�p�5�<h���U&�ۗ2n�l���a�o��q�U�r��3��WrQ���0(D2'A=��Z+r�vii�Q�U�W��ǖ�\����x��"����|����R����ژ�5KՂ�x�L���b�i��/α���P/Ÿ׉Lv�zt��ů��(5
���K��� ��5�إ�B�
u���2���'Й��=	M�6��(�{ی�p�	 r}"��R��d�t���e�<pl�%����Ń�O'-F�-��-�3� �so�������!j���Q׫8U~��ӊ�>����:ͱ��~��ie=/M�s�^��5��ځkT�"c �� ;Y�$Gj/�u�_h�G@\t �	��AOcb�8���M��"���]�b�[cN������3?�N��
�}>�U���)��Y?��y� �K PFW�!h�g����k�7ݧ�s���)��zsq�\��e6�;ϓ���7U�o�IaH�k�W����=�C��Cc���	$h,�M��HQN���z�hFr��±/j;K��XR�������UdwhO����RL�^��];�W�"��:Ŏ�]�#IQՖ��N�9']�����E�'p����;-����'���8�V���-`]�l�S*�S�w��կd�J� 7 &�7m������>�I ���<�;.<x�@ڜe�Nj�{^��%Tf�vI����t�Ł̎���ġ��H��&s�U�V^�!��M��Ag��@�mhқ�-ŉtS�����ʫ˔N7�%�� �ӂP�h_�~(�w��i�B"̳&���I{{ʫw�u�nz��XO̵��3Հc�OSe2i�~�-ڎ}��Lc���M��>���Ø�ّ]d� H�z��fat���z��O	�C$'e%���é}wPFg�;z�L�q7>��{���UZ8p��F���b �1�PUUF(�.%��a0P�ݎ�aDP��_��0���	9h�w���<B�ݛ��0��m��7o�6���Cr4y �i�Mg�#H�ۗ!�,��40��4�����b�ɜ�N�U!L]<����~X;șY~���LS�6u�V����dID�V>Y�좮L�B���*��2�K|MG��%5�bD@_P��%2��T����e ����@,۩��E��4VF��B�9t'��3�?�[{|�xU���>M�\�`#�����)2��AgQd��e��Y���k��j�o����廙��r�:�8���������D��hrF=T)1b�"�����$h}��X���{�~"�����#��C؏��p��:0�@'�m�`�V�P� o�Y��2������,�����s4��G��C��:6u�j>�W�/����j����I���6�pMi+��Ղ�6OՋu�����4��,���(Ӑ`!�B���ZT�=gO/t��OtG�<���0R#V�V 0�d:}D]3z���V�$��U��G�H���. u)|���f��źr�Y��xǡ�y�S�@�p���'�q���KJnS�}�`3ͳb���rwB7@�Z?�Y���x���c�fwn���?K�6��V6� �XqdL�C���:2f�]>���Er�='��/"]�fW?#��@�d��$V� ��ѽH���4Ep>�����I���?�r�3����yH'���H2i�<��f'���q:�Z�+���L�s�<��h12���
��'�������;��~�erm�9���jF9�`�����װoB�YTY�IHeoY�a�f��\��B�y�@]��Y����W����'Τ�zy˕��MY�Xi{��֛��Ŏ�;�C�_{�_�#Va��y�ۜ�����N&��GJ�� }0h��̝�E���i�����L΅�9�*J���ѧKg�zỪ$k,����@���>ʫ��8� .�y��r��Q�V���]���RjĆ�������8"��M�����'�D�)�0��	��\��S��#�&�)!��!M֕F#��X���e�qrX?�'�p�h�=�e\�G�M���K�w��ݿK�p�Q����5� r�d�q�*�`�	��T�<�yz�����67���y���$*�����X�UwES��d����J?��<�5�h��(�+���x"��L���>/��p�̾v����mZ��3�Vr�WRX�c�Kr�3e�E/� *��j'�m]4�OqA'(IP@H׊1*:wt�>}�tH#�V��u���2���Ae���@7% �5����i��}�&>h� g�B2�o������Z�&gk1�HZ۷8��w���!�'�1��/�H��,i�%�,�*���]1vҜ{�p���§��v:I&��������������o��Ro��Aof0XIBٿ9���Y�`�N�k�+z��`�=W�eT�I��v�ҖȼE�*�$�mO]�6��~�h3&X�M<�oKl�� 
��+�'�T��Ƣ&�ى#�^�Nt�t���J�H��7zsg�s��Дֶ���ǟ�Ϝ����>�Q�t�fw��큳n��Y"���e��ywN��X�����4�?��ͤ�U�� b�$w�IY�<*ٹU��3H�~�>��A�W-���B����M���+f�`���˜k��+�&mK�
�}�A,�W��1���%���_U1�un�3�L�r�2|�}��3��3������c\S<��3��@k"*�04�^�;�ļ��#4qr�@��#���9�cT.�6/yPU���;a����9۔*Y*Q��U���h}��p�!�F@�K�[R�8XwZ߁�(�2Q<���a��.���M���@&$�x=��6��@wKX��S#^n�ܜ�� 5�'�E$G�3۷�A�2K�#���W�+���Q7Wx���������|W���M�6՛x��$l�����S�I�M�WY�φ�{ʆk��b��呹�yA���\��+m'������`�B
a��DJ����#�𨴶���!σ�_��?<����e�֮�D?B��̋ڴ2�j�S6���"S-w��XM."X�_>֊P�+Y�«b�'�.ߔbڻU�����_�
]5�B��n����ds;����%��P��:~�u�'>��EeQNq�a.��_�6l/!N��\�m.���C%u�g[�k����H<�]㯲�D���r"�+vo`|�Y]6�\�KkQu^��QVٍ<t�0\��%}��Ơ����(r�U���-���5�QN��wDՏ�J}YR��v1q),�
�9���qm-�+n�4��3l����z�K(�������6ܓ�P'ڞ��ac/�RB��V�4�e�/tb+x�O���<�<\���c*BuOI�:��5�&g+��+�>B����wV��hj3f�|�	���~�U���ז�B����я�#HO�����E�
�~��&�L ��Y��`y�;P���+�16y��K3艪Ђ2<�wP*�}�ioC �*~���
�����	@���$��E�R���/�_9���ӕ�L]���� �e��'a�#����D������15���?�1Q`E���Z6�=u�˼6:�$�^$h��w�:1W��N,LX�C���D6���^#�Lam�� ��GjF5W���vi}땫䨫{'U;�㠮Р�ǔ��){�\Ć�@GbL�'�r���z������Uo��4K��UiƊ��`|��(�t�k�Y>���z�;6S�wd����~q
�B��F�D�5����h:.{/��~�ۖԬT�o#�Q�1^a޻S�VG�Ӹ?D��G���v
��Y��g��X1O�����)`����!�t�7��?%��CsqI-��`����1�H<T�Y�}p0V���s�Sj���FNe��P��$E��HW2g?6�V��������������+����
_K*
Ͷ�D�Wdu��ʲ�4�G�Sʹ�=k/��z��me������VP�����O�9廙��<� �����𝯴qs�Q�E!��x2xٛ��Yy�&_j&��>��W�j��A�M�/���t{�V�ǒ���Y󼊲����AϵG�M��\Js�c�b�ƅo�P �|4����<񮥦_�x���z�C��=q	ĄT�I>Q�����-��~r�%v��C�ONjUyb#h�O�4�)�Hh�NR3�% 0\�8�<�Hע�>Ҕ"kNS��)a���Ī��)�C��J�:��5_����(��v{�F64%B��xQ�_��Z���������ƙ�Ϗ�&	�s���%{0I٠g�S����k	�.c���ƍO��p)ȇ/������C(��+؍�	��G�s&q���D1>W6j���+�Р4����+�dh���8��|��/q6KЦ�;���[����(���4+JX��==��s͎�!,B4�%A��+GF��L�G��0��o #̺?�ގ��x]`��z�q��Da�^�Ձ�ذ���3�x$o덝ݨ"��X�z]���>%�����֡��xf_(F�+{�:%ى	��m���嘝�ڿ�t�3�g ��є��^3��z��]G����BR���01���^C!�\9�9����:�JONR����1��t��f�R��R�p��jF�[�H��s�Z/E�*����ok<@Z �
��
�%����#��1%���AZ�Ȭ�M8]ĒP�Q|�Hۀ�~��!�r	��=��Z�P���HJF�^`e�O��k�������q�D��W)���mv��$?Vg��2R�0�%<���/o�i���.��cwW�*����Pʗ�zu-�#e,9+�הdB�xCy	�j��$��"��%
����}���ȅ�����iQ~�?�"ېTf���g�P�18���>$VoI]�gE�ų%�C �:`w�+H��4}|�	݉�,�؄m)3]0�&��R�k��.���#K${e0��L{Z��`�.�;�;�O5���4�,�'D�12*ʯ��ހ$�/}�{4	�^x�ϤXx�J 	�e�?��^�W?�yϴ/�j6� �9��<���m���ʒ�	H�/id��n���B��z���؅9��m'��`���0h�$� �"��LW�J��:�� ���r@��@�F˖R򩞍qT6:���ݸ<2�d�u��9�o�Y�l[�%�nM�F��PK���2�k�fK���M3�>�� X>�a���L�m5���:!�[���uy2�%g����..�FE����0zS�qHaɴ(�0�?f?����Ӻ���,�767�ŗ���ك
*�T��c�K6��i��㵫�?�Qp��{�7h�j3��Mc��+]�8��=~�>�*�����0�u�LDI�s�Ca\HE�f�<@{�]�5�<<Bk��Aۿ�5���h��{Z@���S�5�q�J��롉S�`����!�`J2�iI���u5쬡�#�B���8L��V�w�^
�DM��>u,f�qI�5օSY}E������8�V^^Y�qA|Ѽp�#�������
_jƼ�J�/gV{��5�Vi�,� �o�v7�6���������VqZ&�`����]�T��J��v7U�y?��KI��iX�в���2N���DYG�O1^�����Nq������?_�Ix�_e�p���l��#@��UF�xM����^���W�v��gy(s}��o$;�@ /$��<�%�C�Q�?�6�p���"yE�����ք�Q���u� ��P��r<FQ92eFJ�:�������kl���ۣ��Rp������WLx�Yu�6s؎�TВ��@c�h�utbY[�T­�~�՗j���ĉ[���r�-E���}�T�b0[���^�dp�k,�U�dL�XC�]�z���
D����"D�ͽ�.WФ�%B��j�
�oŴ�O�"�7A+�nP�ɐ

�&���0�S��|���@���L*�(g6�E��o�J��*�:^k0�;Did�]�W��ZK��q��(�<�Y�	]��h!������c�9�9��>�+�ӯC9�$�l���5=�����a}��n�=\%���$œ2�z	Y�W`K�@���y�}�2�Xd�ߙv��"q��c��o�aF*�*+�V^~��$�ze,�4��o� �R�b*������|"��hs$Cg,d������2�"��bKMO��J0i�h�u_@�(�3ê6��]`����W�`Fx�+�ΒEj��G�94E�Kj��r�\؜����o�L`��x1Kv�J�r���b���a���%�tY���)KJt**��.�MӇt5����?���y�陶����7Ͳ�%��6Ĭo��TT8��ԭ�+��!��JA [a��M$97J�K� �~�q�T��������5?�D�l�p�g Ҙ��׆�0����vj3cu
����6�PN#綍��BM��fs����|�qK6�[/o ���?����E�B��wp�K�|�� ;��#��s�����1��'M����#��W{!�^�w��1��X�z�ҠZ]+9�e0D�=��2,GD��N��P����9��3��"�P��š�X�-��P-�.��R��)��=��A�K�K�;|��=B�6gP�oV6�	��u���l������QXI��>=�\ȃX��Ԫ���eʛF9>����qЩ�D/�R��A�y��e��VI%~���8.0���Ш(lT�Uq�B�,�Q��ѹ�x�U[;!����(��wZ�`kzv��6\������M�<����mT�^�5>`7����e��C�9j������tLW�U+��f2�1���z���������|�#��r{��۠�Bɟ���g�ZP�.�V��s�E�f����{���B�\R+|`�~���%m�E�@�*.V4�`��R��|�J���Mۨ�v��EYݧ2H����$&ȗqo����'g�����$g�&	�"�օ@�#�^�$9�z��F� ���$�J�q�%s����P���]_�Z0�2�-p�r �|{��C��]_��(�g�!�l,����J�\(�Zȭk4��aPP�$SG�YS�k�d[������p�"ܮ%�a3|�8��EV��RbS���uz����F�-x%����%�?q��Z��,}���X��c�Ej���g�JG��\��m��j�fx��p�pp�-=�m��9N�s�,��-����m]@����r�	ħ�%����騷��4y��OW\ۚ��3 �`�2(6SM��i��L�>C�
��O����k}59��	�z��]��ţG5X�S55�����dp�e2od9f_"x��ZE?�[^L�C�ү�*o�>Ɯ��-v����\Ɲ�p��nB%�q��쁝ք�����%p�\�3`ĠH�^>��[��* �z��p���{k4�q��j<�N��Ҳ�2	ݕI\t�|R���f��>#½Q���Й7nER�-wӶ_4����\Ac.�H&y�l�z>B�c���ȉ a�������
��q�
��#���,����$�7_�>�F4������l�]3Rńh�J{� =�$2R����o��Su���-��3;�=�;�{��ږ��|���Vw���X"��B�)�~L݀҅�XRe}<�����ag�$��v�:ds֧ �G��4`�޿&te�|�n��X+�)c�CH']�t��Ӄ���r���|�$��|��2���g��8�RUʔ�΋��Й ����p�k�6]]���C�\ �oSq[k�Q�f|UbC�Ӣw���2>�=�_�7�mt'�"X* �q%�ڑ�!\���#]
��UYoz?��c'���c;lGzO�u��*D��7�A�C�P��@�$�j��W$�[���]���1�S�0�t�}�*�/L����]�8���ݵ��W�>E��@~�"�E~-͝ѓ�69H�\��\_H$�n~)�%_�ܽA�vC�0G�Ǝ0�ޟ�����+-ķ^k�F�L��6�"V��2:~��ؽ�l�3z����]���D��tb�-
�]r���V��Ϳ�N�K�������������RTX�F�2 ��|4P��R?�^ɯē;%�� ��2�nh}��ϻq�ۈٸO���csLƣ6.ɧ�N�^�3��Id��� �לJ����h�]j/�)�Oɻ�u��Y�	�|�i��c;�*���ola�-P���cC!���gZP'��F�%�:q�oj��2�o)$�R-�?E����`R�����P#ͬ�D?�pZF�������%'�s+��ʧ ���Z46���`��E�ʑ�%�R��JKBi�30V	�k�2Il��+�p�B�[a+�H��H^�-a�Ak����/WZ �)tf��UC^�q=����Ur~h��<��n&�D����.EA���p��7+���p�;�M��A��UoXc�z�rg�l����u�3?V֪j*�dZ�75!f�a,�.��UQ�PŎ�Ă������;��:��	}�~v~7��	i�]�<kn�n�/�鶯2��~N"Ӧ�㨟5��m5e ���AG���������|V�Z#�6F�|�&Z]A�$���l�:��wj�n1��V��*=�g���������&L�O�cq\Gu�M��U{g�YW��2�3̴�9Ǥ��q�(��?iQ�"w��\�k�h�2'ed�jz𼺅9�}��0��/������@��)�?WSR_��ǁ����l��S9� �	�f��-^�?��'MM�\��ӊ��g\�QY���t`s��D�9�ǽ�z��^֜�Hg4GbO�K�Ӽ^��J$�����͙l�g�Ym�-�R�mq�c�~x'���+g������,<�������vv7.�ڸ��wQr0�~Y�~/y`�&�]ը^����F���:-�}Fx�u�o�Oz^�&�(x�q"��r��풨�\M�h�9���ԪA���j�m��>'*�>���!C[q�L��a$��BL��A�Gz��q }g{sk��b�Y-d��s��h�.�Hȴ�a�bj�,��X��7Vމ	���m��>8��Ul�*[ʙ�!�]��x��6��4��X:��c.�a���.�Ψ�
0����9�컑�����hJ<�[���i�~���9^��t��JuJ8��h��p&����Q���;>�F���-��^,NyJ�V�#�dZG#	��f�,J�E��W¸�-��;���&���� -��䰧��� d~���7�|<��s@�8Ns{�,�l�w��]Ƣv�q�<J�52\��d%��r�y$O�.�H����[���H���f��xN�OfV�����\%g�ݑ��e��?�[���#.k��A�ES J�G)E�v.����d��ȧ�n/{3�꿗��>�d�$(c�P�@&��w�2J/nz.b��r�x�x�%q�����K��&�%L���(x�7��m�G�M��׮f��D��fm4C��핏���"��^��e w}��#!�G�+�-�����(=��WU�����~�]i� -|�EE��z;6.g��%%�������<��hˎ�����
כA��yƳ���O���(��	��͎��H�Q@�G���7_�,����|zf��
��YJ @3$�e�=K}gƲ^�l������a�O�4e��(%�����?��u&e+�K����|+l҄�w����.G��gF��zgRL��5N��xۢt����'j��f^�a�I}WQ�Ӎާ��GҲl"���Uxa#R���s�hē���SSNako����/b�7�Xfo�8��7�j����^
��'�w�L��6���|8��ۺ5/B��ΰ��.��p�z�R柫��ټ�VZgr~�e*���@��=lC�\�!4���6'/�c`���U���R�^����Q��.'���b�]��'���n��y�6�M��cw���� xie�Rh��KM��_��[���P}�W"�O�ϫe�*Ye=n�ʧ(�?S���=^\#NV��,/^ٱt_`���3H�wE����44��b�"�D`2��>-���?�|vy͙o�^���Dw��d�N^.��ک #&(�l �����@4P�Qm���;Z��[�	��K��ѧ���ϐƅ�5e�*�isPO��3,/� �CS��8��>1��8��NI ��� �Ԧ���ߘڔ��L�5�=2�Cj8)H�3I�PJ�b��\�F�A�-������)o e�(��Ÿ��|�|�x���H�Ҟ��g�/(����*!��d����g�Y
�2����k�,~�h-���J�v�v@��S��O�S�E�MѤ5�N;�}���`$���u��:�S�(J�1r������qFo=�Y�!V%�	q�Ǉ?���:�z�@wQt231ƈ-�����>6�X��l�B�),����ZA�7�E8��~!�^Rq��#/$F\�����d
'��ԫ
���7_-w��X�Άw�I���`�K� 6���=b�.<�J��Y-�'65� ���a�Iǻ��݁󨕖Y�/���{^͆6P�
��.H��}�H���>J��8��=�&]U(�n����*8ɻj¥3r�Z��^��"DHC,�B��;�� ��]�?k�F�'1�n�yV�	q))>Ћ�����W��jl��qS`�^+l6]�����}�0~��w��F��*�Ng�_pl~���`P�s�}�m�u@�S1�8M�	�vm�b�'%���y3���qT��8U�gR�67�F�=�$��nTX���/�)���J��q[s��n���A�����g��54q�ر��O kdӐ^aL��|f<W�)�=���ha�-��q_�©D�§-19ˌ�҇��\�B�"��;J0�G8&�ҭޝ|%����%PL�B��!���������Vtc²9�H�"��C0�u����^��k��ý���[=���gɌ�Z�6ߍ�)ұ�P��{�%�`���2
Z6E9�_ z�����p//
����X�B�;Zz����\d��&���mFo���boS���ro��ə[���fԘ2:�8X�ϴ��^�{%�I�MX����2j��M&�����-�j7ˈ�cÙd��>f�dB��o��w�$�X6��|���{��e�t�|��(`oLl�V����Fܑ
1��N:zxB�@�a��rA�ɞJ���@0���ɩg$�n�M�j������cC�;���:�K���,#�7�L� ����2z��
R���.�Wmf��wf�"Z6~D�����.r]�����$�� ��#���h��ʙ�D�Ô��P���_'s��y�N�.^��Cb�Ӊ�Oqc/�8��׿1rFzj���E���U@��m���KP
��$�vy�!=W��1���^T�op�oz�Ά�n����8��R�8mym8�����F\��	"8���$]J������E�F7p�j/����� 7��'h�^؄��N��:'n4��V�l�z���C���i;�0}:��Q\��ti��MG��j�����m�|5��D��t��{�C�csj,�<E��	��D�{XH(0�;�(qí�Z � x}Iv~��r�BW@=�P�9�#=v�w��u��[K\Y���@^�G�tf�S����x��sa���bt8�-Gb�{���+5B.V��/��(1���2��9�˸� �$���y.9��^a��T�oR�������mm�Ai�O{f���j�O,-Ųcvf	^�X͒]ꋮ�%���.X^���X^�܇�s"����{W�(��I���e>�-��FB�:�ٔN�0��^W/�S��W���ho �%-n��9:�E�("O�q�,8G���B(�ZF�WC��D��FW\f	�lX�N �^Ӈ9�"@W��*�p{�,���T�~�bX8Z�3h�A��PC�X�������p��2&�=�f��Y�؅�ǌR�d��8��+/�u�r��m��]>�FL>3h-�S���0,r�Zq�}�$$��
�,�9�*�m3P�M1���F�Ʀ�|m����ay>�h]K����c	_:'�{X�rm�e�v��jju���Ӑ����U��-��o:�IC3�y�Hb0�ρ�箔��U���0h"�8�wMۙ��K��S�,d�����DR+�������C�\1ƿ�Y�WFMJ_dK
��a��[��ؽ����!Ǣ�����d�`�g'a�y�@���]� ���C��9�qW9:U�˃c\�ŗg>a�� �~i��A��+%�W�טV��hFo�����s	~0zKX�@OW��G?*�����ƞ`�+ۅS�Q��]jp��:��X8���[��Ӱ��K:D� b��̣��s?I.���T���K��b��߹~��P���-V�����`�錵�q�c�n]��}Ḙ� IE�f�]W@��@4�~���%��A�		��D*��g���8��\:[M�Қ����I�Ql��jԄ�bMW y.��9X8�߇����9�d��,�L���%{�[*���b��3���]A̮'�,�z�p��tfK��:.���:j����$QM�!��W����}�Ӭy��
&6Q-6�[�Yd�'sRn�>�_M���?]U�S<���5a�`�0F鰴=:p�-���"�W���}�K?�mK?�~�
�\��|���빓�FW��fB*������vP+�6�I�c�L�1�
5��#�j�@0AQVF�݀�xn���x���^���F�������������^%|�Q��X@t� �ߠn����d^Sfu�E�)|���g[Ů����۸g� �F�{Jw4��y��K�d��(̎�&�,y���銺�A�	�]�e�>�d���
�
c��/lڴ�+���eM�BUk��G|�:����\U�*� �ERRX�� ���X ����^%LpŜd$<!��&'`�(b�DJ����n��	C�z8N��7\5�fn�f�\I�]CF����kR��:�ҥ�U��7�ʩ�����CM,?$/x��ow~2�Yz�}�;"����Bʟ#	R�1M�L���M�x���K�Ka��:�$�b0�k�G%
+7��y��q��x����h�k�EaUԶ.�A
��~��
�[u�	�s�ٔ���Z���O�ɇ��DKC�I	%�)�&p�o�NR��=ElI�{b�=���4�֍�;,��E�ު�LρWxOЈ��5�� ؗ�gn�hw��
%q2<ۼ�Z1�]�@@V�\���^:l�}l]�Yv���#ķ@#p�@�w��N�i��	Nn/WH��F�{i��<�q-a�.n�Y��;�.��xS��_��[��;{J���*��j�:p��^F�3,�6@��p�
�v�<x��e��
�V���,�Q!{��Nt 5��1X�l�t�X(ù�m�܏d�H�	�%��	��#J�J��Pt��S��Z������m̮���zK�`-*3k_h���!�G��5��3�CG	�&|���;�"�.��v�����Vc���v"���J��~���q#3�!������.\{�`>�=i7���h��*.�����j���QL����Ӧ�j�����D��QU��>�3;�o��_�$�H�آ�6���y6�B����q�q��]�[�Z�:Q���/=��z=Z�uG\�ݗٛ��W&L�5�ݞr9Hc���r���hR
 �X.e�k�A.�j�F����<&>#EK��󍴦�4�>�.�=��g�ߚ�i�
�-�GG��&�b��1�0��IV*gθ=Z�N�)��{E
Y:}�j�{�l�оY�������a����&��8������ڗʖ��7�C�NV�dx�q� ���Byڳ�:is�/-��V"��ɦ�����`�Դl<`�s�Hs s�n�*����%���In�E��Z²�������k�oc;��$G�,v
}��J2HN�y�� W���=_���ԅ\>"��W�I������ö�����j9V߃��#�Ɍ� .��
��Y�K6��U*�uz�YL�h��9 ���Ѻ��#��O��:I�ʄʎbh�V���_eJ-<�p�-3������mz�ʄ�A�B/c9�S��}q�?;܃����I�p�Z��l|ÿwȠ�
!���b��z
ǈ�!FY��7��mY���Y� X!��g��:�h~��,f�|��m�i��J�ґ���>���͊� �f���Q���9[�*"@��O+�e�5'Ws��c�u��"�G3�r����UP�f9��mT��׫�Ms�qh�OF3E�@��qOy#0����ZL����T�|��.9�5��ٔ9`K�{�BI((E;(�����������Uf�G��{��ԊM���s��8 ;勔;ⴎ�K$,�G�����=�_��EU:����X�0�_� ڐҋ|AC\���y:_�s��SV	�(&铚r�׌��^L��65�l���5P��d���蟪�``���I�թ�6v��#�%4��P�7z2d���[M�d0��	�#��`�{���T��P����R4�#'pc��`����A��
���\�YY�_.�
'0��j2���� �)�C�)]Gǜ�/�V]5���&�B<V	�rk���gk�/՗�vQC2:���-�����H�M:� 2r	���d�Y	%t{	�-��ct�:yuY����
�b���_�": Ʃ�C],¶#,�ׁ4���$����ft==�dYi�q3��6���F]l�?�E��BL�e^ծ1ɵ��(k+��,�ü���W����X�ӏ�����s���^ŎK|�mCW=<Ʒ�]H4;�20���\�&����^�5!kG��U�!�l��H�/w?R^<
E	%l����f���T:�=mI�V��*���ap�b^�'���b��t��O��,P��
f��lL�*��L������V檐c��n�hBIw��M#lֽA�*q������kx���%{���aI�0��9�5�6�t���[�9�·M�3!��Ѝ[�/�dw��y���S� J��F:�;1�8�D@�����'Uc�Q4k�҂����P��n�������}b���'*�=�t��9�����Q��b�Uʠ�{��0��e�;���5i�v;VLF�,�[Ot�9�oL�a�Ft]i<#iQ�>5�xN�y�~} C4���'��w�k��%�z�7�}W�N�����ð�Qr��iP��8���������1J��E��s�����u��艨����g1JIl�T*c#�Omk��9}�9� ���`py�+8�����K~'�yD�F�,*����*�Vz$���P�S�_蚚^���`	���|LRfr�O�"t�n�bC 9�o��(]�U� �tz���9�|t=Tn��F�Ʌ�z8�����!�)KpU����7��6� ��\_�LO�C�R��~}����0Ғ�{�B �2Ғ�:I̙K���9v�)�v��@7sa�Ȭ���}U6m�X�����ˉE�L��E&���=!C����S��������a����!�G��s���o���zR�1j������8$'f"��(���['Zf충!o����q�k���PAs�n�; ��Cf��y�3"
�BuLD��L�7�A��7��K��D3ek��+�D+�����e���Z�D1%-�@�<��3�T�0�S��96*��q�H���\��bHN��U�# ����dv�$�y�;(�d��5���n+t8W��I�Ի>Պ�DQUy����~Z���g,����0��HTy�_̀G���Z{����i� �Q'�3���D_��j�ü:mW7 ��+�uBŕ@^��Lq0dQ��Ehi�C����pM��Ʉ�/�5t�����'4ˈ�4.@�ʃ�@�S��D6��a�ň[}+\8�^�IE7���Q��(��.���K��2�4NܪE�x�!��t��$*�e�t	�-�¤�kdeџ	�%֥T��!Xt[�*-�l�Կ�o���DD�ɞ7�mB<t��f��ꢢxf6�^��v���ML<lh�#�R(!]�s�E��#C'+��A����M���W~7G ����y��1;ڐ�H�We������rQ��-M~�Eg�& $�3���},T��/�Y�h@c�J�p��^�]��f������G���B/�C�K��HL�b�t=�oLhV!�6�`$(ר?md@D��?�U�Ԑ[���>�)d�MU:�׌�����z��Nl`�TZB|��g턕�4���d/���ݚ�c�rEv6���%K�q�:���6�>k/j���-xFJf�~����]��$:��&�� �3(���S���:OO�5�C��Z �ؤ�F4�bS���ǀ�
�釵�3N�ՠ�驂�cs�όj���Fu\r���Y:,wN�@2�C,��^���@������Ɉ��@TnS5I��-�����җ֕'a�I�-C�>�zc�d=�|j���>]��LCk�f�s�$!�>R�$�J���\�f��<y�7H2����9yjGyT<�B���k��J7����L,�C�)�@E�G'����g��*�x���ڔ;��J�^"3TX\M�)��}3'��rvhwZG��S��jI�Y��E�'�D��6|��1?.��,��04�Iŀ���"�,�$j�,i(h�T�%u���[��'�����E��A2�v��]w��EFMp���s kx�#_���}����0AC��{�A�����n����W�Q&*��/�����yњ�&H��e=����>O��a������A#����4��3��m;�d6K)0����>�9�ݭz3�A���E;"Q��n�^�p��&��h�+�i��@��ܶxء<�i��m|��(�����+�j
���Ï� ɝ˃61��`���'����s��R�+��u�{��+�M��t�'V���M�79�a��L��G����������Pa龸�tU�F�α48��*���w*��Q����\#��RQ���h��{�H���x�o?�9��]��#L3�o���ç��I�Qc���vV2u���8�q�-ƭ���;*���G����R��xSb�?�x�I� ��G9tXL�ӝP�F��K��u�z����׭�0t��~�
��
�����v�.c]�!�9\C���|�+vX*�LY�A}i���,�ˍH;��[�����*�Հ	�Q ��W�C/�~�A�'��/�'��sܾSc��Rb m �����U�<����}���4�ŗ��|�|���CF���=�b�a��'���pf���=!G�H���B�f�����&]5b��,+�[��B)/�[�����;���|��Hs.%�����s�?4��^�0���?Nt��g�S"J9!��s_'������EUsJ�[e)�p���t�d�@Ǿ�;��O����W9�	�o�!W2K���H*��u���A�q�7�`�����v#6�H�i	��A�Xl��9��q�+���?;J���O3E~t	�w��X�jcƆ�k!���:�{ɥ�X�g%�z�Szύ��J���������!?r�;2�_�2������(��U�(��
2t'�^��{3'�ݜ�U��x��C;����@o��G��JF#E��*���N&wco�(���2���2�iE]��i�
�Q?(!�9$��½�ۅ�G($�͋o4R��ɦNG$O����y�4ʸ��\C�m�q>���=�,����Pф�,��h�c��������W� �0&޼�W��h@��y�s�e:�@�V��q��~�]ʣU��B閘p�]�����~�������e�Y������g��2�zpX0�	���ho���tt���Tm�iB����P��eƪh�Fߙ�[�"�Ѫ�fWwj۟�_�5��I��u���vq���6�P5�2�)�_؇ݠ�����1�!?
�Ss��F��39;^�`�.d�_z�(�֧��ŉn̔��$�����������$�ct��O���{a\�VdUi�}N��?`��T�|�1����3���
��e��w��\����xOSf̶�9���fL�WrZ�:������D!���ז�r��*��4C)�N17�DQ-LE/9�r~�KG�D��#�_.q����$0)����z�j>?[�JO>�7<}�kŵ�����s�P�5u՝G定S��U־�U)�NB�{��糟)�Z��(�����T?4\c\��o5M�I�'��N�K�/�E��۶P��8'[ۻ����?� �u5�Y����+M�<��Ғ��m� �\����ƎX��%�'��K�ԹT�Nw��z32啡��y��������Fg�uPY�t*���(�Pd�}��0�1�`�C�}�<�� ¬����`N�����C��r�(�Y�K�	��E��2U�U�iEs�"�U8N��Ga0>��ɝG�	�������4�7a,A�;.��k��K��2<G�|"�~�%���i��Y�Hm�P<�O��yn��]�0����+��;����Ff�>�^�l��ԇ�0z�՜4�̬�?��%Xv��X��;�
n�f��Z��HZ���Z���	rX�~�m#�s��z�A�G�v?xU�f��C�{�u8�'[��1�¾ ��ܧ��T����I��"
>��Ŕ�U���;�S<�da���cR�{08��!1��_:|�.$����?ўB��̰����G���C���wMq��41
���R$�'5��xX��.�|�b���y4u������)�k]WT�JZ5u�0'I������t[����7ʥ�~e���Kcu�1���6�(���❐�}������x�4��W[�����҄zP��Ɏ.ӄ�aNЦ��1D~K��u�*_]	s��tߵk(����s�Q�.�m3�ތ��w�Ta#�P0�)����6�Z��3Gd��������9��	�:�k`��sU���c"��@��/���(�}0��	��P���ss���7�	�����]��/�����4ۃT�9yjbY�k�L�����8be�+��z`���q��'HTh0D����d�+���()��5��pw���~+�ɬ޷����<$Q-^�8W����]�$7��9VM�~l]��'��BMρ�Q���YW�����u�Fd�������?��I
ݕ�=O�É���nGuە�뼟7X����Y0������)k����s���BM��Sr��Qc���g���r�Q�򅫙���S����Yt����+ٛ��Pc�ho)AԵ̐U#��Az�xÞ��	Ӭo�n��s�����a�%j����A�1�~_7�Gvc��`&��>���7�ד�Kơ<O�"Z�|��5F1��A3�H?o9�mS��Zb��l
��*~��Y+"ѧ��-�Eʓ�9�҄9�أ�<�7l��#A7����G�L]?Ԑ���Pz�w�o��&o����;j�j�8ۭ��J��y�_:���R�hʊ�%�E�5\��`IkU�������/ue�`?����Q�g͉x��>kp��
S; �5^>�y�X��K
?�7���h��*�˿-���C���KE-����*cf�|�0r�p|Z�9�� ��(v�y�|���I�F�%�p�ʉ���G�;�h�)������r���qW�c#�0��a87>�Ԩ�~�P�Q<�b�3"$«�Z���>�Ш��=s�S�a&��s���}�l�$�e����Uk�Y�	�ő�Yp�O��. u�2�\��6"CV3Ŏo�O�F��M�1t�j	�z�,7�����=��!�P�� ڼ��3�^%��<�8N�쐯�$r����Iwv�
{u4o���cX�;ASزLBUˆ��˝,���P=��_j�N�h�QFa�1sf����iFK��7L�Qw�m�k끪��ƛ3��P�������'��}Ō�ފ���<v�O`��}O�������B��]�$1Q/j� ig9}g�tF�Z�dw�¨(�.�����E/��x�%�<J���B����#����Y[`�O�7[v�[P�#{��_4����K�OΩo7��-�����滪��)Y
Қ٣ry��mJ��-���A��ׅW�����Q�v��@�� ���{���c�z���&"�����OT2����׆ҪbV�l�D�l�F۔{�ԅ�\�'��5�O�tC��Ô�ub���	O�������h1���)5��W
Q�.�~Φ����Y78�������U3ce3�?_�
�q ������~�p~$��v��cn��f�BY��5Q���;�����tn��QMŀ-t���Spy͠�S�3ȰKZ�K�d��W+�ʰ�)�
���h�{NJU��!���F��4�xd�`#eΦ��W抡�)�!$-�[�Xv��f��7�����bd!{s�㫱i6t<�X�Hȩ����:M��	2�]�UP�9�V�HF��)zy��]�b��2]k׻TgR���ɏ�ėӢ_ެ �!��6l�!Ɉ��6��Pn��C0�;UM0�
x��L�}6����x��:3U���>�k:r��_7�$_�#� }�@��4|77߳KuЮ���|GM�b!G�al���EP�O��j�^�#B�d*�P���&���az���
�έ@x"kTd�2�yVU���ҵ��Lzr0E�B��
zޣ��ֳ@O{��j؍�8Vd��F�������w��3��Du����U�V�j3yY{z�K��w����6_C������ߧ[���n5fu��>�jF�0��쮘�	%���/%*]�B�C�������y�S.�&#��b�����P΁�<@�	W&�a�͖ϻ�Kٶ=��؊<��-�op
�x�L}�,��%& O���6���U��=ф%x](��VT��ҥ)��ed�>�2ȯ�8>M�q��?�����S�,�at�{�׼��E Z�$�`}8��M� >Y>�FS{}K���shθ��v1�#�7"��k�=���U^;lΌ$С\�D:&��X�&�=LG��.-J�\!�[ �̚w�E��V�nV
3��-[��Q}�gn�V��Kdժ�I���;�]$GX	P��9���}�$�*��dɧ�}��
{Z�|��=X4��vg�Q���FS|YcOep����8������c�Nd�m�X��J�#����|�\������(�1W���w�s|6��8��
��(���ӽ����:#��+}3�^�x/q7���R?4����õ��(7�ǫ��u�2X�KV-�zC����Auo�d�1 ��~�n&��
.N��b��e���<�grϩFm�x��%>i�ҒdP�&G�Nf Ɩ!��.kJ0w�%�lI�i� �\��>U�,��Kn�Urэ ���E	���A�!w����.g�9^7>S��T�.I���58�TCW�?�Z���uN���܍�HY�A���qҝd�C�w��R������LݷU�{�_�:B�)fx�� �:�=�u�c�Q��Píc W�+�"��-����[j4E�;N>)z��0tV|�qL���	*�NC�_k���m�~#�;�Y��"�`��胧�k��:��.��U�(���g�w�>!�����[��@�At�����O�����0-����\A0�K#��G���U�Pk!��;����l�fIj��|Z�|B��l��&h�|�;��l�ivu��;�.��� p!ͱ��-Is\!lB~�1����8�Pu�eh	� ���|���/ո���1�z���a��<����!O~�o��H�5��,!$�;��6���_(!S�M���2���ᅇ3B�̾z��L��^��J5��M'�)1� +�3�|V�j�+��^��s��Z��s���!؏*�tO��6��ȧ;nA��c�Q�X����	y��OUtTI�����b0��3���P�TF��&w?�j:og������d����MP܅]��3�rP;H\ނA+�˭H�;�,�[$(� �瘸���б�_��)� �f��� ,�������}�l��=U����U =g���[2��Z������F�4�O����޵�gg���]IJ�A*̍�K ���1.g+3��4 
�(������!e_ބ.�K(�QB�i'W�^l���W�(�ծ��M� <����́-2j��/���1�7@������,�BQ�۾ݹ��w��tO��|����3�#M��U����/u	N%:<%Q�Y/���������Vv��e�gc�i�:�C��dζὒ)z���_i��)���l������aʽj�;^�w3������V�BDze����r��_d|���5��R���X��<f�sb�kk��d�#e��.SYO�J�'��u��'�&:��M[�3Ȯ�ٻ�H�Ɉٸ���G,��1�g@YgC��P��)��F���i�ژ.xEJL�r��C���u�bLf�}ɏНZK%&2�Ñ���H�$��Kp����3"�S��Y�܉��J�V|}��?��?n��� X���%Nk���Q�3a��h����꯾#�$�D��*��t������G�=9O��}�(�z�>;�J��JiH ��:;�p�{��4�<V�A��P	~$�,�nz�h�F��\�:�%��XO�?fb����-{n��<+sF��_k��F裤}یg�.�� w�XI��uR^~v��T��A�h?�|&�Gm�1U�[u��vQ�#J�Y[�]��^��FW�iy�-��T�[�(˾�u��}������B�U��W��؅\l?��o#���W���b���@Qr��BK:ĬU�f�%F���{<ME"�[F_\\���{u�"���#DB��"��
�D��E�ς(L")l�T.8<�d}�vz�]���2����PgqŵR��eZ\��o�7�quF�㯧��3�JVI�U�pZ��'�8���L��q!����(�h1����,��8'�i�9^Y>m�K����gS���:��y��~5���/��۩h��~^c�z�+������z�\�&�d-����ki�;O��Τo^�앏- ��yL@��ilqК?�)1c⢷������4��|&`�?��A7r=�9��n���˕��16��Sh�Ϛ�6�2-����OQK�![qltz">]
�WƁ[}!��������V�Q�p.K3���W��ͥy��M�T������Z����B9���:;�4����3;;�y����%�@k�:R���+2Hh:��!&��B�I��T���O6;*|����#u6k�?�1cd��1\��t)7{�m0j��o�##�T7,\|i��o��^�S��u����q����]sFhcrx�)�H�ЕC�"�DE�XL���z�^�f��yG��.����p�Y9*����M��{R��UEx7�:�U��^;鬳C珏\2.�M9ӆ�en�=�Cg�󹵘"���W`l�&��	%����гf�4��%��=�z�r<�{|��;����t͠�$�;.���	�Ǖ^�fA6��x�� KG���j��2��c���G2��k�	c.���9?��z���MK �Mo�-��F���,m�ޒ�~�=,���wlЈ���i�w�/� $�S��l -᝺����sj�"^$=0�=�������.-CT�^�I��oᲡ`v�w@�ʚD���=�i��i��)�;[��3^�N�6+��2�q|�����3��5_vL��,�GBC���'jЏ�TSJ~ݏ�0�$[b-ёo^X17�a�|�Կ��F�1m����$�V��>l�%�0����d���q�>i�[� �=*Q;�eD;Mt��l%��h�5�K��g�[GL�������e(pеt�A@��1V#�ݲ����3�?�ͨ�P@�ڲ7���)�~^T�˚����%�.���<�B6����8��btݚ���:7٪�����^�^+T-�ٰқ�{���q��g�H�XE�;s�����{��	�G�.�1�����'R��Rq��Ї�)����,��&e�NM�"*KM����`����$Q��پS�:���Ӊw�s��:)1��VO'�n\���aR=M�/�D���H�,M#�;�[��]��zM}����NH�Dz��S�����$�S߀s�K(�5����hG���}!���~�=m+
��8��H�>2�$n���k���Zp7��gq��+Zu���O�MJ�E�������憑/Í��1��x~�{'E�1f}W�ȕS�:)g�xJ -�1c���ɈZ��g�;�*uU��ڟjZ2s�ӡ�N`3��=��SR�y���o?"����|s�L���9\�붌��
lp!XZ5\�Mp�x�Hź�ۯS���n2=\�0�»��M��2t{�O�)���AĹ�'�֍�h�_e��cm\�������#�8i�g�����@o���/�ա?Q�Ś���2��P{�u�ExO2�|�s[_��Sǣ��Al���@�\����߲�	�t>Wf�3��ʾI��^߿2�3.��j��ڳ���#��H+D�~�%��l�8�ԣ�>��hG�v���5=}�`K$%k�D��Ζ��6k-��rF) �ո��5�	(�4C'6�V�Y[������Y�2m��s"���wpkśq����Ȳ��D��Ym�)Ȱ!f�S�I�o����U?�����`J�L�⳵�j~?5f��9�iU��6a��r�E��l�4�5	Q�B�m������m�L�d��T'|7�G\��&���KU#r�	J�T9D���O��������I�P�T8A7I��m������i�U�ĐeD^�g8�)��;oPt>Oёmт� Vx��P�+��喘�b�������<we��O����$�@��2�����r.��$r��͟?N���I����)�b,�2mk*�,�t��ׅ�8xY,&�Sý4I%��}󌚮&���%��j̜�h���o������
u�٨��v٤U���8�:ՠx��l����D���a�f�+	 ���H�b'Ǿ��)"�|�0>��X�s1	a�G/�/�ĥ����M�݁J�������£�＄N�:�x*��!d���ScaD������2��"�oCud(%ݖ�g��{���G��D@�]��+0�1��߳2�b�8���a6��u�U�2�:���<�[x��+�fBa�"�|�X B��6��u1u&���:a�R$��]� ٚ���ӫ�!k��S����J�~?n��ec������E����\�KCå�';j�i (�t	e0A�O��`7P5$�v��:b�0�6�l�f2]{`�h������i�8�T[�DmH���=t��Z�z就���F]#u����Ϣ��d<�eO#���K�$(�g�Hy�q�Ns, ������;�eТ���5����i�����W��Yj���H�����cGQ��TݥMAa;��R'-��WL�5����9s�p�!�?�RKrK�E�}�#rNt�ފ�=�|į���\ϧ۹*3R�5t"&��9�P޲f��N8X�m��b�]..�<b�lj��$v%f
��.���<׎4dYH@�/��\��2;IƗ?�r58�!��T ���i����86��O"��R�y�x(;�6�C��� ����D�A��e{~[s�9��ϡb�6������@Z�#kGYy20�O8�| xg�Qg�g�|��}�4fڏ�њ���6P{~�#��8�J���6�}�V���bZ���'��� �����-O���o�WQN�i"����	����@) ��=���'�|��#���Z�x�2��S� �;^�X�z�{��ᗂ��<�:�y��"4ϱ��n�0A���)�6�L�Y�J�����w�VG���_I^��"�m�rB��(����{;�Əo�箜B׬��}{)���F�aW,J2��ɩ�!�O��;$MO;�x{�c��D%K��c��?�%Ѻ:��ȃ�,���f�'w����>-��M��?N����g��y�c�+�дs�T��mW�>�Zc@0+SP��Z+5H#vy�=je'��f��Ƙ%�Jc[����5q��	}1vL��Ƥ�^%�q0g.?�'��k}�̷%L�j� �_�!����Y����0S��j� TW�����	�ݛ��`����O��u���R���������l��K����;���Xn޵SE����%?9z��3X.i��r���*��	��U9���*b<b�;�h���~D��3����>��Vfj���ʻ�aYϥ�!�R�E}F��((-�o��D�����&[K$y5͠V4VE�s�3���<���`O4��/��<HdˊU�G �0��v�L�6($@�x܊��?E�K	��s~�� \QI���O^ދt��$�9~a�N_�޶_ei�Q�Q�?�p��@53�t�hE�����6����d�%�~֗��z8Τd|�	��{�pI�dr�I�m$�<Y�=��}6m��@��V�Ɍ��y���S	��*���Q�&���5bk��`{͢�����8�AZ0ĿP��r����\������*��WIn�ڡ�ҹ<X�7�?���GΒ�H�ݪgArQ_а�_���әߍfW�d�BV�P�~���x.�_dF��hb�c��1���C�1�A0gv��X�PE���Q�悒Ԋ��hs�#(C�:i�S���?2Ж�-9l�����R�{8�]��l��b�c(}�}8P.�&oD_?C���<��Sd8�kB|����Pڡ��2���M��[���ȶ�?�UN������#q���hq~W�3I��	W:N鉝<�LG�b�EFz�J�۾��3G=��D���,�&N{��6�&�05��h\�Ꟁ�4�#|����5H�<#N�'���T<�^�#�f����0�|����ڂ�#J$�Ϧ��o�K���x�\�G�� �������;��EY��r-~�*��ɀ�
j(~nm������j��	18Z��@Hs���P4bmVg'��W�a[�����ڤ���H�Q���	?�θN�+l?������w����V���NS���Sg`�y)\���<���̟B�
a���1�����������9kn����n|r�����3�绊6���J�N�m�� �!�<,H�.mBy�PD�(�$d��&*�d>� 	^h��L��Eu���E�R�Dr��d�Iׄ>�:i����K����R��ۥY�[zj*���!2����^P�l���^O)0��">'��Ŝ���$}c�!#�rB�.��b��U�"��d�*�G~�eo����F�H2��2��qM}��q"�T�+Ə�0���J;A`���]�7ͻR��y{:7��p�}5�r`�kɩ�yK�a��w��,�GK�C�q<�'�*"�Al)b��UL������ٮ%��+TJ>��Jz��!����x!tN�4B�/��,Դw�Mõ�b�M�� ��b�/�q��1l�%s��z���;Kȅa�����d>t�l��}�d�I�D����t�+_�s�}���2�	Gj�Vُ����k�>�>Z�*�]�@��|�N�IFQ"���If����V޴���l�ej��ǎm��칳�T���fg����8�Ǐ�t{�ہ�x[Oo]+�n�L�v��\뚕U���E�'
H��"�K ��(�K�"
�o�O���P�����5�#!jO���E�9t��A��8m�\!�X[Uݫ{�X\��o�@����j��	��I���+��6�N�>`n�>AF@�}�w�ߒ��_�x�G��uKa"E泀V�)�DC���_��3���=[�ԉ����@�w�v��BVq��s��8
ql^ISY=]= fw{S������� 1�F�^��7i�xg�ZIz4DD_�/wO9��S0�<�x���A��|���1�A]�]w<��߼�SUA�瑣����>=7��l���N�O%!��r�N�`&}��0)��"��9���)3�-K���w����f�L)���Tǰ�d�5L��E�Fǒ��m�2z[ir����t����M�-��+�	ю�$��@�^�@j���YM	�8��0�pg>�*�^>	�?�L	.'΃��� �l.�롬*�:�d�!�6�L8�J�Ȱx:��3	:�bC����Q�����}?z��u��|��H�?����h$@�g�ޤ4"_݂�`���SwP����q�+$@?�bZ`��������t�e�6	�����)k���J.Φ*�oy:Ea��#�\�0J"�n_-Z<q�|�$G��+}�e���Q��ʶ�p�!��Ls�r|*�b�~�v#>�S�!ư[��gV�c.��S���(Kӄ�NZTRgV�n3*�-1�����qvU�yTS�ڋ�b�OQX�қ]�m���s�A$hpFN�k�U�%���0�}P�������֢w_P"�y�D��E�dgG�j�4T�Dx��y��3L�n��i9>�^���|dO2(@�f3���VB����4R��%��a��0�;�p
O�H3��ѲƬ�`���M��XB�8gZ�[<��;�cn=����+4�,E>�� %�=��"mx`vW��$�u�HϾ�a���Ź�	��r��m�f�����F))����!ya|g�����{>��/�@A1������#�	@�n���|��+f$}�g8p��$rs殈����^��,g��N坕j"# ���>��|e�տ��5��dԺ�>q�ZGk���S���	ڙ�];��;X"b6�,7]ү�����̹4vA�]����{����I��*�nw�J���M��][�jY�Oʏh�/����{��Ήb����|n���-����'F�4����8�� qU���(��E\��mQ�TQ]�M���>��. fmZ����r��۝"���GS�������Ϭx�hes%W��J��Q0��O����6�3�\��2q�Ƹ�i�vZ>՛�gr8Z�V��a�z'�?N3����0\@o%��vk�~S�B��1�����E��c��Qa��!'^�B�K�GƲ���l�z���ADs�x�.}�[d̻a�,e�1u��/q�u	�<�М��:�Vޚ�J�:��\��k�z�M�V@��n{�&F��x�6z�բV[� ��ؼu+��~o��	0%�D��-|�v �zc��~�CUI8����?~^`w�$aɏģ`f�F|�j�r��~���G����7L��F�����}oh��n2��C��a!h��M�h����uJ\M�\��O�sbns���O�e�˕.�=��2��MH���O%w�_���9����i#�%���taD�O5$��b]<S�ǫ��Ҙ�V��/��P��Wc;y<�:������xE�A9��C���$��kd~�"�)+�!�B����d��o�F�����x�%���)�S~)�&��-F{A17�,Oǁ���Au�V(X�=��V��Ϯ����7>�g~q�R��Z��vr��m��_��h�;�	u�V�Zp������z�H�=�?ٝ��q����<�R(ˮ�b1�c���䊚N�����ޔ��і,bS������@D���a���h�������$0L���3ܧ&�c�7"qW��"�P��oTd���M���S*�1P@]�P���j( ��Yh�r�� z��"���ew�b��mS/��$�*��#��T��9d(����M����!=��K\�؝�Q5yv�*\r�Ď��vN=��R~�s~#%d$s��:���Y9 ��`�a�iL1Qt�J�=�����Wאc�+�&�/(L�<�s����g��&oAC�}@�B��]ؖ�_l�MK�ޡ����#*�ٺ�t��?y��t�h>�ϛ|5�>!E�(I�s���:{G��A�D��W��6Mh��s�r����dF��~\�ڐ�k�Ṭ-E��f	��� �����'�쩑!+�l�Fg�'��v'��(;�̛�� ��Y��쩢�!xw[��~�G-<~An��t��1���Ũ�`�S��@����hX���s(��)�˓K"�z����
4��B��z�(D��y��*��ʾ�mu��ച��/��"�Ì��,cCX�\��%��!�C�C����],�{��**���5B�̭�����]������j�p�v�4Z�+�Y`�~�(�&kD�R(T��X�Q@���#���]@� ��"��F;v�]n�ChA�M���)���
�Æ0+4P�ő#dj~�d�kHI�1�������t�H,��2����f��g��/{�������O�<F�x�� �l��Z1`�SQw1�\��-=��n�K�Q��M���ُ���,P��@?ϖ}�����ŅS��MӉ+��}�c�����b\�X����Q�����^�w_5��D�g4r�AV[��-�I�q�P����ٳ�bH��I@Aٞ~��+jZ���� ��Ӎ���py�=ﻟ���V3o��0�C�#է�ϷW��v��mq^����5����������0
LI����j�/��)?�t�d�~����K�ȁ`�ەHV����~��း�7��G_�@L�!�kJ	�]���! 嬝7�?�}��c�����<�A���g�PmL��n���炁�Ifd�7h���E/�b���&&�� !�,�X�3%�$ .v#I�]r�%�KJ�T~~w-̓d��~�>������U�ʏe0mP~�çݤV��@)C�� 4�?4jU�Zȵ��8��Cg��S+���_��CSK�!f��"�̒>��^su�
YgYP�g����s���1���1�%5�\��-�V{�l�Y����\S*�~��iQ�7y�@�����JPK	�I�R{T�l�	r;!��C!C��SSH߼(��O�>���Ѣ�U[v��M8�^�M?�ᣔ>��ʨ7��a���{�b�T��QU�cE��TS�(�,���9������KT��d!:��_���p�gT��S��Źc��$ߞ�ڕ$T�-c�=m����!^���厑�H��gX�d/C�0�̺��s��0��j�F�%�GNU��q.~�Zʝ�0����b��xK����T�Il%;#�?Fd���B�8/>�V܅%���p��i=�U�ݿF�mV�ĥf������'�MY�K�Z7�n�I2�o��4'g�����mI,�=�Xݫ�2�Q�c��j�׉�d����)e��|ۋ����{)��+4�V�&��k7p",�)Y\Q�Rr�j���>L����)y�W���\�%<"�Y��rA鏴j���C�Y~�5�N)����x��n��S��sR�8���wcV熇��GO�|O'!�:""�h������Av�%��d&��$�qèH����'�XyZ�yv�5Σ&�*�x��D\E�Ģ:ml��v�	VYO���x,i\����m)Lc��45��:��Kb�@��nE�m�kRR�Aa�!2�R�h�\P{���	�6�)jI�>�\�@H5�s��R��^�5&��yɄ�)W��a�:�����i�7�Θ^$5{� /���X�Mv�R�8�z���8�1]h~yZ���ü��hl�h2j\�+�u�6��#�m)���ZA� �w�����Y!�^Ï�k�N�&
�u�R�+�<B�c�X�#g%�"�T9��`�"O�,]�+�"W�&lN�R�Ǣ�|g��Z�&`g�s��M������qn;��	�n���\��YJ�������v��A�M�ޏ���"1�};i%��97�����m�F~�`_����}2!������<�.gE�t	*�wʊ]W�I���124��<�2�rh�]�k�)���Ia���FH2�(OS,�*����	<�n�����������b8���:s�"��U�G Ǭ_����������Փ���ü��Ocs%c��}��KwL6�tl����8=$W��[d4�Ҕ=T��#�C��cTM�$���!�h�{?�7O�3U���e�{�š�j:/hM,�m��+���s�>w��%�4>�M��TU3��vl��P�R����b�����l)G�މf���ER�Ӛ	a.*�c!-��f5���-<�X����A�M���s���j:�~d�ɖ��.��em��)�{�s	����G�=])W��|��)E�ݵb��>7�]ѳu�2#����^���{�?�Y�w�j3<�vR����IG����-2r�B������&'<�YG�H6���%�mI��7���:u������M�jb�d�'!Zu�%�A��T�M�v�#>�T���ئO����r���m6>|'�G�)��%�����Qܒ_����(˭����w0`#ҵ��Ջ^K��c�덊V���q��>z���g�$�7%׸u`����'��]b-�Y�=#��t{}I�f),���ã�%O�ǑκWp듯4>o:�*�io��f�n����RM�9�G�΂[IX���R����%�'����vc�y�-�j���E�=�E�+Z�F��b)V��W{E����"�11�F^�g%��{��|nt�9����/��D��Q/X���Y���A��e� d`��k~�j�؜NB�lNC�	�ظ�(,�Nꨥ���uۗ�0����!���ӑ��pӾHV�UW��9�Skh�}�;B�"5e/hE���cO����3���W�|��fI�:��8W�A��NWcD�5� R)]:��
���%+r�u��`� ���a�&b�נ�1���Τ�\�}���#��9��'�jR�ǲ��@;d�e�� �������ǭ�.@� v�;�D<l���D4�gA��t�g�Ȑ����ݝ6�WE�!��m�8gt��/EK��v?�P.�Ԗh��դ���ISNfO~u�~V�Ý��e��C��<2�jư����g�F"bDS�5�}S*"�O�6��c4O?.e|ծR�܊�y=��b�@ɭ7%��*�!�H��}o�^͝��H�YEf�	���=����?���)/�0_1�Sx��iʹ����N`��I�Bٜ_?�S6@��V=�a0�W�Ԁ{�"�OP��ҕ1��.�.��-����C:�"s��c���a�����������ttGt� ����+��E��ԁ7k��dgk�� �c��0��|�t[֡['�++���|��]�ī��F��Џ�"��t���E;Z!�U��k�N��nm'Q=�8�t?��ʐ����;��P�&����[�p,F��Y���M*���e�2�6�$wz2̏lP>�K�'4~�`���o!�qg�Jt�}xW�}8$���E���BYȢ�M�����~:v��R�%��x\OvF,Q���=�5Hh#,G�u�~�3�}_0�S��H�^�m�:��� oK%Sˤ�N+ɰ�����:�!��H�6cx|u�zn�����R?7����'�潦��8K�z?��D~����b�=[$*v�=�|0���I�	Qm�NT�u,��M��N煻9"l�۴||R{�S�/j���@%�Ѣkj�s ӭ��hF*G(��m��C�Eq���B��GYl��<K[	�2��Jܒš,���1gSP@� T�Y 7 �H�ny6XG0�����2|�VN�oA�9?������'#��r��u���9�������C8z�'��k�܂OtV��٤��M�?s./-o���b�8.^�o�u�0�i�O� ��nY{�-�>�h�����5QD�`yF,���Uź�o2�8ǟ�G��hY�6Z�e�{D6A�.$sw�>E�{��xz�ﭯ�6t�2�4��}��N7���Z(���X�����*BՈ�(
f��+��iK>Ŝޓlt����g%��
��	��L�H�W�/�C$x�iB1���Qn�[�π"N���+�e��V�+;��y}��2C20����a�<��Ì ]����i��ڗG��>�v��[7��jy����xь�����L(��r�k�9���~f^0�]����F�����E�R�#�
#��FP�Ӯ�\G���¸)�
ۺPC�VM�q�ke��=Ԓ��4,�",�'[?X�^�2�[����f]3�.�&�.��Gz�j`E8Hq^}ᶂW�}�^���1�ؽ�W��7����5'�=I�BOߤ��9�������\
���_s��Zs �/*͉ ��G���2(l���c�~l�~*f�~�P��k��1��M�������u�K���R��*����Й$��g�b,M�L��Y	�j��N3���H{��}h���Fٿ��?w~�~�v�_��B��2N�t�yئ�I��L΄�f�(c4���	冩�i�^/
����L�'����(�x���Zh{���:5c��%d �1�D�fQ�$]���ͫQ m�3+b\1�L���r\^�x#�
 �/X���]!�a5<G@
����L�w��q�*񇢱Q�F���d���"m��	C }���3��C����E�R%N�A�`�|h�|�Ft�hzV�cszB9���hr%�f�Kģ��Ç��8��ї�Y2�L%j���;×�4lR�YU4�K��a��j��O���H訁���{�M�ζm]�\�m,�q����:���#��J��ϛ�2Ƀe D�����%~^�vZ1��q�[�[�I���ëJ�s�a	Q�(�v����M0Wò�g(��9�0qS��8�)����������D�@�[md<'/��F�u�Q!��$l�_�"�6|ܣ&������x��w�ƚmN>:��c�r���H��@FWf!R�[�r�p��&��C�%�U��
P8~�'8W�3$��7����k�
�]4�;Dĕ<{E��x��Ud��D�d�F{�"�t*J9�ϊ��y�N:�k���1 �i���BAZ���'U#���?�o(\&�}Ἄ���*�h$�P[�`x�[�!��|��#��7	M��������B���FU��RUr�OQ7�J���)k�3pF f�7��ݘ�@�R�M���	ѨhְK +I��g������������ssm��s2��k�@B�Da��|�,���0{v���]<�F%w\tF��@�Z�21e�<&�U���(�#�##��:���v���G�g�����7/�t.����~�#��_L�A�v)ACer��)[��g�ot8Eq�-��h�8(*�>�J{�jъ��Yz�^���b�3C�6�حhI0�	�������3A���	���ϵ��z�}�3x�rB8$��`ǺɅx�,���
s``1�7ܵ?*J� �(��O/Rp8�
�/>�����Tx���si�k\�?V�^�ݙ�
"_(���V�,��7� ��~wX1#�����L5A�p�`;�p�-��H��U��)�VI6;8�;%��ä�g6��!�%@��]ۥ���h����9n���cU�cD���ɠtQV�. gރ�2;Nw��J:e�&+���axh��e�`M_��Ӆ˯m��0�OTu���bpG��UF�0��!Z��?$~>΄7T��%��M�W�F��^Z�CUKf��u[��Ɲ!~fH�r���
Ȝ."\{c=�C�����f��;o?�H�3�q����jp+����Όk�x�Oa�)瘶A�0�*l-e��R-)����xEΞ�J�� 6cDS#ù�7�:��AdkN�3"=a�HEָ�{�Ύ����i1�v�V�oϪUC; A�*j�aNRo5�[�K,�����`ȼ��4%��V���P4�Q�@�Ʒ�"��%Esg����C<$�vt��ww��ݺ�����}���韐���m�[�5�5y[�0����p���9�	�����KG���"�O�����$9���JV��������h�-+Q�G/��!0�E�Iދ��CO#���)"��O��!�e� a�rQu��GlE�"��!��/c�8��c���)U�o��)�����%��1u�S�� ������3�8X����pl�x�p;O��DL��p}k��X�������{�����y�;��*\�%�2H��k�a��a�]
�/�v5�J-���-�{c������D@���Pg�%O��wm�_n!T��u���ny�|/ �&����z��>e���a,f��K�i���p+�os1x���R�8�P[_e-��b�.��²�A�39�qO�������øW�x#^DC�em��k�����i���ۨt�(�$#߷(?�cM���F�k�t�^��GZD���2D�(�����2�&��4�����&`���M���JP+ �/�9��uyeeA�HMC�؅�[�B�$���5%p�Od��9��Z�_�P&%	�ձ�%�M�}��6�n�~��(�o�����1V,RA�,�ۖ�[H�1�������nj� ��@G�f��θG�b����"KϑBWg���"������sz���4�S
і�{�1�#D�ކQHo��ʚx2�N�د 8������I4MF8�z%e���[/�_%S���\cl���H��2��������G���j!&MZ&U����9��g���\,k�P�QF�A )���L��E�������[�w\�"�-�)-[L�H�y��p��������������!F�a��k-+�d ���sau��:�g�Ͷz��ij�1��3�����q�bЀ���%a ���:�m����O��rf�e��'�Z�n\P��Ć�3��8�2���^��X1&�p����ѭ/������R����d�y^H1��Qe�xM�o��`��v�xu��!�F��H�b.�7���L6�v�~0	�"��!qg��^Z��}I�C/��U���?�vq��+�M\�l�7cd7����|��|,��w0HmP��&�Fl+��D��>�"�U^	)E�uS�tho�16\=���`S��ͤlR晼�	���/\ш��[pm�]������&T׽�6�P���2q��,�w�#�k7���e�w�t:kWn��ԣ�[�X�@����vWoqۗ�_��y^yE�4F��W}ӥ�:7��a�XwA2 �'e��Z�l�U��a�,���0����Ɵ�	滲o?��ߛ'���?��\��;�gϚE�A&�Z�zHW��ֈ���t� R���y�O	�?c�|7�b�Y9X!��ʦ�+�~*��T�¢;��x#�aP����l'���h�h�a���s�>�^%��t�ˡ���,�����\;��	���7=쓝:c�צ��2��a�0>Vf�Ak{�Ů�٬3�y�EE�h[SQ��Nv=�%�QX�)c���>�$Y�a��M#���y���{9��c�/ � �\�crQW����E��Cj�_]� 6s��o��l���9��������GT�3�`ook�Jf��G��,O��r�:�X�l���.nl����4eÝ}�RB�B��x&���H��?-�$�azO��K������|�<�â�j$c�ԗU%�Q
G̱�ɔ���J^����ܰ����T,bfx�b/���W�Yhor��L#D
^����c^%�\2�<$nj��p�s�P��H�*PJBI����5��\1=������)���z\N�?� �.����;�p�q�I蚔����!�K`¾��/�1AHR�cwDk.�#t�x\��Y�=���dB'D��.0�����!t0vp�]\��猘dO���Ȁ<�'�Xl��� Zҥ#Ü�v^q�3���g�G��Qp>]��ED�D�	�%�F�:"�C/�>(��ciP0¨.��v���+M������nP{���ᄅ�œa�J������1�����Veb���-&\T�M*�m[�ŝc�i>|�K�w-�q�f��ň&��i���*Kf� �!_1@n'rLF]��}��E3aJ��@bb���D-z�GɊ�8�8[�y����%�����Iu쯲����s�[l���2m5��n	��{�4��ƣ� |b�S�^�:?ݺ��v�:��U�O=�0�?���
�T�'Jy⺖���_���g������aO�_|F!'bl��G�2-����;(D!(���_���B�w���s׌�*���@cϺq4�?,��l3z�J�~	��~���� K���>��p �y��	�0?�M��1��>G��y`Fh,%Ջ�jȺH�����D��z�ʘ]�t��9�-��]l�nVt^��0���~���)<,X�U��>�g��Aa4����oº�I���e�W���y�_×A:![��-�<ÿ�[�%b�r����su<���n�5�a���^fL�W�\n�5��������\���ڲ]cY��������$�Gz'��#�6�HpYלI��+y՝s�s�٣^kZ�l#A�.2���v�q���iT�u{*π����R' �'^zE	�{����:WR�k�7�"��Ŧ�T���X	5�ʧim�2��f�%��\��A �g�?��̟�!�E��1Á)���C�4�� �VA8�c~c&�=�v3��HVOQU�����Lj9�q��A��}���+p�h+�Q:2���勬��ɼb�����J�`DVv�ȯ�o|�*df1�n�:��5.��>;�y�B(i�^%����/A
\��f���9�0�w�7i�`e��ȴ��v�0�]��w)_"����4�^%�:���X��A�ǽE�E�����;���[���T�N�" ��fN/�-Kﬦ�j����&Eɯ�w�ef@��V�:��������fG
�
3 ;��S�~.s`��O�e��)� j$��l����9}�%U����>�Ȕ<�!����BT�n: �/R7B� oos1�c�Q�$�2/�'y�
��//jZ�n 0�Y�s���|.B/矾�lђ*�+
�B�ι�Z���� iji����;��Ly��>�A�.n���>���{bOWv����N�Kc�s�J�4���]�?�WY��p�Z�:S���nm����d@,�tZ�'XY�_ͥ��,�9�i�}�*���6���V�>����^s'��⹂'�}�	��ʻ�W� �I�)�� �Ϝ�^K����.�Ͳ>�M��w?�&.�[j�B&�5�:��Qئ�ȭ��I�lj۔?�{��.)h{mY�C��T���>�m�sû�����+x��u�,C� ɡ�Kt�l�N���n�o�J-���YA�~g�	ͦ�]N����B���"����nr����ê?Q���>ݑ���ʴ��^��&�mv�y�����������D���ۥč�bjY���I�h�;��\���!K�%��/���rKB�	��pt�+CN%��������s�V��r� p}�P�$ah�m��	R�&��4l�*x��;��?�`󭃖 ��s�	�:�����p^~, �T8�/��cJ�y3¯��A�.	o%'¢ ���1Ң��4�@�p@�Ŷs:9��`
:N!��m������q�ގ/u.�U��t���%b p������
� }��>�!�~�a��$����� (��4rj@�ZE���Q|z9����5%S)&
V�`�0���M8�—�S��KZ}���&�{�U����S������Eu�����	��Z����.\/���1�X��=������7�~a�`oq(i1��J�]������*����iyq�w�����88���[&,U'��?,;d���(�v�_D�j��4xX��j����!��#�SU\@�(@LW�OV��-��sV�)���amls�䳙�����r�/"Ǣ��l��NvQ��}�xNy��!iI{M�{yH�@���jBz��R+��J���O�H �̧\��=����s��8��A����1ܚW)�JQ��d�� �Ll	8��R�z����~)�ZY��U	�������z|<�$�@)�W�\�s��)?B�;P)��l;Y�p�w�Ha�+dg��]xU���WC������V���=S���U�݁�l��D��6X�J����#8�������C�1����+ަ�T��L��!�e�%7���$k��z�n�}^g5B��5�8ۓ��M�8I1��<~���ٞ�3H����Ee4ү�����w�!Su��-�tmd�cd���>AX��)�x�0����.q L�Ƥ�[Aڜ��*�-I��;m�aϩj.���0��������#X��%_���vX�Y��N�z�4c�=SА�o���P�Mw!T) ���ڵ��$$|�t���b�C0�쁘U?{&���s�~��2iA�9��O�M���pc��t��A��wo���Ul�,I�Fn��o����44������LyĦ�5��k1�C%�A����;#�0����w��>��MgP_�i���S0^�*�YJ�ZY�g�N2�$�z�!��cUl/��ABݟ߷|uc4���ٵ� R̜ O�,�q_~SY��:�Z(	~,���3� ��D��2�Wr�1�qf�>R�zi"X���e�#�`�o@�����7�)�s��� ?Qu�����&l5yL��3�$�LxI|³4fѠo�p���uv��gG@5`��Z?�t�98�M�ƪ2!zk�%��_�����~�zW����V�G��rO�����iI�^Ր�~�v���A�Ѯ�>I��H,p�w���,���;�g{��%�_�.��:[���FV�'���J�ܕ���J�Hwkk�Y�^�Ԅ9���e�S�p�����g�S=6Wy�#@��$���ͻ��Ѻj���0��e\��IyU�vz���;sxY�=H��n���y�����s5���~���"�����B���V��B���&t���gb�����+���@$<�'�&Ќǳaz����y��{�=s��d�w�*�ε���yI��%�)jW�vdw�z�j�~�����K+��!)g����W ��?3q9=ȐMX=�ut��]����C�tۅѷ�,�杺�La�Ǉ��O���rPY���j��xFs�ӳ���	4�N�2b)���"w��=�HSL�M���%݅��M=��Gyz�ĩ�3R�X��\��-ۓ�Ō����d�ȫ�q�):<B�7碑����e)��۝;q�4�˅��wE��4�[�1�ƪ�mp�r�TA`NIH+�T������p\�,ٳ��^Zs3 6�*-��N�-�Gb�i*��#s���)�w�W�O)��@8�㧜�~�,��5�ũ2M ��C�k�@�a�3�E������>�9�_���z��v�|&ܹ3[�8/��k�&)xlQ�/=i�J���H���T��n%�G	;����᭯ .|5����
%��MrZp�����}+��#���� 78�LB�V��V�Z� $��j�ٚ����Ǟ���m�Q,���O��'{i���>�
"�'Wl?��/Z*䠲���no�I:������aV$�乍�a׶O��	�^2a�V_��b?��Gŋ�����b��A.e�R~���>7Lݠ�5���d[�7Y�m|���O5E��_
�)M�A�=����`ES�����`6�i�V�M֦C��c��/�f�v[�⧼M}����w�a���=/s�����*ɀ=>-�R�~�-�O[�D�;�d�b l�r�+a$�n>-Ҍ��x��/��	�B,�yY�"EJBeY�Ctu����ss���_B4M|Ւپ��8������{�`�t":���qe)~B~Ѡ�:�"�1@�E8>��% ϗ��se#���O����s�ZA�B��\���v�r�&��VCR�Gz� ����&kx}N���&�q̵�1���!�J��)�Ϟ1-��[�T�К�Gjs��~�0���|�4��g§���D�"�R�2�(�ӌɒA�����. �EV	��Z�K��T�Bix���2q[i�p"N�^�U�Љf�y�����9'�g�&L,���Y
��ȦTn�NUꛫ��*v�[ԪiܖTټh��dd4��7MO3�;���Ê���Ʉ�hB�Wѹ9�^P�\}��~m����V�o]i�&H4
٥G~��,3��O�ų��Q�8�ğS$�+���ң��cq��s>�u�[R�=3�n��q|�#& �9~�M�e�/Z�	S����8 j�}����fk�|�[�V}F��|�hV�E�-�!E��VJ=ȟ�T�^��ߊ�^4��vE�F��z�����B��Xp3Ë){F� �:5l�Kb���i5�������gg�S�� �g6d�"���<L� ��`x��,��&�K��'N0,͏��F��	�w���w'�LC7-`���y��D!;<52�Q1s\�+C�t%�?���P�\��JK���t~�S`��R�$��S�4J� ���J�������뱿�G��x���H�͠��#M�\�|���2��PSU�b��*��9+8�r���Ȩ�-�ʏA�	1�ŽM�aKF��P����{��ii��`B��K�Vz�;}-��aO�n�j&Ae�!?�;!g�5H�!���vN}:\'��5{$ok{�HZ7�$����w�T�����5���ܿ��zșRR��Ȭsc���2;P݇`������m���rP���L�w�|��\�t���#t0���tK�yœ?o([W��6 ��=r�m| �,+�����N�c�{\�]Nvƃ�<s#�7��Z'#4Z�(�����|��}� nC��y}��[u#	��[
a����F��N`��K�vZa�[_�^Ɇ�<�:j]�q��W�_��zoM�:bY�R�'q9���*�kUn<�!Aj�����l4�#k�h�s��; 1�ǔ<u['��("�X����D�
� =�m.G�]- �r�E������\_�F������4�ﶡ�Qpw��� }c�����"�OX\P��=�K����cM���.,�%J@��K��>�q2�À��^����W"�@���IŠ)!� ���Hc�f���"խ�I-D��7[Τ�9"��~G�� �
+@w�j�
����=��K�!Vi�/��o�U�]��q
�i��-R�����[B�Pc��tg$�6e��v���cF2��Ux�+x��!���?_�W0�bb��.Vۻ�pȈ�b��<�	�Z�(3�j��%�܄�����+b6Ȁ
���˘�k]�cԽ�`�<T\^�x2��e�;�j�z�r�i�����E &�	�PU���������5�mނO�9'�~-�b��~�G}�p�'�.\,kc��o�0\�����f]�We�jf'��Ȝ	�4��t�|�~E��f#Yzc�j&��+�V�`����%�L���n.Y^- K���H��(���9j�1���yX��fz�P���9�����ghR�)48D���-�%��� o�-504�D(75:�Yf�P�μ�JQ�����UQH�9�,�3"b��e�AF?Z���e���R݀
�Z,��#�*h@l#���Ojܧ5�>��{ŵ�vv�*����ӉP79�g�Ǒ��{�
��"~ɱ�]>�+�Y�C��=^l%��_.��*�g�^gq�_a��ʡJT���Z��55G�<=W��pp2:��RG���[(��샞����f�8�On���Q2F��&7�'��3YS1q�k�IR�L��U���I~@K����.0[q�)ӊ%�I���o��}�FM{�Hk�gZ�E�U�W��\�?+��l����7�\³��f�f<��^��V�{]t�t7I��3�pn�KtfZu��?V���s�,�vF͏�Y����$���L6�*-�/�Q;f��c���(]: f0�����x����.X�&��0-���2�Q �
ث�����i���͎KT�nϤ�4�s}˗g2�~iS�Ŭ�F�|�!�)U��p}?�D����r��UU��<a؎��
&�:\�� -r�ؚ� C���xNd�-P.��?mp�N�6�ę�����K����BN���2%��b�c�?�PZ�#{]Ku�
��w���}m�`������s�`!�\�����C���ɀ/ S���	�\�O��bL2ע�	+�u"�Q����p�#̋��WOz�)�l�pw%�q_up��ă�h�N�h�MH�t5�{0Ɠ�g�O�i$>,�KP%��ʒMnZJ��/e$��Ը]��W����"�GBP��
�$c����7�4|2B>���#_��� �~9�i���"������-�!y����{��J�?�zQ�e ��drYW�r����zE��:LYz�w}ᘭK���J���Z�(�!��REhY��+�ڝ��#��ߎ����F��s~!�����ۦ����D����]�����i�U���E�R����{��$��@l�u:�x��0�S%�n�ɘ!�(�6iBN����PFB��ʧ7B�FX�F���*3���Ћ3�I�Z�ٲ:k��a&�H��H�7�xk)��9�PCJ���^%K-���,�d�����#�K�2��oݒ�X�HWM^�v�^DU�Ǚ���}v�O/��JK��&TE���|�,�EӸ�AHCZ(�C�O걞����|]�E�#𙺟�uQx�±`���߳/��0�J��E����p1�i��4["��L�����!`d���l얠����"�c/�j��R}Ds���1B��w����}�#f�B`Rj���o������wlޞ���t�gٹQa��#���l>
�)A9���y�"c�s2�ЀTt� �G2��uU}6��=�2�ww���o/F�P\�fiY9�O+g�o62�ǟ���6�򲣀���;y����"(��2�.yG����$҉�r�m�o<��ֽ��U���'��Ԧg����r�c��zw_B�������z���8[��,�.	E�1(��k�7`��XS�d��M `J�*��r�{Uq�����Q߈SMU����Fu���%��
�CʏN:i���H��(�b��n��,�5���~�Sz��=i�=���,��si#�i�5�P�T�6�'E��g����)�:�,�s�!��ۋǩ�G����m�� ���.	������ ��� ��,���h�G	�Nz��fvC>a��������}?�w��Z��g:�`�X#s7��h@Tn�(���@��'DFB�8�ܚ�D^B�JZ`G��Î3̒����@4b�g�ۋ�� �F��\�O��1:�Z��P�TE~�H���a���*���|@��pq���,ÎPg�v$O��B2+���pP��I�j[�nv�Z����H��jY�I�޶�8;5!{L�m�fs��q�:���}s���i�R@�<?`@�c �X�\d*�m�c��i���=�&�����0YĶ�l�?˯J�Kk(���H�,���6�j����d�3bL��@�G�:�z�P�v���{�əb.h���"�w+��#�\%�b��h��~;�r�v���k�$Ř�m7T���� �y�C�x�������ź�EK7���$��73��4#�����T�j،	��]�W��c.�ܷ\b�^Q]0i?h�Q	��9��+�R�t��n�3�L�ˍ`	��=a�U$!]L-EZ��t�d�2�-Ȗs�P퉟�H�p
ڂ���+e�f����yT{�@"���7.�S�L��>L��-G2F��Wm�2&\�{(��!4zC��~�d���2�f��gj� 4�k�+�G��Z�S,�!�B�;���c���Z����y6/7UN�B^�E�W���'?!�%#�Cw��DT�p�y�� �#X�gV��0�r��I�ެ��[pEb�y���8�����c9�4v���_26��6��魅����`
�&��0^���V[�������f�Zj�&��<uj:ٲ�t>.��eD�b����#l��|��McW�G2��q3+-8C�?�g��i��|�FT�ͪ.ogb��|����v8�;��Ek��;��B��Ҩs��iF�kS�z����6�7�C`�9Ri6�<��ǒ�k�|0��5�)����S�"��gE��7tp!M��t֓�0�����e~��FE��3��1�J>�R�{\E��&��U��i/��u3'���K]�(G7�M�gס��0�b�������#0��n�DU�?�D41�3�����:���_\ ܲ��ɸ���@Zi�<)�f�1�c�7��mm��������u�-^6@4U!����E��x ��v� �A�?u���{�ǩC|�c�$��ށ(3`�@��bh>���@�<�6:���<	���S�FA����C�<�yVy�E�9@&�Vn���ù���?������s,�D�p��#�K+�9�׭�o���5�Vn��ߤ���Z-�$��(%2wz�V�c��ܪ9a�_&n��Ǽ7�o1��=:�F�T^��Bt�i����0f$��j��Ow�	J�����g�Ґ�N7����P��*ǆ�N͸U!��wT��ᾅ�F!�Re��N0U�	�t"���vUx������^0�?�,��(��.̲�2�d>�&9�jf�ױ�O�!�2��`W��D�35��>~�f�Zk�&g�]�Y9~_ōI��p ��Cv����e��j~�7!�G�wW[�
�k]���<�K��B��_���ٹ ʎ��
����s��d�%�O	��? �C������j ���?m@d&dޑ[6�r�Kh�����Du�����!Qw�_�c�qZA�Hu�P��]\y����7�� �7� n�j�D9�ņ��#�k
c��}f��[8���!%��_�{��z�M@-����@:�_yv�}W4%�7yic;������d_ѵ�B��H��cuc"�g��)<>32 �������]��zY�S(���b�s�v����oߍ6>#��L�?��w�fT�mD�]�]�Z��mu&����{����̾|���@�
k&�Bل���Un�/ٶ��m��� F _u�s�Lڟw��s�CQBL��Y�����g;! v�,tw��2��H��6A�ʟ�5���>2&����@�j(!��h�p}�T�,�]�[�i��&ŀ��R3�A6Б	�z���"e��\P�2�T�A��7�v�X����o�K�-��`BCR�	*:�32-� ~�0��J�ݗ�ԴY�(�8�5@���'�:�FT���멡.�v1��Է�� �N��/J/8�:�T�F�6������
�ր`�-����=F9�'�ǎ� p1;�	�d��-������,\z6[�C���#�
���s�K��jS�,��6�6�����(o��/��5��I�t )��+m�aC�1��e�֮e��V���E�
�.F}� ��������0��C��a��4�x�B�(��P@p�;�v5���	�t+�
:ְh!�ܨ����0�&���1�3�	oOKk^v�M�J�".���QV �=�P>��}�_�(�%��6L����È�i'� M�wCNIA�V!��vd�g=�{6��!:�HsF�	:��D�dT��C6�*������L-A�f�oI����r+�X�#����$��bI��pL�iB�|��|�t(����D��-�'Io��TwZ�yIW$@�b�	n����/�2�:t2�����!9�J�T�װ9Σ��/�v�@�A�Ϊ�ET}�R���x4@�K'��Q)������h� u��"#�r� �LsV����Q�4a���5�]��V	}�aˑR������8K�7��c�2)��51��?63�$7�6K��.���R�v+&�'�v���B-i�����a'�8j�G��������I6y��o�	��c�i]}��0/��x6��0, q����Dc=A$�
�$a��ćߛ9Z\�&>�V��~�D,|����ߝM%)�`Q<L3�e�e�|���x���˩K�#�.(�p�U`�����<�4�[���ЙJ�j�Y�`�,��]�� ����dsUQ\�޽'�Tz{�p�Q,�Sa�X�7f,���{K�M�a����ƹ�	�_Ԕ��a�]xD9�r�ۅb?�#��ɑ^�b]8�*Q?�Frqb���(ܓ�1�E��}|/��M,H,�#�XL} B�&͙�]V�^ex|&��=���K{.��b#by7���l$�)���?j�]~��*�l�3�0�o��.~3�>�@��IE[�~���T��ꚤO�-�����x�M󦨥C�#�'q��/έeL*t�+��	�ؽ���<[_KR�̛ç����u���*��B_��>c�Aηj},������Κ�����+�/��u9�A�>���+�xc</����}�Z��.��?���Ǫ���O���[�i��h��EJ���yn���7����f��:�y����۶�p�w	��V�j��`I��pk�|R�
�OOa&�ǡ�Z�� �l��H�W��wm��C�ـ�aeE���y&��-!�YI�ZuG0߾���\{&�V�>O����:pހ{��~���n��Z�3�w��ԋ�`�c�a&�XCc.P��4#�3g��+AsNͭ��8�M��}�0K��P�R+�a��; ���A�SRQs.<�ڕg��UZa�j��Y�WL�e�������O -���RzM9�U�"P��4�<mE�����ღǸib���ׇR�ö�YӼap��$l�]D"��ΘY|ϱ��g�$ppU�N�T�(g�p:~8^�>�6��l rq��	�r����ׯ�_�K���U �뵴�|�D�Oİ.���	�i�RA�8�m�Յ������q�p�U� ��^X,j�A}��쐘~��_����t�p�J�=`�0��M9~�Vo�R����]���j�7�R��:����Ql�)D2���ɪ4a���뿳uo哼���/������2�����c�.D�q!�����,&���A_�f$��S���/rG�E�U[��/�f]�pɲX6c�'7)p��٧�3��*�b�ޝ0����r:�&i���`QJg�f�]�ja������i*��ߠgO�q�mS�bp���)tu�2:��M�;�lwa�wC��UirY�Fk��Œ�K�ncC������9��h���s���P�>.����=��j"��Af�\N.�+�d��*�:�߈&�/t}�_赩��7����&T~F͈I��l�p�;���i�Bo�bgRc��ȥLC�����b��\��Tr� �9
���+�=�5�hΩV��j��?���xhb�t�i9,#���[$���	�V��P��g;�n6_W(0Z�X�@>W׫>�+61~o�#X�tר<����\�q/&���OYdRs���M�M[���oE������vu���	��uUm9
�������>�e�U��euN�U���!�U8fS�$�]��S*�$���.d�n4�0��_�H����
���H��hf,7d����t��1L[�V�Ƹ�*���=J���$L۾�IP'�^��4�R��p��ܬ0�J$�����@�1����b�(]�%F�0���,|�EM��_&�)p�k��+
��"�'���

��ʭ��V��.i1,V",;��5�' E� m�jϰg��/�[��aKq�헣��� �F�i{
E!{�U{�êY���<.�����x�+��E�\4"8:��z{l�e@�o�"��i��F��1��)n7<=�F�dH�3hf��t1��KM�Pbi��3��HN~Q~�Wv9���'� �u�4M�Gp�w�V�U|�`>TU���[�f?��"ou>�^�������A���W3�/�)�޶=F�\���J�]M�t�)]��9f=�>�y�8��n�E�z��Tm𵪵�{C���t�>�ڃ6K�ċ/�鸗|��=l7�clp���l"���4\Q�m͚�%-ol��M*,{G���g�L���p�]�p��1��J��>6LX+�9ҹ1I�\�4J,%Q�����|G��X��89�A����)�w�*�3o�~�����]B.�z��D�c��?F"�#��4z���s���/��F�~�'��;��j��r�}��D�ʑK�(�,����;��X@�=�+�����9P[]�q��d^(M��T��O�p_��=�؅�1��xA|���t֞M�����t���:�vDg�[j����m�i|T(b��g Ji �,@�Z����FpmM���m�/����ɡ�P&v<����'�<��?��)��|����?��@�*�$g��V����vsr0=��"��[���HrČa,w�s���I��PL	��<W��0�.���n���j�P�/Q�E\@D��s�8��G�*�#�n̔�����&�2oJg®%�-�0�ͺ��m�9р���B���^P�� ����8�vl���h[%΃�{l�Ȧ�w�怆��:�It���v�
#�PNL%���N���w&=��}H��Jp�G��q֨}O0b%��Ӕ"�3�{ T�R^]�\^�)Z	}�_>�B�u�{�6;������F�$!�U��M6|M�&��g�l�-��&zD��B�2�k��_M����G����X�B�)�1���dt�"f]�@��3�/�UV��E3"ǻ�%���_H#�/�Stص.ۛv/�-K�z��&.��V�w���l�i\Jaӏ�#�;[��I��!e�Z7qc��Kp��,��<t?Y�q�J���mI�R�@�Ƀ띮+:[�EzL2i�7�^�a��7�ȍ��XrEV�O�W1\˴�*Y��K�v<���o�?p��u˹8̔��| �X=���s8����~4'�:�Q��4�|�)L�7��'�a#p������M.�c�묇��VUA���<��+�ONd����i.�� is\Z��}�V�r�sE�_�d"�sw��NF�D�YK�:š���W@v,~��+ݗ��"E��@�l
��q@�U�3���R0�W#�a	R�B����驉4�!KI���Y<E���엝XRʙO��A���^)�R�ͻl]�<��>XJAVG����e&v賘�{'}(I%b���	��C�x�8�!‏���7i�
�˄�\��~EqV?6�@����Ֆ��
���R��E��h��Z*6٩O��;���*��d����zᡒT*��O����-W/?�Ŋfd�ߺ����e~�|���kqasG�ÆAa�9M�_��BF�<'�uĐ��N��n�����z~^���>]�z��Pߦ�7h�<����%98l�cΜ
�>b)M�tO���q����/�V1F57��K@I$!����M'���)|@�ҭ ��*Iٕ=o#%�:��U����[��� ���F�'t9��]�aq�Dpd�N��V9o��[P�i�`8����IR�Ljߨã�i�.eSA`��q՚ O��eR�� ��3�z��@Q�E���{
��p�[�U+�_9M��t��X�.��*���;�'Č�c�౓���J����m���b6�9�1��B.�F"�g��qk5�5��T��l�i�Z�ًU�
�c�)A�;�TW�2�FN`�~BC(/\+h�������������k4T�ʎ�z�� �~�Q'�\���.�yƍM��>G�_��_��@R���5�!���|խZ�a�W-U5���eBzդV����Za߫&����E?���c(OT���
�~4 ��|���Ή�����K>_a�
�֛�3kp�h6��V�ch�S�JO�[T�̨{Ppҕ[]���7��Y3�+�_CD��@��uW�/�P^�}&|���&�&'':C/���R�m�n�aL9:��޷�=�[խMC�JЍɎ*L~H}IZ��,�&�U����Z�Xյ$���j��0v��j�n}\O���t��[���B_�G���A�Vb��J�1~�KT9n���ݎ�*D�3t]Ѷ�Z#,�e�>P�8���������>n�����rD�쎥��@��$+�P�>�Wؘ�)hW:(�j�Ėk^���Y�d��t+|���n�y!�~kklP+Ӽ�m���'G� ]h �c���2����լV-�3�j
�n��&�@�r'qG��~i���Ȍ���xW��5�خ�
���з�C�ө�Jd��~�c�%�ƻ�5����/Fu�Nl����Y�<I�%jR�6�X�(z��� �|�K�"��|��
��ґ��ʽ��l@Ud˦u������x�2����w��(#z��J�})�'��ƠZID������w&KG���u �７�BI�{l�؝����Av/���>d�¼l��}0K&b�˞P��NQ%��_8]ȣ�G���elB٧�xf��
/.Ee;Z�A�j�D�b�z�)�@�Kn�)�H����uZ���U '�`��:��K��.㿻�됎�����u�?�`���.XM����s��Y���\�D�~hCA_r��nvO�`�c4~%��P6��5��S������%��y'YL -e���kM�m!4���~X᠝�;~��c�2k5�����MtB]���`��y�w�y�gV'���܉�WS�9���a�θT��i�����
f��^���:y��Q��`	mDM>�⠬L�.<]�,C`�����
U�F}K�d��Od砈)_3)� ����$9fIq��Ru���W��!;bg�B4���/��D��g����AK ��Ѥ��R#k���������ρ�CBE��\ ��r��hb���9,t��tx�.(Kږ��Ʀ��x��o��z��^�ja��0-�xB�%�����hC���B�s��DL�Y9���&E�%�.�~K@��j��H�Iv����!ń���hQ�te������(��$#Zh���K�Ct����[vC��N�W���K`�����Gȸ�<*׻.��d��r�랡S��B&L������H�$�(q]��C_���pAH@�m6�IuQxI�/>HZ3�����	06ߨ�3�wt.�y�9%�Ði�R�
�O	�7��i�8�j����;IL��."����g�JE!J+t���`+o7�&�b7hfH$y)�k���B铣.e�Dq�ė<l������\�+�c�=s���Z�Mk�*��̗S�bh��ņp�0�m_����ɩ"�� ���5����u���PVf:(��2��?���|��Ɖ�t�x�5�p�ۭ�q@J{ܞ���8Q�U�6�c�EI��%h��(��4c��E�r;�;7�hR��J�mul����q�9A���W��`�U���\>;J>kV�jݘ�R�Z�N�ex�_����z�K3��eJ�b.sT���q��5!�!u��L?�Z��_|@���\�Tǌ�î�;ۇ��r񧉨+�(v5�Y9�ɽ��%}!�x�3�3����J��&P�{��EwG�=|+'E��fQ'�^8�n�\Co���lJ���q��W�յ��\[ӷ