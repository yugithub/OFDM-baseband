��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6��a���$Bh�����hul�^B��9���&" �Lyy�����Z;���k�~�ʧ�d��Ūt�� \&���Ų�6�t�ۿ?^Z�|n�M{�EU�Fbrq
M���s�:��\�S^����ހ5OT�/ק~ez�T Rºե�L����	�^j.�TRe�y&T���?�ҀJ��ޔ×3����
sJ.� &)(f<U��*b�+�*���C�#�.u$�@G6��ݳx�e��`��b
����P��.+3�go' ������o �U�����1!�P!
WggF���y{d����/v��5��t)���n�
���wR���rG{�
�.��t�>�݇���c2
�Q�#�`��A~��`lJ�u�)�zQ�;�/�-L�:�&n乞��x
���V���6O���`���n#3��<��<"�B��H~�,��o�5���	[��td��ӅpD3	Ʌ2��.����陚T�@|����'�S���}H����g�g>5�,Q���mL>z�`���n�h�5a�j́��g�`�*b���Ȯ"��֝ɽ�r�'ޞ�gȰ�
�0aT���K�7��B�S�q&nԌ���>��q���ZvQQ��$z���*��q-0�L���"/^a|��@����B�L价\��Z؜@�8��֭|����%Uk��J�ѷ�FFZ���)�~��^��F��m!C=�^�	�%���h �<d�+(�'�#�}5�8	��y^�aC��Waݱ���+���a�H�P�%�75��O�mʎ�tX���'�9���T�+_ �oq�%Q4��9�C��eb+:R^o�̾=@0�A#�02�:�d
��!�Nos�2�M���}��눎ύ_UIA�H v^uy�xvi��R��U��;i��Y��/�m�}�+����w��+�W�`��^�YO�~z��w�!X	%�*��v��(:��ɭl$�S�!VM���>��wR��Z�K�jTX��D��a�u5�!��[�C.��:F~S@m���\.��wa�gI����#��z�+�W4:��Z�^6�[<�H�"�6Ʋ�毘�uiU�^��|��f̅��B�>�=)Bo�dZl�5���(y�(e�x��W��9�^X��D}"@�#�ho����Zd@
�$�נ6���-����@�H&궮�4�9��3�S��Y�]��?���6t���n��u��1=�x�N�θ��.�9���^i�����'?�[�=0Q݌P;J�M.��Ɲ̰N�Ґ(�5�i44zN��} b�:�I`����a4��4���O7�#���6<���c�%��؛9�Y�������.���=�00��e��ڈ;�o�E��@&��ĺa�tzPkL�=Ku	��ӠA���F�W�:�(���ک�q�O�	�l/0��e��/�c8�!��������Ća�_I�J��2#\:{��O�to�{B�����.p0;9DDU�`�ԯ��d�FJOK�ܖ��O�B�Df�7>���iM���Օ���ӿ�)%��{��$H��xۚ��!b킓�*K�9�aI��){ަ���Q�]9Җ_כ��q�={�(Qqw��M�О^�B��z�f=��nz��>
�;���m$\�l�ql��*;M���J�ǣtx�e._F���]�t/�R+z3��G~�����x�H�d9KDg�q5�ʰ���t�%�&�H�Jm 2������|lS7�pW}���V6�4|5~�ȩ�Q�q�,o��9T{�?׊�)��ͧ���J��Xdgij1\�+km����n�ٔ�����o�܃�'xO_�x#�LԬc�H�opH�zq�|U�d^H7�m��ʢW�sxہ�>˗��.G�@l�
����׮Σ�1��Z���	㧑��H�F��w��2(#�����y�#)O=V4|���9����g��K<�nM���OẆ�!\:�17�@h	�q^i�f%uo��������3�q�6B�3�X�КV�?�	�|b��H*N�fi�J�=��������l����3���$��`�9߳c�ԛE���
Ad�6�_rF?��e�%nʃ>Po�\ܣ��e���B�?1.b�S�,��V�hn�ocQcgj�
�xS@��7�,���q3�0�g,RP��?�hd�`���WHk�L׎3��r'{�PV��Ǧ+��'Jf��Y0�ͳ����X�q\��㽄��:�����	г��x?���!u/x(��;\�:c��Ҳ�+����5�;�L�xȍ%
���n����nl�*�n�A��D{���o���
	6� 
��Π�Zʕ,�foϪ�s�8�k�͍7���w{~����-q!|�(:s�+�J��B�&%j��K��0G�W �l�Z����#h��^I15b�D�+���������U�d�A:BA�y]v;]u��b�Ù)IN(qu����KG>C���f�F��[m�Xw�=����.�7d��5yo�����	W��";l	����aUø�+�\����n���@��{?��%GV��;�3Z����{��g|R0	���'-	{�wQԣ�8�|�Щ\�E����K�\�(61|�,W��-u�J4~�d���ك:��-������9Y:��Rp0�m���W?�Vl�}�����q�}wm�fN���t��Ic=9m���Q!��nH�J�	臰�C�&>դ=�f���h�؈~�t��G�m�;u`�� 0�S�*(��f����s�<̘)=�	�Fa���׆�Qթ�΃�	UGV�:Ioo
�Wv�w�x9|v z2y�i/SoU V�@��v$	�'�b}-��4L1��V�QvwY�V��)qN���G˧m�0��� ��T L��ic�TIS��#�f��j����9.ڻ)������e��#����b=���J!%��m�w�X��fܧ��W�]N�S�툓���Ƹ"ls؁yb'���]:��ŚU\�~��pL��U��^�l����zuL���s�^*n\
���&/J1�,�j7���Dlf�k��FBz��Bϔ�JB0Þ4}���mhss�;b&�k9�Lb��7�J8(3x���
e�F/�5<ޒ��Qk�J%�T6>F�a�YS��dJ��5�Z6_�QO!e�L��/��S�N#S��{�,�_�m>4_|!2]�D�'��!�pXu_/t`B���-+-�ؘ)�K%�?>�TU��K�pJ1.1|;�U�>m*(�G�6��D'���H��M���t�	e�˔i�&�^U}�ϩ4�Z#WR�H���x��e��#�� �{��Yay^|�&�S�km��^W!�WvPo�L�����n4�DNOK֎iO�$~O0��)�5�#)������c��� �}F� � `��dՁ�S���>7��'���|��nGԝ��Lu|
����o�/��Q����h��:@z�y9��Q����lRu2h�Z|���Igz`˻�pj�U�Ţ~��t�\�ظD#�w��m�
a���Bl�h�=��x]?ׄj�V:�����B��j�y�~d��a,�2O�f=�ulk}@�����(t/wc	����o������ُ�`���A+�`��@�V�?x}>�x3UXC��7ߥS�������KWL�N�"/�ɖ:����UV�����XѫҲ��6�j�h�ۃ���[��#�Y�:u�)T�m�$O����l:+AM�DW�r/�����̱����@��7J����2A͵V�˥�w�*[G���`�9w4*�@���Ԁ�n� �{��p>F�nx�vMhQM��NT��`@__W�?
=u�$V`N԰�5G3��:_�H8���NuD�)�>����-�_چ�����k������<�c�9�$�b��63�/��]�M�$K�����&�y�_͂�U��Ŷ��}b�%�#�������7#������Y�.!Rp��Ԍ;[��Ӛ㗧L���iɎ0G�3L��ؓ��uP�.1�)�-qCm2:t0[(�.�`�WW�ġ�+h�&�*;{�m�MȠ�*�#���v�#���[���5�S�/��f0���OW_,���"��l)+@.'���CZ�L:��4H�H�½�OD�&�]�DV�Q(�ŝ�k$_�S)�u �o�Seix�vrk���wxԈR�����^����CM�1�O�V�]�k j ���}]�����8�"�d��XyC�\���0��ӊ4,��8^��F��"�8�|T�O����1{��@b�l��H��L��e4���EDsgj�&W��o"��_�p�h�/d�8�R���{�	��jL�)�l=ԫV׸)��'eq�����HV�i�ז��M�	�*���y���w��3��Xs��3��c���J�#+�r�⊵�"��<���������7f�ue��C�;���3G⣦%e� 
�AAtA����2��]��x�j��I����hK:�/��_��'���Gf�0��O=Q ���T���9��њ%�߷���{�(S0.Seⅷ���T�����p�`��n�Ү�)����,w>�Ι
��R��a@drdv&�Lm#N��a��Uި�3�w�'bF�G��������պ/H��@v �e�>_�����W�K��!�q���3ep���i��F�}�}�_p�\��I�x_�A�;�i�T�vR��յ۟�b���u]q`:"�1��I�<���>l"+�,"�ẓ�I������|�]�d�?H�-8�ڎ[G� �c���.�7&ݑ_eް�������zڧ����+��J����u�p8&���&ڕI�.���V���������ZR�Bޥ2�D`a���-"t��eY#�Z}��`���>Q6M��#�ǲnO�(yT�?��iT�i�`L�+&�@������!jV�tpQr�EȊ�z�*�Ģ�=�p��(O�^�J�!��G5����o���T�@�H�j�^�˰��=��+k�Ё���Zo{���4�������.�'>��5~v����Ùr4y��ߩK�l��X$΍9r�ʲ����[����$��П�yx�g��(_�Γ�Ѧ��K�~��F��G7�^AN�Mӈk���P�a'a��$�<!ɗj�
�
��eպ��e��0��&&ǩ��S�2M���û�ュ�"gDupp
��{��W��ㆶ�.�"���s�Ϋ�N������4j�\b#�g�*%���=f��۬�����@�Q3U��/[�(Ҏ�#_ԡ�kp����!U�o��^�w��`�ky6�,@�k�A����a�W-n-���e����RBHi}�Qj�8要j���H�?��A�.$G�
��6�%X@�w�~>�f�0��3�EL�6V[n��N)�-��P�Y�*hAW�mզ�r_�z5�e:��P�؟h�}���h�D��'�N�7s:�`|(�����aUg�dX�
K?.>���ǲi�������h�&�`+	
��!�U��xܞo� �R�7�G�T7�R{gI���D}�VO!�7f`����WB� �M�m/�
�U�%g��pف	;H��KnK�u#G���G4Ul/ʇ����wys)�D��[��l������J�b�%��N��P^*�G�����ړ�U���RI?N�*�ka�#�F�9������K��V#�.2:�,K���IF:���L�O�!��ʗ�n p�g��̢�y�xgz���z��`�o��T�TÛ\7�yiq��v,���ӡӖ�Lgy�eS�/x�Yv�;D몥�K}�mh�x�S�A�#|��Du�e���un��(-���&���W���]��g-��S�����赩�t����/:�Q��9���]MX������۴�$���O��@X��'[��,ͪ��~����2P�?*K锆�J=t��|�5Е}������Gl윖}���d3�ƫ���P��TD�j�"�_����<ވ��ˮX>��rjQ%���R� �0�Nf�h���&�/x�pF�	KI1"q�}W���l3A'��֡���d�Nm��W����%�g�]��ˤ��,s��/閊DQ
m����B�ȕ^���RylZ�gL���?=:����f��8�oɳ:�uv�1QlO�b9��8�u_Ǌ��wWs��k"w���!4�F�Pޡ��Z�mG�m8��?�6�H�Jөt�$CW`lg������C[�۰$)���?�`�y#�U��g,+���h��:��`��x��}5�ػ��d���ԟ�/�Ӥ�\\���sͨ�
�h���㜚w�����H����Æ�h^�:%��ČL�=�<��Ӏ����k�v��L���$�/]ϊ��C_�Q����	��r�k�,�1���q+�
ui:���Gb�F�)L�?��
a�ƚ�["�Mݻ���*;?���6.���� �/;.�G#6	��h�ӭ�(�5���*���oYL�7�����D
��mL�d:��a*�599��Gd�ҧ:����`�ϥp+�����7�CM����������0	��jM�����y ��W��,3&<�"A���������"��{�������G�j4eKq`Nהd�DN�%jz�K��~����m�͙��[E����9��Z)�л��"�l��!�_&c�Av�S�w>��Q�W����hjb❘8��q�mB~�C����oK�S�j���M��֗�q�)Xl�dG����C��2k�~Z�ݒ�M�̞e4L4�4u�_�nz�Ɩq�W�<�撰87JVD'V�͗��Q���3 Ύ
�C|�R'�N������,\�y����&d&a�f�Kdb�|t�o��4�}��x:���G"����N�0X�8�1�W}Z�	��{�^��7�h��1���@�U��t)�!_��=8���L~�B,�|����9l��%��m뼚�"l�w�6mВ�7R�Ңx?�����]8@]-��p�����?1C�6�~���1эmt|�C�����n�'�w��֏��X�ޝ��#uU�L����P^��@�K��v��&l��7\X���EƮu�O��/�e��'#.�)Z[2n8t���Lgl�oظG~�;�d�#6Ȉ�/�M!�R_L>�j#xz̮@��k����a?�?!z�]'s0���p��p!V􉬌'W�A��i$z��@t�A����.$�5M�0ڕ�y2*�9��*�5�_�������dB��1~����N��b�<��8m������AZ�)��F���Ax#WJI���Y���ۏ�����#T������X�׌�.��C	gH��!�^���e���`a�
�^���H(�r7�]}������]A�k�V��������F�|�N�\��SS^�,�^��t�ab��9�x~�s:`R5����f��6{�WQz[`�}��t^��X��Jfe���C�T��M��_L�CJOG @���T���յ8��&�շ�!D�X�w�w�^�W	W����.J����ٖvk�S��/�u���6j3�]	ۄ9�i�����P�|c��E�%.E^�L��b<b1C�=�~���:�S�j��8�������;��9��(0l����p���3��Z2���<�{�qD�\�w�%���H��Rߟy�M�"�cDՂ��-Lr��׍����N��Q�)��^�&��c&��뉆^�p0��:��[��
�JI�	^�(�\��Շ1�G��cOp_*
�"�V2�i�Z��3bP�!�b/~jR�v˔6j
$�B��*�E�\	p�ⅷu��S@F�w�P�N��n�z�F�������ڊ��9��յ5@w˴�+�r�ͯ�?��ɼ0���g	�uʇ�J��?�%1��Ԁ﯌�C^;qJ8W��\T\�06�����J�j2�Q7Ky�Ħ���Y�ye2���������x�!�����cM�� w
*.� �@�*��t;ґ��V����A�mD]��@���������lח?-LuǍ�MbyQ���;j�Z��(��7"m���=bK*��9�є���Ky�p��A�~z�Hiv�"\�5�	����>ҩ�̒&����1�hvi馕4u�tּ�ߋ�������B1m�NaD"���^���W�H
�ʃpi�I��9D	f��C��Ԥ��+���"����<�k%����0���p�Z�&U��-yJ�|�.fh��R��m\�,�������3C��@Z��30A��P�dj�/����-���2��^��G0Tyl�TY�0����%������K��{��fI(���П�1W����K}�*�����!:ۛ�I�u	�r��=�<7�"�7i�h��Qbp�Vk\�BT�S�/����|r86<�?���^$�>�VT�W�!��F�߼��5TpB��@V,v閛8�BB���3f�_7�ŅG\� �Ia{dәau�Y�Ӂ#�I�"�2(7]�b*���:�$�����g�K�vS����%��u�"'={P'�N���2��ƈ&��2���եiqgF�����q�(̇�W���p����5u-D~�K}3oGp�\�kĢ�ʬ%���.I�aa�l>�Elo���$�}�%�ܒpW��º���ga
�#��{�4a'�C���1��̤�[)i,��`�U2'f\]���^����"L�`��7���H�����U�e��G�g��@5P�r<c� ԁ�i�� �#N�˦�[����=�)����ߝ� ��=J�\/Ig��������(�DNX���HWد����  !628�t"�V6����\�~�d_v��ݚ��3�C�Q8�V"�B\􁢖�������M����7
J��_��mg�Z����Qg�P7�v�_a�d"��
9��7E��)����T�Y�7�К�s�.)��vƊ�P��U���Q!ww#/%�ېWqS鍉�ѐS@Ë<dZ��D9��xVl9cwB�6��kWo��q�y��{h�������Z��t�K�vQM�ɼܙ~��4��B�(��O�8ҷ��8�S�=�?(�-�AT�GYrj�R�Vc�tcۜ��޺φ�H�8�����X6~�� O1�Bݍ�n�<8֬�2�!=�a7T�cI#�iT!������#na��3p<�$1�pV��V&��VxB ƌ�yI0�Y�b��B�*�|1�%������| ��Pāe�9u���~���-����}�3Uѹ�_J�׬U�?��e�%{�w���rG�R�sZ����j`��\�'����<&h�3��7(?8s�A<bG �I�b8�\�mkQ4�ؗA�HGY4.���=;���H�i�����C ��e�
f��0uiJA��m:6pϵ=�d�����e���!GJs�� R�^4fi�V��<����=�{sP"'�[��^��x�<B�;�$�����W�N�F�3��81܏���#օ8O~xd� ��0���NI�k�J���Dj��Yu��x?�!3���{j�85�"�fB)�_��s8zb�@�ʮ&5�:�����_/��H|�1�i�R�oFV���@�ܫA�=̕��ɬ�OzxS�?Υ�_���G��\v[�L�?7��?���"�i�qCͰ{����}�x�|6;���K�Z*�T�|â	"S�����o�F%n�4j���9����T��;���u�髹��𲟘�#��� �����7܅�=�w�0ݐ�kU?�����������#�򝶱�_�Z��t
0H��Q�n����BZ�b�Nm����c�I�>�.�K�
Y��-�B��̈ђwP���S%��a��0�'R�q�c'�r�G��bl?C.EºKX7U��Α�{
�q�_D[:���=�A�So����;�Q�g�Hh�5�/������:�2��ӗ9�"r��Ԭ��'7"DD�H�Ć^'��jj_��h�������?��x��]k�pŨ�x��b�e�ɉ�z�5w
v��Z�g�V��J�-��R�~���M�x�45�	bY�v�����Ī;gO>�/&) 9��^�dƫh4�t��e����8r~��*߳SV�*���1�����.q%���-��e,�	��L�� ����}�o9���O���,�����2���ejPL�1Z�ބ�vwl�"�1.Z�Tev��T�	+�;�1F�+/��>y�M�D�S��ݞ3�������q��3�<����4T�<����1Ě2y�//�ђF�Pq����خ���aw�=���pg���ʘV�^'L]~ѝ��݊U�l��5q�Q�;[�K�YI?C'`��V�Ȣ���e׾��ߜ2*��[`(��V�OӏC�*	v�/[�	��O�u�q
�Q�[s������ȭ�OK���#��ϫ�,��'A;����{}�fgm��*<"<�peǈs�R�(���G�[!b���+%�C�բup�©��!�ŹC�����4�]eQ�g
:�?� X�e�MO�p� �7
5A�����n��9/D�R�;:q󂶐�>6���V�:��1m��$�tMoR��dn�U��wZ�&��U�m^S��T%��i8�P}�Ԥh^Tn�&�ºB��b����Ƌ�!jAȜ9`�����Wu��	_����j�p�mfC���C��d4�F���d���������7���:�������Hӏ��鎫��.*v6�!����L��£�!�$���x�xI������s�=9�צ�k��ܨ[�ģ@�vzcŪ�@&]�=�2����<�ܺ���+�6бQ����=�CX7Q�@Y��� _V�)ΛΖ�]���8�Ηs^u[��,�T�#11��j�tW��Y�yo���A�#NJ4�\���Xȑm�\7�u�`�dCI��y�������\e�)�`s���*2��Wڃ��
M���kvyPA�-�s�GӉk��@���/"ݺso�f7�!��$�zH��EȰ5Q(m/�%<�GbZ�jʠ\��6�d�F�XJoZ�i�:�a��1�Y��HR��X�y4<Uv�5���x%�u���x�(r���<K�y�Y^c{��N�7!m�b"��n�Q�ߐ���v��*t�sF����е�I�߽�i�Ch��F�oL�e���Kl��@j���]�6�A���Z���f4�`1��8�PD��尖JJ��k��2�P��gNd?w.�QP�D�+�I�>��M�8b��9�8�9��]Z�kRrN/�}�W
�_�?�;�)�<��Jl�(��u��t���=ѝK��,a	�T���5�u�6V%��m٧���r�53֨���w1B�7���ħ1�������k?��y��*�����`*a�Ĭ�Q��� ��v�K���(��,#Kc�3�p�)�-�d�ԍ\\��!��I4A����\��rPZ?/��Y��Q����n!&X�EN;��'�6��"�����)�9��x�L�z��yoA�ɝt4׷f�Q���%\��ez�GO�/�3類w��+��E��fZ����}��0�"7��A�Hr�	�v���E�eH�B?�4h��jѕo7��]�#`��k�z�u�Q:G�`�9�����ƥ���(R�(�ej�2ɂ�>�����.��ջG1 ��?%;���R���n,�u/I��6���7��.�s�=8�dkJp]#Ҽ3�x1���VV��(��%�@��GXv��#�h�@����}_�<��B��b��f/��-ټ�C4�(�{�1K	*V���ҖF��#iY�'ب@�43��m�:�(=�_-����`����a����tK���.�Xdӭr)�O}ݨj ��d�d8�v����l;��k̚e�������Qf�+L�6$V��f6�����`���u�z}�h3)�i2 �/";�C;��}��3�B۞,�2��j�\
���,�����iœLBI��S��tu2�ۉ'1<�>�&�����3I���mP�����%�J�s"_dM	�+yC���
J!}�������a�M����;[&W�Q�Sp˭��m��{g[)���j�RڮA#�	2�k�p����ųυ�9^M��}���TPEľ�Z�Q�>DD����vU
bXfR��r�=]P�)(����;�|y�ǂXB��I��V��Qn3��|�x�f��*[F4YcVhun��D�}�!�kN�$�K�X����XD�狨��ZJ�]�Z�J*i���Cs�΍뷒!8N&�Bi*��8�m;ur����W5Y2C삏���.f*G�h��ߝN�����é�R ������:wK}S ܌ �*.8�����n� o"�٠|#QٞPɷѷ~6����?h��#��bw��n�E�	/~;q�=��ʓ�}�]txm˛�����}&n�}��q�k70l�/eR9�uY>{`맿$y�B?�wjL�!�u�ޏ�}�ߋ��1����?��eA�\�5�ws�� [�~�oY��-�{D�Q�mQ��N�6�dvqQ���}�����"��Q���};�"��)�e�\8�m���ʀK\g�n��P��`�]��vb{PȠ����Iz�S�t�#5_rMČ�!�q�qvg�r@K�k;R�.��ȑ�1�X�i��`��Nv8�1؃��Y^���1@X��vfz*�G�6�����@?WgyB�gd������o�,W��Tq6�$~3Cp_3�N:��F�L�'�7P\Ցt�g�TӜv�K�&�4Zϩ@���U���z�>F L�5�I?壬���@@����ˠ���l��UQx���x��`I'�~�z^�e�i3�=��ƕ� D�ul�D�pD�gڴdl��$�&Z���c�`@�`+�\��_�/.T�bBEL�<�g���KI#�-i���?��t�tE�p�����o4�Y�H�W���}�G�	�u�<�(S���s\��6?� ������nS`4T�5;��������`�1a:��@B�V�������wW��Ka���e,+���������ڥ����p���+t�U� ��6�ʭ�\.��Ǡ��o����m�*��9��s
0m~�v4�6}#T@�s���`�p��\H����l����~�\��Y:R
�O}��;�\P���U
���V�GYgn,˂m�}�V�E~����H纎���~ܚbx������2�<�J�60k}T��Kɔ9�����wc�W�����	W��t��;4�]q�zp�k�H��o,רR�b4��qWP��/&�ce���x<���s�Y�<�E�w&m�W"�q�H�Ma^:v��Y�H�>-�iK�S�2f�l���e���_���Y�AΤ��ϵ¤�T�A8���>�n�]�Ga�b�.��_�`v�{��'D�}�5�^��u^�����_�����ۢE�+�!�0�I����dF�������[t�I�+<�dr$�a�T��4�iه�K^c��5��wŔ��D�U���r�go/�ϚD�Z���9�KB���}+j	�K�*qF�&�՞�S+H��pJ�۫-�A���&�[�M�Qe�)[f�TTA�f����j/����Jă����N[u��U�U$�q���n�!�E^,��[/L�wn�s�ڒ~<-��F��ZLm73(�B��9����1@��m��VzBc|���5J
F�j�����=�q�͡<h�Gm~�����k��OyAh>\�~5<���>M �0u�P	=�Q����^H��-u_ٚ�r����m}Ӡ�Q���S9��en\ 4��U����R6����xG��9�4�l�%
�y��� �j�(!����fO�Za"��C5/m���A����p�Y3Iݩf	W!p{���z"m��M��+v��n�%̜Ӡ�LF
L�Q/�����r�F��_��V�/�U��Y��lUd�[V������>tr"�u���ǥ���7�T�ǫ9���*{%&o��"���Ԗ��k�t�[�&�u�/��0�ј�wX���c���.yZ�P���n��-�eR��o^E��\"�����5}��E?���f4�P�%dC�%��wn"Q�?PԚ?%1�����Wf��SWq4b#,����Z����ʣ4-P0zcZb��b�Юo�����=ⷐ��4�"�u�<"���=��!�f��ڀ�6?���Yܘ#A��^�Z���7��$Y������O�
W�T�
:����_dW�cm<$An���i�F���x�.��A�H�΂:��6��΃�6ʔO�P#;�ƴC�=;�=K�UŒ�-��Vxm��}��y;I�:���Ά��͔l7~(yi�����|�}��o�n�֏�`,���Z;	o0�ٝ��>n�h��ؿ��7W>�֩N�M�-{_� �񝽽ڒ�]g RU��fl�!|�ӳ���MK��h�D�9���4?��>�k�flWIZ��;$�J��LS����O�A��R��V��ϱ꽍��G�)���<A���@#�_җ�)��ܽ�nù���7�v�����3Uby�³!u����FY�����h����í��j��˳�O�Z'�X�Վm��&�Oy��A`;���9�:��y�x
aE��{�AW���x���V�����4��YiMj�w��@�Ns"��Ա������l� ��:�,�e�/91�ź:<,�Ն'�Z��e��o� ��bVÇvy�ʌ��b1A#i�܎�T�%������ w����%���PY�8[k[,d��L� `�f]���O�7�w7�������;J߷}��I����č�Ty��T�:	$p�1'88��з\9 )т]����Y ��~��Q�����r]����+^��r�*8���Z��k����%�N�sAߒ�b��p�cP��Ex�H?�s}�o![�8�j!���-N������>�OZ�n��S��mlѢ�H���O�~��lle�.�+o0����%��:�W�'eDu������E�r痄FЃ����D�X������ӳ�>�:>L�3>E��ho 't�v��K�_�mW�>���{������5�g����^���	�^7��>"
�Q���𺑤�� Gf䨪�ziB*%�q!��HwP��(S�ܝ۸��	 4H嬀Op$HR����=�v����f�q��:@�Z��9����t�������/0��W���@ǕNJPP/�3r$.|J���6�&)��N��p8Dj#͆�A�gŦN�2Za��(T3�	@���/����m��"p�B�6PCh7Q ������p��A�s� ~�����N��5 �f�G����d��FA9� 	u>)h[�zfP8a1���?R'!S�PJ`�6�#�*+T�a��&�%\WپF�5����b)�i|p��*����ZwѸ )E���Gm��&"�e��U>_�u���'Sݚ�_WG��9*[��n��Ā�MdI���K(�-ʖAЂ��8�=���+�^Xت�:{\��Z�c�m��'�1!"#7��]7\�,������p^I��	w�kHzw����Ҭ�ȩPV�ԩU�ᢉ]��+��E�WOl��_5��$n��`��ĕ��%��t����Y�مٌ7_*���0�zg�!'�U\�����(����5��NfDb��� �v]���q�/.W4���6�2�I��j`�~)X�F�I>������Wër-Z����H90��%��nT�>= B�1Al�6���4���#y�N]x4Wf?GN�~(V��^�7�P*|a#�(�8Aм��9 �����q��,�2����1&٫�|��h�Uq!AZ3k��<��"E|V0�����f⟦F<������O	�
�Ϯ�,��	�t�d��Uꔝԟ,y��C��'��`nAm�!�E����k2I��pc�2�9*��t߸1�	������g�'r��DA����B��0��,i���'^r�����J���N���)�q�r����W1���
u��,?�^T�bߧ�G\��qx��d��ɍm[I�6�oҦ�{,l��؟;��V¶DT[�������4 �7&2PMx6i����yj���0�G�Ro�i5��f&��!��a$���k���Q.�g�ޯeQ5J�XE!W�'瀽��~o�D{<7�U�þ��	8��������P���`U�[�*q�mZw�O�{h/�\-& �!V�):qD�_��(�=����G���m��~�h��������Ŷv� �<�UBJ�0u�p�dsU�����ne�zy}�\�il�\̕}��SL/X/�V�_��S>�c��90 &��G���+��c(5MQNeR$�M�G4�Kba�H$yD��Hi�3�]��j����'��/L	������{<�2g�g�N��UM��bm����F5ΐ�A��<?�n6u�o���aOa�C�mP�D����sXK �f�[�E���X='���fS������_��@���t����&fp5µ��,؅���#ւΧ+����8p�p�A}8�Q���뀕���������3�u�":��j7��K���Bx�$)s[�kc�1�
/L0�0�b ]/�M'm���ݮ�hH�����wc4��1S��]���0*�,|w9�����e�+��î�A�M�Ƹ?�
��|ْ����l�}��5lM3=V�"]B<��e��ÉAYq=Ed6*�l9�W3�[o��������)�+���Dw��e+D&y���a�Ki"�՟�"�U;�Y�1��*^2nY&F�ΉBG9#�Z2s�_��#�p�X�}�����y3��x�#L��A又�[���@f�Ήl���L�z�Jg����Y�>���wic�-�,�S���J����Y_��"�fƬ)+���V��P�h�6��C/���@�?� 5k���AW�_�բ�С�RM��ur{V�S-��0�U7l+����돖��Yۯ-W��Vʸ���(��ř�)��x�K�V\�P�%jv�7��M;^�©�����:��C��b%�����1� �k��3㶬���R��s�*�]WB4T�x3\�	�ށ
(j|�=�݇�3��j��^�����_0|Un�-���ta���dŰ7�U�+�f"�!V_{z�Vf�Ƒ����Y,�)	`��CFf��υ ����zđ".|�|L�V��M���E����l�I�"��z�阘a�t��K��:�v�m]}i"i�����}��}SXP e.��Ҝ]mA�rKԌ3�(�X�ε*u��l������.�ɓ�=S2-�NOi��J,1�1'w�
cJ��c3���]<�6?>��f˲�{���+�K���G�|��� Y?��MqOclq����0��'�4�P�C<��z[Ɗ0�R���~7�tM�wQ;�	t�]��;}4�< s���|f��:�Sh�~tJW{w����(gf��eA�jJc�;�����Dz��~/��߮t��1���3�z�N��	�'�_ȹ4��Gۢ���E�q�X!0u���|{$ �{wb�ɻm>ɘ�*_�IZ���8#�r���Ó'�� �Nk�V�����h)���e!�~�,�xe����p������.��6�l�up��g+�V ��&'�z+�R%�<+�-�n����`�`��/^��>����⇓�O����+\pŜN�Ue,2Q7����>v�M�a�d��e��T�-;[����J�[�Fju����ga��w�A��I�S��N�uN�#頼,�h=̵rV@�Uu��X�:����Ӻ��䙢���)�S�fZ~��p@��9�6|V��|�=_:o�'}?��C`Yڻ�c{-���0��[�7n?D��k7��k!����.��7������-���D���+��,��9�Z|X	5��I����}��k���C� L��9�9���( :J�]���c�̪lY�	��ˤ�#�<QJ�uRh=�f��h��^ף�#όe���B	ol=�{�b}�O��%e|E}r�<�e�Zrδ!�n���h�:ݟ	*="�-��sc�C@���?2��G$D��5ǚ�-�R,:&�\i$��ܿ���ܳI7�����Y��O(�7�Ŷ��Ҭ�-@�:tM]��ws۽�%��#NN��|�o��ݷ��'��ʓ�Y�H�Ŝ^���hMD������Eь��}����z݆��	�ΐ5�yu������?��f|Mh���C�*�&eA�\��VPR�U�9:����<l.�$������+u�����X�C�∴C�	?�fBb������?���min��d�0����`ֲ�`(�";Y\	�����~ΤtD���ѥ��젮1����s����/���d�EQS,�Q�P�~z��ŗLo rtS�\Qm�N���<�v�Rd�p�D���-`S����5��/L}jGňA�|K$���q��[GsIZ�w���a�Tw�<��EB4�wj#�����C��׼��a-� ��|r�NU�ܞ"m���`��D<� u����-?p�t\n�y.�7�hjụ�>���F�L�݉C6,و�����Ƌ������2�&�Q
%�U���J�ĠK�i(v���%.�4���{L�\ħ�S�|�_J������V�!�uv7[L#�";�h�~���Y(�=�����Fjk��g��a1X���{���q5�9�^��h�޽��لBҸ;��U���C�&zVܰ��<��ʑ�~VCA���l�º�n�tqgLn7f O"�sV.�O�E�x��GaW)�����)����:ɑ��т��nV�������P:1h|�?�w@8ICa��yܸ<�"�i�HW��GCFVSFL�K[�I��r鼒�TD�7`wB�LX�.��{p�(��@�i6�RSSг8��M�R>	�kA�<E
��Wj��=:���B���b���)���]-oqUwe�#,�E��+�W�j<����TN{�u��`ۻ:(�)����E������חL�-x�T���UCQ�I.�K����9xn����n�#fg��ʤ��
ӊ+,��w��W9{(�3mp�H�4�P9�u���Ns�MC6�	5`�+��V9#	����K�'V�8&J+W��`����p$���u��;�>�N'�|���?ɯ�h��q����\C��:���:w#�	�����.6��Ǭf�@v�qs�(�v1ae�F�iǕ�$�{~X|�	�O���E��w�0TɾO�+�`�����r $RNƾ�(X#"G8�Ww�Yi��^�j�I�ނ ���R3�G��5�븕-����~6�����so/�ݏW�H!���e��E�U�Ц��4�>�J=��ĺM�s6kt�WU��)�n(,�$l�Dgd�L����PV,QP=�!,�w� `�A�Z��~'�p��ځbw��D����ɝw�e���A�V�AD2)�c�ܑ��]�1O�<Lf�?�7�FCȄ�{�� �/�UbU�+�������TUP9T�*��Gֻ�ҫ�� ���A�3�g����c1C%���L��o��� ʷ�кW�Q=N�l�?�ӨV@b*k���j�@����{�ӳ<v�|�buM{�-mR�p�>][��BNK^��R��ҙ!�F<>�_t�7Ef���t��jT��ܺXm/�+;&zV�1 ��k7 ��/�u�#W�V�~`�xU��{v��؜_Fv����&ݕ���G���x�*����QY�P�?I*B�[c��D�M��{�2u�N*6E�u��P��J#��ℳ�K����P�J���a�r�ې���~lV]�=AD}��FX�����t2�p	h�a�_GV��%�9Ak���s;��^�����m�;q"_�S�NB�O�����bM�=W�&!^��;�S����ͯ�|�l����hjmɼ���G����@�=�Mw�{����R�K�����`�R�n(\�_���/1�;��N��%��(���]F��3Y'
cl�� �u������jY�'���z�V���q�z.�~�5>�@u<[�%Cۡc~���'��M����.�맡�^�2)k����!&�bC?�LV��mW$$��]%:ĝO��cԷ�6�|����a�2���l� �%Z���Z��Xt�q�|Y�\����9?x���������FW�M�pP�ޥ�����H�W5�.Jc�8^,��mŅ��F���g ]��]�>a�!�cq�1�ex9���#����$�ZMڗ�|b�R�lϭ���6�������Z�;���c���T �`9f�dh�������sY���Ĳi�W��D��vNjn^"`��i��0�H�Ls��L��'�ka�"q��DYpc�����u��t�r
�?  Ꜭ�hi�{�����yT�=:����9������>^D����?�*�~jc���6/0��f��ҋ���6uU|�Q��n#P2��:�;�i����nP�rb2:'Z,mw?����F�����'J�@R��M��������Q�v���%�bs$�'�2�E����Pr�-/�vG���� ��C�9(�c�t0�`���W�
,��!�Rw�o��e��ٍ�}�h�17�U���h͔� �[-�t����)��^^���OаXQ���f/Co�9=S��%�[���U� �w���F�p@3-%"�k�PQ~]���7m�������������laWk�⑄k#��4i;��URJ��Q���o�b�(Y�����J�nB��m$�V�G��P�7����b���қ!��A��-xB����6	�ɸ5��a�e������q��hq�<D�,����.l�]�(o�ܪ���!��xY@ٓ��P\�#C?S"`��� �b{�:�MG��]g���o�A�s�aՐ���E�;�)9l�oN���R���;-�7+�_guH�ʼqm�z�Dl�ܙ�Q�uv��n��k��p��D�� �n��nv2	Q�S^�;�zW
�5;��S��bŭ���S�M8A��h.���z��W
U�Q��I�ķ�;2�%�F֡��o��B���7�s!�C�w&��P�e�3��$��LƄ�d���%��ʖ����&.��ڭ��68��u�����R���8uӶ�p$�Ռ*�vQ�ׄ����QW��K�`��B�T-T��,Ў�0���
{�Y/4)s��]X2F,�a�!��5
��~�z����1�&ۀ�I`5����N`60&������^� ���������#Cc�9Wx��b,����V�b!�v�<f@�H� G.��o�o�Ճ��Z�|i�!��8ǰ�=+uD"�T��9J�� ��q|c[NfE]i������CI����|�����=ͨo�!�����V�0]ð�j����b ��Nқ���a�� ��$/�y�o�|�05I�Տ��K 	���6�R�E�����?w���H���:N��F�3��SI�f��_��5S����>�c��J�ܾ�
0��~jQyr�z�rW����9�OMST�o�ti��X��<M���_����Mw���GsS'��A:̢C1h
I]�Z�
��R}d�{G��'w(�W -U��L�&e�|�	:ɉ{HNt���e�A�*~�6J�虲�cQ!�W��4ō.��ɕ�S���<zm�v5���h�=T�b(�Hl��q)c���2��ցm���5#i�{�Ɓ��2�T[Yǟv�k��F��#}���L�y�{@l�Q�J�ZUt�-��l�ȭ�cZ���u+�0�5)d����i0�0�cL�%��މn��lG��*����(H���ٗtzDVs_Z6T��$���xiɟ�;Xk�dů���V��?��Rj��{H���].�>�&]c�*�Z��E����]��� w,Ey�x|Jt������wF�'���7l�Ni��&�I���K��N#1<��pG�=�}	�h�r�!T]�x��{��H&"C0���q�J�cmlOǗ�u��,��A�u�����@"����Vq6M��f�REf�N�ܿ�a�)������ޛƇ2^u�x�t�K;��Af8�	S�	�"�t�9�)�F4�����ң�^iދw�y7�
x$V��Ծ���?`�v>� "�y8��ɎoR>AѤ{��=��r>���,��o� ����8�<�\��x�n��`��@d�i#&KlI����_gJ�MK�'�[�#�La��μ�i�+�T���uy.1�$x�jԾ!�X��r!oO���R-v.��Ҕ���`�U��"�}��݌�G���*���G9�u%N(���
5����+s�o��چ���%�|n�?P����M��3Y����4uVrW�4��[8G���7��یOnt�	�0l*�॰%y����,j��I�@�я>�r�{��l�r�V�C����4��k�C��X�k����x;�oMG$y�˶w�ƣ�9.AD��OeN|&R=��$K�W[3l�'��8;�.h�΢z]���f��JРl��#��1?�W,��6p����I�Sϡ�}�3�sG���i���{�2ʊU0�8v]����꜃<����/��cR��e� P����$}
봹������$��S龿� s\y2�F��a��S���j0y�z�PuF��>Zk�>_���(��lp���@���T�����!�r݃G	�XL4��]�f��6!9Z�ϲߙ�f����U�����]�棸l��Q�D�kTXJb�mdQ!q��#4�W��+�W+=v��U<��zF�7���d��]��J`Z��/�Ĳ�#`���EB���V��N$5-.zEsk�-R$�{��|���n�<M���L�f GX��R�f_�����d��U���Nk���=2ӘΣ�ڒ�o���v8%o���GW����$��KU���5��Ȫ�3��6��Y"������������� ��B �h��������0U>v���n��xBu�4�mU�����5d��G62r%H�O��:���e���1����wk�y)�����У�;xG(.R��r�jLUO3m����UTC�[ټ��!��p�KD���Sƌ =�T�(#�v�������Ck����#˘��0+ԉ�x�*��N��|0ր�e(�7�����ةd�y� �PW����z&�L���X��j!��A�'����ؔ��D�^C$�_b�R��e/	������eJp��ز�e5^2p1Mt�՞�)�!�Y� 
�Uժҫ�ӂ���s?`�
�"��	����qJPuH�rձ�G/95R1�A].�ӌ�����|�Lo��N;be�,e6�6 !`��2�<
�5�}���l�����P�
/>���!K�?�v$�R���Ү�"��uy#��*��_�טAS����A����:�����ؾ f(T3>6�&�3����A����8�z�9r���noP��z �-�>-��Lp��lk�m孊�^������7��̌��@8C��%z���Ӫm�W⩮ߖ��G��'F�9)8�%��Ů�m��^�d�Ǌ��g�����Fs���ۂ[��>�َn��L�)i)���r�w�Nr�Vhxi��"Ntn�a��>T����R�{zS��M%6�d�
�1�(6K#�I1�� -���P޺1n ���e+��M�&r8�gv�ԧ1�����G�m6c���Ԫ��T� ���&�C�@ʚ�k��i?�|��a(E�-���6b_����w���~���z��)�\�p������V�.�g��4%a����� !7��N��lo����|*�Z�A��յ������|DY؁��Rż��($P�o��9��Z�����~�ˍf�� R�M�����t��έ��MC��D�芾Y�{�O�k&�&i��⋿�%�K�!��am�U�}$�h%�B�����d	�Fo�e�*��Ɓ]�R;}h��A�f��!YJ�6ޏ[�S7Cb��P�
\��G=�t�^Ը2T�rk�)p��E^](JX�"�[eb��쌯����F��l��:�y�t�/a���LP�е ?Dʥ��a�)�Q�^�,��u����.�k.�<6f+s�ª�`�IꕔP,��B|l�n�5��$�;�s�5�w�H�g����1T��1���VQ�gsOp�����$����N\�u���8�1"�
Ʋ���@��̧�Qm�c������k�˾&AMօ�S�D�d�ʷ����M`��\v���ގ2�=L�a����e{ͬC �ӵlw���z���F/���#���f�w�͌��.!k^�L�UF�%�KCDy���?��M4@���8W�1���ǫ���.�er���&�Jy��
 mQ��D��jq�u�RV� Cp���j�%v���5�R����'x����X57�0o��엺�ݪxZ�#���F;���ɠ�G��i"::���V�
��zw �"}���~qYՕ~'ͼe)OH�1mR~e1�0Ԫ�U�d�캴t{�g@�ȓݒ^x�-�p;��֒ߜc2-��<u�����\�-3���� ���y\��-+�Nq���J��*�+/�0^/Bp��O'�L���G�8*����P��N�=��'��>�aM�S���,m�����{��}�ǈn)�_��Vhw9�k��K��M�U�����2�,��$:�Q��q( L�Ra"�����@�~����}AǛ�Nxr��w��H��9��4¬�5!�db6w����*����)�,�<zꫨ�	zH7����	�cN�ӗ'�KO97���暡8�l��W_�yC|x��՝OD-�n.P�Iq�(I�)���������ىx�{�A"��IOy �UBY�zn��v9��_���?�+�I&�V�k����??�b�/����@>�u����ժ�{&����
��~?�Q��WЭ\�����W�{ڠ���;�Ԁ��H�g��M�"T��^��m�=~�S�\�'�E��ǈ�<�0k��ֺ
,p������i��O\�%v�$�[�HԤ�_�	t���2���&d�����[#GK���CT������[��<��ez��7\o����_.���7r��asx�bP��؇	:c�O�M�y|^��x�_Sk/�����;�$\Th��Z�̶�x�}�@�D@2�$�������Y��lL9�(O��˙C/TJ�����S�,ȲoF�j�BGʯ
�2��e� Y pwl{�$�����^���!�
�aZ�:_���M��4.	0Dd��<\��{<����2U��p6�C�8[3P��9�[�q�h<���M���f׿VڸlV߹s��kt��*�k��B���
��X>X�^Ⱦv������3io�w����,��\⓫KI�o�(�/UQ�-ɏ�@���p��>=��xt��#;��r��U�Th�����z0���/`�o�¡ث�S=�ra���]�鼆-gXػ��"|d���H%8ʞ��~�ܠ�'�HU�Z�H����ȥM"���ٓ!�G4>���j�gd��OhC�P^n�bg� �Ϟ%�8��B��2�+"�U�}AtA5P�oZ�h�,M���5�����>u.}��谁�9t�C6�o'�|��P�wU1��[�����|�DL&S���XK�0�Z����$~-zo?�`3����F�$s�j$��x�7�* �,09��Ԝ|��`(�%����[��<n>�x�8�������,���-5�q���`K�$�3w~�Y�v4�� X��`���<.��V��� h�Z���)�_�	Mf�b��i'����L��Kκ�֩�s�����^!��e�z�D/#����L�ßdn��kl�lI��}�k�PK�0��j�)v;x��Gʎ&��C9)b5�����y���e�^��"M/�z
Z=!�2����	��L��azWi��q�cY�r�%;��|d���v�t����4
aɧ�c�#����r��J�kS��q�B�7����Cw��%|�x���(�`AQ25��vjr��$b�=Ib_o�R3������{G��j���5���m+���ͮ�J�y �Q�ںA�|t+j_�P��+r��E���)��)��rH�)���o��pd׀mq,���A��6԰4`NC'M9���j?��a��W���km�&S�(gS�����/<�^g� %ԫ��X�/���Z�N��S����VXs3�R'[��m�;��� 7[ }�����gӠÁM|��\go��?���RtK{�W����A� 1|.���^��v7U/G�r��t�\_9���sn����*��F捚��<��%�e�H���������l;���`�W�l[����g�HA}��UF�X�P�����ᯐư���꺪b|�F��EM���Jm�)��] �ڀέq�Ɖh��Z����Zw���J,0L)��&u�\�/����m~Z����QZ
u�g�F��,b��-�nkeԑ�t�,-�IG�c?��U?��?4�Ω��*5MZ�Ϡ�(�+Hvx^�x�ήs$e!C$b̅��8���Ԝ��v��a�T��w3Jf��� h�͓5�2&b8�/��|E�y���}������d���xr�e^��T68ANw��BT�>�5�X�i�\�i���V�)�TW!k�Ň�F1�a���+���}n�Y��'1*�eTm<.�>x�
&��bNזּ�y��tp���� q��;ΒC��ӫN�������^Ŀ;=�ׯ�.�P���v��N��vt��N�n	3��� ���4mf�N�����<;��[��F���l��n�ɰ͠WJ�g :&�Wv�޻N�4�+��]����}�@�OX��$��վ�:+bɷ</���fE�2�X$<�)�KX=_��L0'.	����?2/b�y�kl�yp��Ջ̲ar1Y©�~B��
���IA7r�PL�B3���������
#���u���í@dl�&�ӈf��c��&���������VPX"�}`�,$��Zt���D��@�4��U�]�p��	�x���B���ᢊ$��{���e�__ߓ���jyX�5͐g��� �0�h4�ɻ�&bji����0���3��}��V}OL��<IN�|7��vQ��9�p/~r%�Yڜٸ������
��}fP$�� x��`�����e,L��W�1c��.^)�QD�ȡ�ю�/�l��J��J��i��^{�_$e�/��
��⎌0�2�!YE��$����0���>����AOg0y��Qf�6Ш[fF��湂����F��Ki�*�d�c�ޠ�3:�h�������:4�_(�	X��$������t�+��GlC	����5��v�s ���\���n%�:JC�+�ٹ{���7̓���|
X�PR��BRф��8��df� �$��������hݫ/����oכ����қ܅��v�-5R�.�ҥ`��nd�7�"���uN3��n�;��e �S�]�*���>s8Ӫ���(�y�\�	���&U��0�`��JwY8�`��0��5N���ُ��������,]��(�$�Ea�_������^v���<����r��[�P�m�K4cؠ�9O���4�A�6R��ΣjȊ�1X�$��_�c�b��ȗ�4N��p{>(fۘg���6��Z�H\����s�?�;��`r���q	&7T�l�>�`�ρ�AS�yh�O���ޗdx��3�U��,���`��s��z%��滉m���QWt�h;���P���8����'�˵{k�!'�|�����>`P]w�<�D�?QĲoP6��(��)ea^L������z.w]���� �|'�>(F�-b]| ~��\$�\+���lk�z	�&��9�ޝ��,B�۲Ze�G]Ny0����d¶FR�vᆞ��婞aֵ ��ψe�C.X}�4v���H?��>��}b��S�H��9`�H���gb޽�=P�% ���G���"���ĩ 1G�GV
Ew���@@�.jo��k�KR-�����ܠ:���j���y��U��~0���E�C�W��������׷��¤����F��yӲ$�ͽ��=�����@7�,���:������&��@�	��R@�Y�[�ph�[C���K����t#��nx�X�d��r��/	~z(��9"�Sc��t��r�PC��r��)tFDDؗ�D������E�h�U��5s�z}��6Y� �Bt�VQ_vCQ�#D]��}��x>��d�U���C�~LXY��􀨨�`�2h}�KԀ��x.c�C�'��㏧k�l��N�cz!j��/W��ux��zQ���:��ɂ�G���̵C|/*����OI$vO.��N�P�ڈB
��"�0��D*�>U��d�
^�yd~��S������Z�S�@����>@���w�;*��ex��R�in�ǌ�Z��"�)�!Qe����v;"ٖ�K&*K���%c)�����.3|KXp�h��i+��nׯ_���K;1��P����|�i�F��e��CG(;�SGmF�����Q�Ӥ�w��?�:BJh�&3�W>�+	���Z��/����?���yPaɒ�[�R��� ���N��_�1��yƬ�r�ϣ�$|��Ʌ�	.����%��H *qkNM?����W��j���8%Mx���M�:M|�Ũ 3���"C�;��
�wɍ�]g鞰}z^�Ȼ~-��ԃ�'�� �I9�ߜ���f'v���].��x3��F�l�9pI�m�eW��/���w�>~�#�"�S���2��N0��4�PM�$�*��Q1'���]:�"]��� �d��Je(E]ՓX�����CX_y/ʓ��@?�(c��� ��"|l��Ă��S7-��6���L#l-����4e�Zl[�n�l+��� F�p����7(��_y�U��K�&��k�Jݖ_�P,Qڙ��8\R�*�V����Z�'m��(O�-d�0�6j�p2}n�@#��Pyx�E��%;Q�Q�נ�Z��V����G�B1>騄v��8���d<���$��{��p��i�� ۤ�{9����w�fN��˳��-t!+w���^WGD��0X�:*��F�GP�����`�3�!f�
Wd��������χ$"�|���P��z;�\�����?�)w�[��F��5fUqu�%�E�Ք�@��#�����V6y�K=Ǟ5`�d�L4�Ұ����,(��. }��dD��@�����R���0� �6J_o9ILy���&M��E������B�~�SN�|�5u���zB"���C����`M��<�+Xz��pJm�ςD6T��"D:��t�M<�z#X~~q⛇-��3M���+�.C���t
��d�����Z->]�#:w��z4P��U�XBo�A|E&�ڔ&�w�
���a��:��hL�5g�� Pw�]�T,��⫹�������y�nJP!�c�6y���8�,4}�2Mj��i!���S
�*Y��PM�5ˠO��W:NX�mP��k��pD��Vts\F�����~��`kOgA���,쮡�Z��^��6�䲒z7�A���W"`�QSaK�(�}�>jն�ve��<&�p03�=�{"�$�ܶy��g�*'62�l��"��d�	O�E�
˴��l>H��F*����Ԟp��;�6"?���I�/ַ� Ԥ�)��S&���x{��*0��3߭�jգ�m�P���ķ9�{����p���-��4^��[�U�=�V8��5��?��ĳ�J׫-���,Hi����l*9t�%~�71\�0G��4�!�_�Z\ϭq�Xհ�؆��P��k?:����h���{(@������,-:0]X�y��و�uO�36��j��.�i�Cp�gx�\w?䘨�Z�'�`!�����ըs^i�;�4{�
ㄬ<2	���Ȋ��y	*�=\�f�hi�t�!���Iyu�B�Ѹjт���w�Dq�G���{�����Kx%.�M�!��x��l����ȀX?NJ�$���U��q\��9�C��Î���Q2j4��үdf�� awr���92�P;�r�d�Y�{�<E �/t�[����*t$S�{�.(r}7z�^7G$�X58gS����������Y.W,���&:�<ދc%�x/�b�	u_���[�R��_�n+��UR-ʡ����.�������
d�����𣉂�L��$7q�ܞUO��x�i+#�N$qDW� �f2@#h�/�����Z��x�������:��E�e��^l�J�<Z6&�_�0gNZ�^��	�)3ȥvPA�{֗���u�r�6us'�]�M|ïU@����Vj��6{O���h`�H����'c�
��mJ��,�C ���Ǔu�h��&�v�Ч�3ާ�Q�!f�hV�ݨ���tI1ب -��O��&Ɲ�`OW3�V��+78PQq�����b��8V��6�ӷ��ώ��y��0|����~k�W;:Fo�	�1z����4ڈ����+Ui~���Ewd�8��%��(o�ԻW;LĶx�d�0�kZ|��wkS�� ���XG���G����,Z��$Ɖ��)(�������EAEʛ�P ~�T:�k��o	��D��&Λ`��>�g�F��-���kij��h��P������yn�� ���9Թ��\�K�:���lq���O����VZ	P<L�,�'�:��-#�n���X.H6:l؝ ]_g���#j��"0}v,�ph �g��t=��zoiӟ�ʮ����gU��D5v!�*d�˧8?.5Yi�ht1WK�qY���8n��q��>*�6(�$"�����8K���w���B�u$0�h2;�}�=B0�"�ƋӼ~�1�f:a��Iu����$��s;Tm�$�w�d�^������W�5|����}������A�|U�mc���2�u��8����u��܅x���_�19� ���X�� V<I�X�ݸ�;����C߶a)����k�;Pom]=��{��,��%J�g�E���.��.�ėfz158��٨�Gӧ��]ܸ��	/��F� @��KR�)+���,�2�k�tS���E"2�떂h�
;	G�g�:�k�s�-8�_i#	���4��2!�h7j�F�h���<�A�����>y�Zlk����л�д������΍e	^�.d�U	$��V��>���ݦ�D	��e� )%�+��}&�ؒ�;~׉����Ё����Ҹ4�2�f1 � w#�bx��rj#Y|W�t;����S�g��=N��E�?�G�z��e���6�4"���u�|�!�2Y�)���}XD��U*ƓC�D ��!ET��yP�����_��ai}������:���F���;�:X0�ϒ�XՆ6�S9�*ؓ�~���΀���	t�,A�w��@+W�ޮ���ǵ�<isq��>0�p���Lx&6����'|:*��yt�z���x��l6:;���2m�|h�.�r�33��@s �$�o��6�+.��}�wW U >�o�"��x'h\�z/'$9#���w�YG渏�~p�J�	����������vV>3��k�	��ҧ��@Ǫ�?�rC���Ґ�+���=���tEd�V�*���5O:�͓��Yg�ë%�ҍ���
�YS���D��ʆ��%� � �8"�}�����e�xk�f��	X{I��e�]�~�ӏyIS�< ��p:�S�|A&q�@kx-�V�AU&7��6ˆ�	�_ܧ�;���`$c��&YÁ�r��CG��wR�5�� q#fKwg��X��C�X��_�ׅ�r��4�}g���ޯݔ$3pE�k\�՛et�@�"G;k��ν�"�r�W���o��j34p?�h�:?�&As����w���f�p���'Y�L����Va�#�h��|��v�5Oڢ�9F�0��G�%�`���ተ�U�Ί����2����Yf9��W�����~/�M�4��K�hgg���	�C�hi�DRy�[��I}WT�s"ݶ���yNtǍw0OO2i��U�����K��9��ӧ��G_gM�%���
�y�A��k(W��nð�ߢ%�CY��	'�n����oA��
��Y��7��@x�r�Y��w0I��v�񏳚fi	G�&�)�E���)o���y�F8
iָ4��$,q
Q�6���۶g�W��Ӵ�aM�nZ⧞+�{��,@�����Ӷ��Í �����ǚtRL��s��_ u^61�����ņ�둮��Ds�3��D4���轒��4�JG�̉�cCZ�:�b��洎�¬��+?��**�ޖH_�1��^�8^jr(=�W��V=��jO�!�3S�(P��1/:V�q�B)�O�e����:Y���l�">+B�T	���	e��0�����8T�����2�}5��Ht�)���h�^N�K�a�Ǡ��/�ݰ9وm�"3��j�S�#�3h����뗅�	�*��n��5P(W ��o@g3�n���c��:u�&nCJ?5����OP���E���8��wM3JT5k)��uZ�n��i����X��ϟO(^J�?Z9MB�M��'l<��x,Y��d��A3T D!���ݕ$4f��Z-cv'���<�,�o��΋0I~�<������y� %K!�!��Vh���cu��wɹ�ˀ�J߰?���a�^H���h��l��QI&�2�T5�2��� ("����.�I���{�n��ܾ���+�ܐT�,�O^=}:|_�+2�X�����orP�M�%Y��[Kq&��p��S�I�>�[��鄞�T�k&�,	��VH�OQ}:V�I`��fyS������!��r�����2�"�K�vB���'3]IQ(�-�7F���<��y|.�Y%�����uem5�8��׉��j���ٔo"J�ͺ�Ι�q�����m6ᒁ� �وoPs?���MqH{�l�i����(!�+MV\u��c�0ٶA=�>��3��C�����^���r_�%ڔ�85Pi#����si7e���q�b��Ť+�-��e�K�B<����ռ��t�t�t��,-@�{q���:�6f^$wxX�ʤ�?oXm�_R���l:��&�f�z/<H���ƙ�@N>j�A�V�L��(�F||7~m7����^Bg�Kc�LQۿb���T����*�u�B�����ah��yS7o�RX�䦙�}���r"�*��9� �1u�:�y*���o�[�@�z6���{hxq��$�`�q�b'mu��h�ݻ#�p� M�R��}Ĩt�y"�����>��aC��%��]�L�
h��%<���b�+���Yܭ	M�{)�uwi/��R#<
JJ��G���^)2r�);bQ89E��R�~e��<_)��1� s=� �_�4�mt;�Ɓ��-sD��Xn�(�k����BTY�Nٔ-���j���E��=֟��A�M�\�Q��vI�v�N�abf��p�x��*����VM��f$�xڣ�:Kh�%l�����2��r-��'����>�'q��u�Q�mF�0#v}9�� �kN��؂	���m��7AԿg����A��7"�����6��\d"{�b����$w���K ����/���!+�BL]-���k����˕�	ZG���88���0x�eÑN�T��h�jb}��u��[X(�*�ku��MT'2�ܴ��޷��s��!W�K�x.��Q* �a�ϵ�)S�a�o-����`�������IF���j�Z�@�k]4B���c[:�ƛ�7�-���H��)j���΢#v�����0�[�
���x�}w�-�q�[���5���K�(���3D\ZUIf�&zo��������G��2��K#�s&�����ü��n�~�51�EQp��,^!1D�k��4��گ㞦Gm�A��L@Sz���{Vy�>7��u�X�M�����);��}����0Ϛ��k�M�?	y�!H�=r�����cul��~���3&�O{�=�_��U���3N��C>ɼ{���-+@Mp �{g�2ƈQv�i�y8�%\�+�A�r���3�0��!)K�� ����0]Gab��zKϛ���+4�\29x����-@��k'�� �?U��f��Z�;r>�Sr3���-�U���z�s~�f��̞VGeI�J��Z���xD�`�	����1P�N`�o^�4���/۬ �
���Տ�3��(%�H
�mZ}nJ�.2���M�T��=u�kCpڈ1� N�*�;OdX�?Wg���o��p����I�z��x9>#�k��P:B;���;'ŕn{ҽ�@��0˥eT�� a����nw�d5�<��u�߾�Ri5�%��4^���:����4"�a���P�/`F@��3C��o�q'��W]����Km}��������g�7��^�3h�UM�ιq4�M�oS`�y$%�7��ɕZ�X䋩�81X��k���	l/�?�7x���z���_:��0����U�7�����B3y����8��#뜃.�u�t*ar���W�u^ ���F3���~v[�%
�~x�U��s�ZRS�K⌟��6���Ö}8=a��^��Z�	X/�,�$"8w�k	*�M��qߍ�\Fԋ��Z,`�;GF�)$~;��}���F�G� �۠Ms�Pп��I ��+����Z7 M�_�i�-�Ѓ�]��z���0.
^��