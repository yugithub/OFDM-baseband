��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�|�V8`|��+#���z���6��Jڦ_��ﶠ�嚍�e�X{
X^T>D�O������:J���Ў�`�N���|�)�О�RޛTʭql}��DK��q������4��_��/�����f
�+��I�Q�?p���c��	9G���e{6�Zg�А�8�Ou)s`E?�&WK�2ғZ��G��m	!��p=hV�]P�|1���#��c����:G2�e��KmM��|��q�?1��uC5��#��/��o�L������箹m��X�jmS4
��2HQ�|��(�Sw�J"��L-�HUx���!_$��~���=Y � �P� C<�>ල%�#��B9���N�=!/��Yu/g� yt�")�@	V�������?�J��c4�c�6W L<a�d�n,$F9����'�zj�Qu� �,�}����	g��s�w�q�dy^��Q�2T�����U�׿6Tx8/zq�u��9�"U� =�x�
�^�7�����þ��� >0n>��c33M.�A�Г�>D��F���]C=��s�������~�.q�_� W���i�"�+���^)j� �"���B/׿<�I���y�[��OY���y�!{�Z(�LBӯ����P�[.`���;@B�ґ��|�U�%DT���h�,>��K�65��b�/i�����#�VL�@w�wO�Ψί6���1�b�s��V��+V"�І�{$�L�Ɔ�~�A���b8t(�I�*h�-���6x�y�g�J�'�{��g�������M����5��vЃ	�˩�4�
Z��[I�,
�Wį�D�F�B���!���B�W���c	(�A�� k�	+u���z�U�g����m��O�y�̶[�iB����KDǱ���C��`COӏ�1
���� � ��#��S⡵����X�,�L���R�j���'���\�2��<6�Tit�h�8��n�F6N���sͅ�c��;TU���v7e�����Cp�t<Uu�U!ͼ+6� ��T�M�'p�T����#c��{y8���b@�V�TP8��rSM���R�~�/�v�98CR�~qb�|M�d��5��L�ha&_<i������;p����C�ڥ;��^խ�Ĝf.��Ɖ&l�Ӫ�B��#-59;sKe�������Mw���땶ג�q���(E:��g�hY�L�Wܤ�Ɨ�_�fo��(�ꍛ����˝/6��:�N��H��"�\�	c�kv�h��k�����ڼ��39�#!����cF�_����w}�]K9��ȵM�@�QaA��d8P�ه�[^��::�p�n��4�zTҚUZ񗿤�G|�|���j@N�\,�� �{'�	�P�,��ۀOT�R�0%��F=S*b����~��Lך_OOƿrn�%�`��F�B�_}�%�:�U���: �Gx��Z�V�����\��5҂��a.�x����E]YT�����Ky��ޟ$m�p��������Ɋϥ*��n�j�B8����
7\Ƙ�]��A�����;E��*����j��B�������@�����J�8�:��uP;�����
�݂�����O�Z[i93���rR~�~"�3����t�q$�W��Bp�f��:oV�/A� -��6P�-,�V��O�ƂhR�YWh�nVh{�+�I�k�m=��\Q��\�ń0����_����ZL���5vK��+l]�5�;C���(7�E�h+�*�.g�������=��CX�>o�j���(K�}��l<��g4���z�A刟�8E!�iu����5�Ab}�rP��`����hE�j��J��~��&��1t_���Ďw.Vv4�~�`햵M�~�,�'����߼W>k�_���G}���u��B{}-�a(�wF&�N�j���O�7��LJ���:"�����R0���Ch��4|�YI&��&c�/�����`&�������*���$�D7f0L#z@>��� :qʊ��D���P=C����??�)[��99�o_�x��D�Z5���E�xP�zfsE�������O�Fv>�e���hv*}>��.Il���a�y��������,�Xs�282h��#�0 �<��>ܚl�z��z��W�vI��I�a���^�:�.����]����~�ק��
��*)gYL:�9�j!�� �h�E^��F�|�ŃOq��?�*��c)o�'��фJ�(nO"iP�έ�^`��NѠRA�F"����!�q�z���ZsD�ʱ���9��*�Q�z��k�uf*��|����߈lz�־/�r���5��f�%�KZf�L��:R��o��U&��q�r��9b�9��	~�mC�4a6��U6�0j<���3�%"�I��Z�䓁6��C����D�M3d�!��n��e�U�D��"+��^By�ݎR��|
���u=�m���͢�/�/c���uk�ʯ�:}��0���-|i���<��-on���4��?d}5�Zh�6	Կ�s��ԓ��'g��5\ﺘ)y�f�4���\j�(Ȅ����_ul��(s�"���B�<*{�t��e��*;v�e�ϭ�$X�ҳ�'�>o�䴍���/���Ƹ��{�h�Dߩ0��H5�RԶs m��?�ҁç�=9��ߴPY�>�[��x���B���;�K�1�b�p�T`w�*��R�]��cWY�SsK��z�t��8DR��hz�M�Ǉ�>��&o�)Ly�ɐ���4�74߶xA��=Q�٦��ܝ'�g�W�'����ߟ�K���`��`���b���1$�U"X�*GŀM��l��6�C��8a���yqE�����E�Vt<���oP`�>m�"���Ǉ�Q�0G� �Xr�߿��V��gy��K9�\l㱋jEQ�d�~�T�M�1:/��Y�%+���O�BL��4���o�j�Cd�����f)A0�Td�8��S�r�D%�=ǂ�9��c����q�x�,��q�0\rԓ���� A�л�Ț�,T���"$jW �k&��?��R���"�^�'�����1��q.�Cs�~
r`w����CW�N���l�bL��;CZ�,N�E��ܰ����灯���V�Զc�p� ��~�.��^M�����GN��������eP�l��j-�?&��Pv�{맋�D�=��\V�9\�Y�>��/�oK�l2��FE��t��Dɻ���|+y��
��N.�X9c}�B�1�U�y��Ԛ��c�����!w�vmf�|���3�+�pX��-gg��o&s���=�Sr=D�dĴ���?�����դv�U�=��9e� ��A��)`q꫞��V�{��Y������q�1�����$��)�zK�Y� 6󰆊�@��@llӃK`T�ߺ�ܑ#���|pfu���t�Wvr��k�"7�P�/XG^�Ռ���5TT� �d���j��Q���gF*l�G��[2y�q�W*��P(��k�Y�CT8*�����eB	�]�Y�!�^��C���_���I����E'�H�rz�2y
�������]$���ݕ���O�al��O�(���L��W�Kd����.��'lH���E$�g7�O�,+߄{6Qi^*�6g9R��<A��+濅�}hq�҅&���/aY��.��MNw�&zOgׂ��{��}aޣJ��X��p΃%�����X����U.Ȼ''p�O��+E����ڮ9i��Y���Y�;1M�5jV�[`�&pi_������)�s��fQ��E�����G�00����'-��Y�U����{f5ä��	F�D���۹�6m���.c��D���No���c!f/��� ��{Qz����3g���-w��W��V��h�T�,G�1l'q��7�e@�o�����1�A8e|EK��}E��5��"ϔuS����u0���u�aT�2���k{�z��~_YB8*/�	� 5�����RF���Oj�$q��ܠ��G,�xl�/M/5	E�K���7��~��(��Y_LP� +#�D=�tZ��f�X�u�(������idb=p	����$>D��C%4K��7�*{€�Ż�ɝ���ȩ2LCr����(4�[�O?�������X�0l������y�B�宁_5�,U�����>l����v�hO�N�hT��΄VV �.r��n�?&!��k�5���Z]�(֤C^ق��C&ũ��s=��,<؉([F��Cm�Lу���8:�(;���B��wH�ld���e�i�6�F��xTAn�੃h�SY � �_��/�(�ˏ~�H�l�y��`�
'u㟶ʪ��5/ҽݑ�|��!)o�b�(E���\����`��R8�#��i�h�;�/��S#�Ȁ���.��U�\�=-���i�O��F�X�2�� UGh+�Q�k��:��ˋ�@v�$�&�d5ɨ\������iqV���� �0��g8�X��hR���T��"261��;������\�N ��
�j$��)[��Q��⣴�$��ǎ���WФD����>����35�50�W�~����JŚ)Bo�y���w�
K���a��g=�j��V�7���*ד@s=gm[�G���xK������Nb�ڭS�`�*�kU%�� ��H-�C��'�\퍫ñ�d[<�_h�\�nP�T�EOs�JG��wHt�b`���������+��x �r�:�Dw����~��Ǝ��8��v��2���j"�.Аo�o�CoȽ��DϺ�Y]6�*�W��y�^�f�4c�ii����`P�O���)--K��H,'6 E˞��yQI�2���b��"�]W��}�3dXkԠ������5���L������}���o&~���#.�A�呲"�X��X���R=��i3�-|�b���cCAJ��;GK�SÏÁMʰť���}|\El��ѭ�B��/SB�O��]B��j��q&h�Ο
'�N�M1�8���	�D�q,����a9?��{]����N	&w��!#�6HG�7	�8�����Aō*�����~U����9D���#��E��P�9���
�ZK�c���9�vP_�[v���P\Vi-�-���9��ܠa�b���neY�4���d�G�4:����tW�A۽LM�i�b윞��ѷ *�&c����j�R���������8?npspy�W,@n_���u�4�����{տ���:���}����}^���jF�� ���ke����\�0�y�VfQ'Nb�n��P�	�Xn�6��'�y'�m,�`�"��Ϡ1M���'�6����DU���ŶnzQ4�n2-�ʱM���1kIa ��r����Y+lR
Zܡ�I&�%�id{���S̺��:�^�fe�a1���)�?^��7d�pY'ē�70���Yi�ؿ���v;0i�3`�.x@g�i(Z��4aȨ��n��'_к1�0Oj��W�ۉ�d�)RH��y]ڛ(Z����ג[��cQE%�n�5�D.�KWk@:-����)���2E[	�↤��{!����1j�ny�I^��}�"#���*���n^���t�T��^o�PST$+����8���pk�|l6�8�A�ƅ�+`\��~s�[�7;O�-"@������<c�G�����H�g��kBK�F�ʾ�3�-��9��>R��M`i
�^0n#��2}a߶�ֽH�=� �wv��OZ����G���\آQ���9��,�$������e��(�,g�
���j̱�-L�֟R"Px�ŏt���#� ��r�)��^$3㓪۴�D�)I�8�),��<��s��!�_^1:ʽgt:��ed4��ݳ��|�r� �\�mf�B3-�j�	::voH�]��,�����~Z�ʝ�?I�ܨI^$Y��'&\J��[�����Yy���΁��q�޻�9�6�W�o)`��7�6���0�]�����r"r3s3�ϻȞ�*f8J ��T#�&�@��ޠ�H(�	W������5�h�Q*e�
e����b��h�����)��$_/� p�����ɮ�m����E�u볺d�)�>���;�W�(D\T���7Z�&�`�X�5E1|N�y��BQ�k!��ӝ����Mwj�G�SCpj���*������3�Z��0ךI3�u\6X��(B$OI��A2��25܀aD�	Q2��w`/ ��s_�za@&<���횄]<�}��V(4�|Z:ɥ� b�)ۏ�=[r��X��QɁ{�S��Y[�.���I�L'��l�k�vo�}���/���Mb����f ���OI�(�>�0yB��.�$&�g�'r[��Z�)R?Lz,x���#��I�r%�R���#��!Ȏ���#[���*�2��r���!Z�4�zi���%�%c{�_Z����������{�����R�|ZC*�`�_��Rf!- :p���0�L~wa��`㱾%�GL�s��7����)$;�Q�	YN�U?��]jf���G��8o�!q>Θ���%^���*������mo�f����V�K�"�򁴝��:�ۗ��Q�\7������������G�D"���%��
#���<�@C��J�W���8�;��Z�Q������	0�j��ѷǐ�g1Ƞ��О'v�U�۽�R�	��|�N��R �B�0������-�@$	s�� Ε0�-��x;R�<��}�y�@���I���Bi_�ҽ���CU�6�=��c^沼�0�<�+T�J�
1�˨,@��E�����ڐˣ��_o1��N�QV1R$m�if�D�Y)	A}w%�¨�B�R����BԽ��SU��F9΁JrGJ���W/q�ՒP[yXLn�D�$V��9XN�f�'�}@�^�p<S<C���PA����t�?ǂ�8��H���~��l�F��au�=ޒ��$g`d��wjVs����ۚ��`��	0ё�(�S+_S�a�|JӾn#읮+3q������%�IQp�-�����Wv]��XH�g8���>e�d;:��������n��ٻ�2����H�տ��+�9*�i=@��k>�Uie���S)
��@Lz�5]L^��̎�1�+Q��A�����y	=v_�q���O�V�=��4`��f�Ə��8��p���`>�)z�y�Y����neM!�t�Q����ʹ�g��6�m1�'�8�*;ܷ�C��zW���wf��uE�U���P��Y�U�W�2��i�8�B�+*� �l���kG�᪋:�L�%K&r���yF�rF�DDP4!���g. ��i��0iڀ��"I<��Uͫ�r$����!������ij�B�,2gm�; �gn{*@]me֋T�K��ݨ@[6O�7����@�5,�p���.-�+Z�8-;+���[�-��0���pS+F��<����u>dQ��l�3���W��MX�7jn��0���5~ᯄb$���)��?4W%����-�~W,Eɮ��d
3������<Z�7�U���\B� ��@hWr��:F��Z��ЇbE,�[	G-����N���S�}Ό��H��@b�[�!�\`��L$!�	�s2��iwﳘm�[8D�.����-gK�ll�Cb�d���ץ �x�Nՠ�y����Z�Z����X��/w���1�s~,��щ�Ŧks�h��L����T�!?{T���/�e���#[�o����e�F��җ�E*ƫAN#�errgI��R���æ�v՟��<=�#���5A�8�P��FVo�<. ��|��Q��''(����-���P���s��OBM�����>����Z�z�gnN�ǖQ��W9��#�:y�^~9���KD��	��1�|*�v��w������f�Ԁ���v�.�K�ΓO�?���� �Xei�=jf8?��/ a��e8�G�3�GiM?a��.�ta B� _?O�Py���:[������ᥬ-�yH�@�V���e���~�Mа2�O�