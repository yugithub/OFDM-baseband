��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��R��g�p3����Apǜ��p�~��!�XZ�1 ��z��Ey5KT�Y�T�cy�ϸn�:�|�4P�G0j�����0�H��
a˄z9��Ә��ZW8�|�C�F�`�'�/	��;��)E�)h�h��L�ߦK��j-��9*��	0��d	�����*=���ic�����<�R��=�ec ��X��=�*lZS�-�����̜��M�J?~^��w4�N��T����Z�

x..s���"m������;�wx�'��b�������>6$!�O6�1bs��4C��>����c�Y�<����QX�B�6xة��b�m�p�ЧƘ���Ѻ}{��8
�s���Nq��&�00��"Z��p?9o�ξ!������f��ż^9����^�j-ί���o9*�bU'	>[ضSb���U��s�z�Q�"�f����f�%�in2Gy�Ci�=�6�4B�e��O?
l��C��i/}:���-��l���@��&�u�S�;�� \�-_�RھK�7Dm�ض�ρ�u�D;���O�Y�,���@9�	g�x��?=_p�bK��l��e�C �졼F��]��ϰ����]�5C��Iӯ���eՉ�*pk�ʨIP��6�(����5ot�i�[�8
Q6C4;p�-dK�͐���6z�{�^|z �h=?Ue������mY����Q�Lf�]�>�!O�8�7��� _�*?g�s�f���7�y���N�3=` �#G��z�l<�s�$!�yX �r�p��#��̭/�yW��!�}� r׭��D����!�CE�ۆF���_��\�ןy�2���=��]��Ê�����R �M���Şk�����A���=}�KgQ�^^A`�l���=��#�ǥ�hкd"�0B��C��+�څh]C���91Twg�c@�.� ��u#����Թ�C���`�����*m����=V��|�=��a��F��3 y���7�v����.�`_Mȟb��I9��
'�n��	1^��xC�-�~�����W; >f��� (sͭ��5��th|���!҄�����5B��l�(�h�2��p�=�?m�g�Eڮ�4W���v[�ol:�1��Z'�v�.z�T��������
t	0m|~�D~PG��h�C�e&wQ��LLREbL����E�4�R�n����q�Pwu�N �A�jjCg,Tm<M!w��3�cA��n���9�XA�]�L �a9I���e�f �q���p�x=w��/e�`��/U+�&����[�Q|_{�d��S�·��t<1��g7�W.�x�=���W)�St�d֜���~I'��tr_T���Y�%3�C�CX�m`�d�h�!X|�M!ԡ�t5���)sԂE�B�!.w�[0�f�7��K�������B�+{���P0�TWX����� b�|ب�>�T��7s��*������	F�}P�b_Qa�'[w䗢@�sU���
rq
>MW�����w�^���w1��8��5�`av���M8d�����1�(}�!đ��p�0��&'X�n��{��P�B��͟����N(�l�;��Х����6��uV��٫��6[��kE��0c���Ǝ�Q�&� Y��]�BڅB�Β�A�=�B�μM�h�3�F|~�.��I��������Z;�t�cK�ѡD��i���Ul=W��4��f�l���8{;NլĢ�鬰�~��&�ŵk�����<�B/�����zu�O�g�@+u6��r��3}���ԣ\��tK��!�=�3IT��ҍ0����0�;_j!��Hp!������k�t x�A���m����۵�e.q?>�?�.$J�V۹��В�f�f9�;��]|�Ce[��.]q33���1):)��͇����V�9j8�� �BgTi�FB��H�z�
�"�gI���T��t�Ҋ0��R{������6C��<�)&���n@�q��ZP�Ü��1�Ư^p��K���T�[<�Ŷv{h!
P�A�綶���*���zTʒ����KW��@ev(J�b#���4r��_l�#!M�e�����3�Z/��e'��"	IX���W���*
ͅ�0T���;�L�M�jy���1�ƣ��"�sF�z�����[����i�xQ���v~`�Ÿ`q�3xܸ�,
�j�w�۞s�,~���u�5u�Z+^��fa&V��ػ�+��&a�Ƿ��W����t6o����m5�Ca�����1�02)*P���O
�^�jΔ5���&����K��l��z��*C��P�6�d�&
�B=�2L(g%�a��[���V����Vw�,�*T�W̪�۫�	��v)V1.���xd0WvYp�>/e�~�,�]�|1`\�<Gx���� ��kC,�eH)��M%�ϲ�[�>��f4J�]۾��s���R�r�Nn���p&.��&��Εh0עl�p�,���0��N2��l7�p@|J�j���Krۨa��f�_��Gs�c�����CNJa��$���4���؜W��8#@��Q�G�H�1�� ͷh�*��#��"��G���K��c3*��W �F[��X�K��xd�?��S�A-3�q����$s(���C��/�9쬊�����Eݯ �p����Eȇv�<9 �ă���ή�Yo�)Ow�:��=�=�yy����ŭù��܉˺n���J���*���Ƣj�p�m0��|T8�S� .�g�ʟ\7��5x�4JxqC��ER�{��J=G��������w��ɨX�vQxwj������`�\��2���6�~k�	"��Ÿ�(� ���o�F�	�в��T�F�����3n��yT��w�Y���qʐ9o��d78�3�J�㢛�rjxm��J��-�W�(����f�Nu9�U�~h�܏��	����<_Ϧ�K��J,W��HkN��
m?���� ��]�1��x���U/MtF|Ν�B��W(R2�@
X��y}�E��	7C�;t5�9�H���1�X��,�i�]��� ET�	/�R,~�>�S���+`�������ts����,|z�f�_�p��7�BD����k�$��`~��t�n,}�Y\�����Sv#�R=��ɹ��^Y1`�8��(�4���N�%W��|��dn ��S�Xs �"����}Q�!JÄ4пȺ��Ge&G5�,n�l�>U5���^ö�5<�Ho�����$���D�B�;�:4�m2V�`BC�6)�5�W>0H�*�	��8d���l�S�Hj	��Nyj��Ë�N�)��Z�ɐ�ƿ���a��ՠt8���(�*�T��U2�_�>[������c�a~�l�+w�Nk�G<s����3�"���Y!~j�4���F��q�f���"��#3�7UH�}�k�����;���[�#Is"�W|⼧�R�ĔK�oP���8EpD	�?����g'Q�mM;��p:F@>�Y�O�z��Be/�����+-�9��@��0�}���[+u'��
&j�k�c�V"��r�A,K�+����� �wj�mɴC-�&��j<1�Dɠ6Xyd?� 8yJ|&��A��W@��i6�9�].Z��>�.���7��tG�"��(<~�c*7-nvA������ 0,�w㙷>D�S氤�1�t0=���}j,��=���a�'�cvȔ��YaI��4���G�"*�C� 8	�;��Xŝ8Gq]?Ŧ��Rj��=�X�Wr��_�{%�Tȿ�-���`��ז</B��K�o'TT(��e�ob]��*gxo��`��,��^DRBg�nFC	��]%��k#SdaZS��Q;�@H��w��c��@����hOʆd�|C��D����6o�
w��4���!��s��X��X)ν6/$%\��D	�(y/F{:7C:�@�r�"�^�ų,�5�B;��|�w��x���G��o�G����
��av���KZ�����n�}�x�<ω�R���ƶ�yl�{�I7"�O�B5�ǳt�(lq��ST�B�rJRp̓�m�TwC/6wEQg�M�xԿ�X�N=-%@�b�,�+FE��T��	4��z� ����,���cюj{����Z���f���sϯ/x�а�hDUǰ�- #P��ͬ�4�%�S����3�6�D�e�.x��&0���{r{^�x�K����Qd��)8��m��Y5�����>���`���߀Z�5 ���iD�?�ȶ�}W��x�1����+H��`��,�,��w�*��2���)�Ʒ�p�S�z�`ri�y�vlI(rm�?=p'���w��!�*�-�8���V��N��Ÿfy��q��<��~�Y��*6]vӖ�nK��U-�����\4���o!s
<�%��?a��3c�i�gb��u�qQbM��᳘n���ˊp�c�HU�TI�l=
��2�%$I�X)�T�����+{�6��\�q��hOT]�w.��)����H?�N�27�cճ�.7��Юd��Ѳ���!�#�~�ꃉ�r����)��$�_pCl�׏` (C�J�lQa�y��f��UO�i{���sb��҇w&�wn��2薈�4�Á�O�-���,x��o���V���\�z��ҝ��Yp�:^��?+���Wl�[��*e�\%k�:�&��Y'dŏ����u4�ؚ��b��8�,�ܙ���{�H�'޸q�@��4��/7~����T�6)!��]�����6���'M�;+6���������7�L���[A(�CV�mܣ��T�5-I$5b6E�4E��scu����הz��<;'�Ш׿����PB�@�'m��ʌ���ѩ�ƺ�^���=k�+.m�iC��f��̥�ċ��ٖd����p�h��11��݇\V�AC��5���.��$�yw�m'+��eY~Ƽu�yA��`��b��4����q��N����r�ַt�k��%����%g;O�І=��e�Y���.p��;�XrM�u�����F)����7<NG���>�����RX���S?nC֫� �4.���:�bZ�N�0/g����r��ig9�S��{�AY�Y�<���3k:,_���b�ngD��9:����