��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6�����F��D��=�*�?N�������JV2�?	�Ʀ� �Bh��S�}Hes�)�r�?�B{�󳀓\b1��N�8���{�X)E� 5 -����@�{�e���0�t����8.����[���2�X�KĄ6�˫5��@�>b(I��+� �1��VV��~Z"	?�R&- ��A��嵗�Y���c���������r���D���d����nC1vg�m�4�عjM���h/yb�|�l�iۋ����	���wd�C���i����]!#��4�h4��Y��Y�@��nB�yT{7�	��8�g���p����y����9h.,�����`�k�(���ݔ�y��=�E�yƱ�!"^Gv�W��X�bY������qS��C�G@/���F�S-x�.pR����������O�č��X>������X��(���YN@Z$`�G�gqA����!�D	��� ��^�����4�s�{O�n%��A��5og� �j9�i�U�F��%F>�s�������e�Nk����n�74�O��$�����.oZG�&���U�����YA��]R����ת>��2�%Y����$�$O��cۺ�����d�,��'�Ad��g3q�߹A$�n�N�D&=�#�2��y����V%�����`�g���'�':�-)��D��X�`�3%*��+�xF�� V%�#I�+�FHcʈѐ_�ƪqʕ��t�&�mr~% ��(��T��q�,*A%��UǨyz�Bh�F�N�ğ���u���Yb>��ap���[��鬃
�T^T���k�g�g1�[��NRȚ���c]�V������Î�@�V�ŝO���ҵ���C���0	�xv��@
��L_Z���ϺL�j^��w��%\T��Cn���4x��r"A 7�����5�}�C�7��!<�|z�VC�+����λ�~z�>��x��We���N���?��&J�ր��QV� �qϔ�E���lX2 wR�H�6!���,$��� �{,CP���/bƳ��m���pY��N����^�Щ&Dݠ�w���^�5Xr�d"ĝ_�������T0�'��� ����c\�`>����������[y�Xmz�f�A�'rY��B�8��O���M͙S�*����D��'ʹ#u��#k&�YRImZ�[~�Z�?4����g��h�`���[�RSo�������W�YP?X_�%BiT\�₟��?o~+	��T�ӿߠ�����Y$���!��+NA�'��k�1��7�xf�l�A.�D�؋��/��%W������_n��
�lh�xr]�z�E [.!�'"W89mC�K�zT����YoL��\}.��EQ�Ī=����Ɉ��-��@�6����ad�K�sG��t�^��pG�,P�02�m�GK�Qik�,���8d���r��͚Gϩ�¿-Y; e/M��0��;�w�m���!��P��,�i�m�C#�:���1��!ȇ]Y��zA����CS�u�knN�w<V���8�d.ζ�y.{��*p�$��h�A�aD�a���n�V�?�LT�~�5Pn:ɼW,qH.��֦=�t��b��0o�0إy�D�p#\D5W��`Q��>��pwe�0$�f
�+�w�!s5UP����+Қ�g�������'�0¯
|1��f,쨡�(�y��:���fp=����JQc�o�?�h��6OPl[A��s�Ev�'s?O��˼3@�43L��h��W��C7�h��>f��У|�L5��#�r�y��BL"�Yc�a��n�O�\Wu{8}�f�r��I���p��I?�S~4@uS���3=�9�J{G�\�v<
h�a�"���a�}�5Wǘ��$�^*� ��.|�!K�qB����V��+v��[gϱz�����UY4=9̺�Z������ ����t�y3��� ��\j|�wk�d39����C��y�+(������݆=�R�	�_I���uf2��Ie�3K��0d�VC�_n��[�4�땼������E'�Rrz�O�6�[`�;���~| �:j�<��uג(�V����qo(r�7ԑ>od/�9k��sq�H�b(3:<a(H�-�*�دs&3�9H�%�T�m��Z�c��r�W+/o.fisg�f/�U2e��c�P9r��:`�2ؘ��)kӅ,���x�ڀ�ү��-�hgU�w%�s��Sy�dj!�'g��������2S�I8�)9���\o0�l���>�',�C�r�3t�:1%� �pK�_t/}Ǳ���i|l�����F��0~��qwA7�>Dj��$A6�Dd���#�~)A�"��QT
��	~<`So8��=��t�q�����\����</|���n����m
�H��*���T%g���Y��J��l��x�`,w����
>�Y�ȅj��d^)P�(0����+_��Z�[�kT��>d����F�*S��|.)Gb�,U���{T�9IVm�Iͽ'���:�e<=��^�����bm�}��v�C�z�k^���I2@�0. � ӡ����p($���������S+�n�V����#�c��]��GXBe:I����YwC���Q�����9G�j������A��^������Ȅ۬Z>RL1*���F�0,�_q��R�G��4]�;����h謉�C�5=0 )��41�x�j
q�����f6E�g�/
ߝ[���ҟ%%��߈!z+K�]s��3�i��P��Ҡ{�r�R�, <����/b���hd�E�{�0����Xd�"�ݜ��5���3���}R�H�ڭht%�ɇ����<e�Z�{�?�$�ܪ���кA�-V�����H^�]S�z��xK�$Icڝ
A�P�%��*��v&�;��3ڀ�����*�So`�b(���* ��s�����ޣ�ٍ[H�Ƞl��ב*k�G"6�\{��*�(-5�dr]�k�[���9V���Z�A4�߬�ttFW&�������7T꟥SO��N��f�N���YHbVD�I�~q��+A�`���﫹=��u8J��Fo� Lq^[�B�Q	NYX�<��ŢUNI�b�A:�F��br;��`~�R�*�D?�fX��²��k�uaL�נ�\n��2���H�}䙷����F۔ ���XI�΋9PH�1��57{��b}�އQ9|�`�+y�G����U�%��{�rIqm�-����t�$gI ���r��*�5?������:r��kLG�j�X��������_l�/֪?X�*ǙX�ǡ��,� ����(H�\�p7:bD܆v��N"n�<��ȴs��J�}؏��Y�p�2���Ih�(�8.�3��g�ٙ;
��%Yg�E��Bı�G���,�i���C�i����<^�^k�lE��dtE-�g?O=_�w��$��;D�Ugmb�Ҁr}���'��a1Xo_�\��N��!�0G�m�0r~JȓOWPc��'�U���Q�F!��.�ĉ��f��O�r��*#ؼfd�yl��E�RH�Z��O�Y�#.0�MѦEum�%W�c�No����o�[��PO��na|֋�cTG}�	������[�R�ٷ��=�s��,vyD �볗�V�Ap#�o���+�Q�9�>p�#w�ŎIg��j����3��B���q��mrt�D�!��w����o�/D�U�h���P��?���M�x�L�]�����C�3�W0,�mU3c����AY��#�%"3��wlӞ����ՅVr�|�uWP�:9f �"�q~Y!M��(�M)74n	 �B	�.UԐ��Q�.#n`��@)*����}(jԋ�8Nۗ҃b�o�گ����82G*�����w����:Z��n3A�f��I���y������+xU9��-h��2���PseZ�Pk�1/2�-8@�4���R�~�G�ۈl��]������_1^0�Q0�OFLwN���alv򊷪�5Z�C�%�.��g�q��o�#�/F����i����������,pБ۸�	G"���(�xOc�*a��PTl^~���g�+=������T���cW���x+-�Qv�=�"=��I�+�	RHkL�QA(�B\y�*X� 0�0"h퉺\+�D]��/1�,��1���x����t����VPT��L^y-if�Q�$5��?([��h~n�ש�ԏ'wYÞ�'m\���Y�Ѱ�H�d"�or����=پ^l�Pߤ���a� �]x�5	Ѝ����y��M�yZ'8TǴ�31�`�
�,]@�|	�C�|/3�6z�dl3
+ŋ0Qg����2sj65��-'�}{�@��h?�#�d
��O���Ԣ�u?��D
��M�i8���a?62�(�l��`&>/HnɹQ� �qN������&aֽ�]��j?��y��So�\�@�$[X�\5�)&�(�l	k3��2$�����=nY�#/@�Vܻh'z�I�Q6�ǟ��MGWT��f�A����<C�U��6�[^Zat���>Y����2o)�#�s�$�̢�EU��L&R�О6k����රE� p���Fi�O���ߗXw~$5���l^k�ȉ��m#�f����eYӽ<�W������E���ܽ<;�
��b�'�Z�����,e�P\�������Z�Q��s~:�$��ض����8�s�D��B�P���N�����z�Y������Zּ��ғ?z:���Lz�����{�ץ�o�Z!��&�6�����*/��KI<7;;d��ά[7?Ø�w�}��l�o�!���JMʑ�c6��O�&&�]�W��8��gS��_:������[�Ǔ"�b�hzVbr�%�D@���������۲��jD���pe�T��tզN�(��ovQ�7h�%a-��BmV��,2��i8 o���k	����G�,�0W�p���3�A
�T`E�+�Z\���T����Lo��(��m�,y�Om~⌯c?�|�r�C �em��3C�����54��D�K�f���3�F�D�8;V V�V�)�-oJu81���NĒ��R�π��dТ;��� ���HLm�8-;DjǢ��ʥ'>�ʹ3Q\Tsʝ��F�TUV�K� �ߍ�6GA�ie����wş�;��wؒ�Ȕz�y֠���kL'������ "���r~�V6<�+tٮ�WMˬ;��!�4��6��LX�,��Q37&ݘ"�?�TY+�y/�Ħ��1�pT�z��l����<��$VF�����m�>�J���@�	�pu������z�ؠ�U�Fn
���|����{��E�pvBۻ�8�X���a{��)���ΰN�\{e[}O7�¦�s&�[��k�c��# Qp�e� �|9Z��bW���oM��~l��Cy��KJ΍"���B��5�6\���A!L�i���4_y�qnJj+��J[I|O�3�_k{��=Xx��I��O���w����P^Iu�3����k�1���hfK~;���颓�� �P�]c�LL�G��Z�E֯��o��bᔡm�8�	AŸ���Q6�S�X՚7�DKS�U���}}�U�ܬϝ�$0��u�?��y�>����c��O,~k����6�
u�Q��	%x�|-}��){#z�aX��y!8?��K�p���"���y|��1����gp��B�O]a�W	E7��MU�C�_�>�>uu�z�;	s9 Γ��� �7�wU���V޷e��[�pF8������zFA| Y��+䫽FlS3�hUN�U��ܬ��j���e�baCP9/���@z����C���?��2�\�Gf{�>�g"=M�lP;[��aG�B�qy���� �z�!$__E�M�iGB�z7��r�+ݘ�M=���J�&���=-���M)�n���d��pv��p; ���4�Ц,s���`7�R�VP�oOR���[݄կs�W!��Y�Ov��"��S�b�r�5�,b��.��P5���:���8���oZ���V�e��+�E?��,��F�(yO���M��D�'��e׎��hj�E��֜����*S���r6�����h4&��|��f2U�<N�oGQ��ˡ+&Ҙm����ڽ_����(��#����:�G���L��$��h3��I���˸��	\��%&�l٘�B��>�L�T�K0��9,W��<��v"Q1��b�d)�-��`"[�'tvu�(q����������1=�)/�����s��>m�3�	V���*e�Y����S�L!��
��<A�Sz�2|��2�0�W�P!��-��C/�c��l���׏>��ŀ�-�M_i����M���>ͫ�S{�c����X ���$��܅��@�^��՗���1�(���W��D��lvz�,X��ԝ.����}V�&s4ʝ���%o��a �H��Gx��BFP�� 0 �@r�b�	�lQJ�t�;z"���T#�.��՛;K)���7���2����T�G��K�x�'�#7	�f�4���3J_rw�	�����4m�����H#�M��kMs��T�q@��O�6jG6c�>!њ�1��q���i����㕙n�IK�����1�__���
k�s�B��TK��=n!6Rv(�?�S���v|� ���gl��psI�噥� ��b5���4M�c�̜`IJ�3�7	�TͫY�WI�2ژy�BH� .�]Y� ��l���7<V�b��B�H /�'k4lK�pD4@���]R�/���ǭ���Q�-�0��lz}��Β��5���Ƥ�q��q6z� �\+3���p�8q����l�"@�TALeN3A9�A��vNGu��i����l)��f�x���T�Ew������ϖ���sx)u�D"�&�Լ�܏�rC�8���Z0z|z�	_������M�N�(��3��D��#������6j���9k�jۙ0��(sqv���PD�.# �Ǣvn-֧���b�������_��ֲ�D��DK�:*� �����;��s���@������my��/���Pk���BO+��T
�S{�%_��;F�%?�_��)ky>tM)�?��x*��O|4�#6�V�{g��K>��	"{�������_�� [U�:�5�
�h��mt�Mc�!��5�i�;O�E�~�M��֟��̭����k&��WmG[|�SB�L��J�5�陚y�д6XO��~P�f�S���k;��/�;P�@����|�w@��|�%�&��]������ѻɨQ�\�����zΕ\Z٪'Uu�7��B�΂�z1�����t�C,��D!Z���\2�j)�9�暑XH=�!nџ�N���K͚�I��Ϭ[�)3�倍#ˋ���m�Ag�vfBS�Bi�o���D�|���+He1�����q˸0@�=x��<�*������)��GT;��8
�w�+�;�
���U�n�[��_W�r5u�� ��4�������d+r�%"�hTN��͙U�<����Q4ju����N@;,ќ&x�cR�ؠ���Z�a8[� zML�8d
�҄[&�p;�O�CF�No�v>�Jk}���v�F���Ҵ��a�Z`O{I;��	�UI�q��%؞��o�>���,W����i5v����8l�#ʗ_j����Z���i�
G|!�1V|�����:���0Z8Ɗe�&��Xj;F
f�wdbT�P+{�$�&QaE�z��X���r�/�W(U���9�m�T�6R��v��ݾ`�=�ԽJcb��3=�>��@�4�&��u��R�����~F�fsҩ���s�Z��3�jlNO.:�B��g�����u�9����'q��ON7}T
~��_s�K?�LWZ���^�S;㟍�0��?�"�|v��$(2�''���b��5�DFtΖ�{w�t�I�s0�ڋ�L�!$�d�� �T&$|]!�ҽ�5�Z�D�Gn]��Jh<�+QiE>U~�G��/x���ܮ8 P0�`�V"�
$f9e�᧣"K�B�ҏE��+�D��2Pb���L5�q��6�L�F�#jTH�%G�I���[O��"3�|l��V\MŘ̶����B�!"�ޒ��+�w���`����$=l��Rc�y�B�%]�l
�e�$��m�30�8|��j�k?�'��g��G�'�b�#����0;6�	v	o�y�UP`���c�L!�e���{9Z�a8�Ť�my]l|�^-�]w�G.N�@n�Q�6[O��<rUא���M�qpl������F���+��)�C�+E��K��"��?n�iW�<~�=�:�zڀƢ�mR�qz�KǓ�4�H�4����/,��+�1��<����>�"�6�ƴ�z��S�]U7��AE��#H#�=�]�V�@�'����n�w�ʷ��Z�z��h~}��[D)W�ܩ���H>2޻���.�Mh-Q���Rr�6�Y���xcj�Q ٿI�ْ"���Ӗ�q���4����&-�"�W�Wo�� ]��ڃY��5�N��A0ѯ�n�HrQJ�:@��Az7O�g�Ǌ��O2�{�
6����M�a������s �m�s�i����}E�9��'�&
�,�%�Z����Ґ�m���d�f�M�*&�������}�쥈}�D�a��J�l~�D���E�?�*҄�@�l�*���,��2c|��}>]�g�2,�:h��e�~$TJ� 
u�z��U�h�(�%�Ϋ0�?%��Q��Fzh[eb�u�>�y#c�'@�-YڂI��1lTS��M��l�V)+b���H��<�(���=~��Ԭ��փ<���4���� ������J"!w��&5�k���8�ÒDBRjM�)ǡ ���m3d��IiU�Zﰖ�s��=D��ɮ2	\ߩ/=W��*]YZ#�����$��}<���7/�&�du �L�0�~���l)p���	ya:]��ˮ8�ۂ����d���V�{�W����?��_C���C���$: iN�����}�lè|[�A���,F3T����5�ʁ�k���~mp�oY˰�}��;�{�x��R�:H������q��"`b!��SV�`���CB�R愭�g��*��Ih5�<u�fVՕ"�*FC�Z�*�k�-`Úe~Ѹ3��Ⱍ[�-�f�fE�ˉ�3���I��{㳳m�־���,��BX�X�!^A��������fX������+�p����ڋ_*D�i�^H�om��3|��:ݖ��]��g/�I4o���Ԯ�d�âƝƞMz�A�1�p����J+��Ī ٲ��Ik�)�叩| �90���Q�A�k�~B����D�-��#�h��s�눋*@��sH���י�AFn��l_�2Wn�kZEI���-��uvU;%[���o ��n���=�~�r��]R��ٿ$� ��[���	�K�1aJ�k\'I%}�Nu��V/@�A�Q��%pׯ���MS�q�
<۠��T0��
%;�K��##�ڇ�I�Y6�(�`"���T�Z42�޾	��[Z2��]���}��#�t�D@[U�[zyٝ�M\����k��eA��۵�/��5��3(��Ilc�L9	�&�^��4fFZ���yqpbBo���P�܋�LMv0	>݅&���Ht��a�A�ɇ�����29�jFp���L�Y�\²9�� Z?q.��Z.a>Yk�%]]�(��܊'>��PH�����1�Ν�-+���o�p�TѬ�&�Q?��.��ѵ����#��ˁ|Sǌ���HYm�a����|���)&}���"��^�~��T����xv�F���GR�H9|yS`4p�`i9sh<�U��.h
�y=��wj��{��b�t�[W�F��@F��[Օ5(;��cօ[J��AD:�ێ܆5g�	�O@�p��s�)-~e�2R
�YJ�Wn�_Ǯ~���d2�{�.���íL|	�7��p�J������1��磠�n
fa�����ň]�":�}5��a��Z7x�z`�r&�o��۪��>.fuO��X�5Ĳ����VZ���F�A^l�n��L����kߌ�Dl���hQ9V�>���0|9a�ߐ���=�b�!�����$���������&<�SK7�rtQ����=,i��ˬ�'Z��qDb�cڏ�o�==�E4���\%KHy-�Ҁ�t(����|�vn���5���O�ӥQ�"o.�-�/'��i�@��\��GL�5T>o$ߩ�7��.;��:qŅ{�bD �#6��`G������AG��,W�U�I5!V[q�W�2�Ո�:���tx ��5���/�S� �����#�nL�_��6ٜ�}0FT
�E����d���`�/��?`���V7�\x�+֢ݘ�s|��� Yv��A�ڳ�����+��/��1�[ZR�4b:�/���s�H)!¬�+���O?�sM�/���o�X���籹��"^n�&G����sѮܿ�,V�[1�W�<s��n�?�:�*��f�$��h*� `�H[?��[� �lC�!7�l3D�@�e�E�,4��I�uaEq$��l�����xG�f$�a���.��`8b�MP
�`D�� ��_��@0��.L�-y���Ah��:�H�O���r�5sP��t��N�2�%F ~�t��҂$�9k�"M|J�}�-�۸g�]�z�5h�'־#k��5_z���)*�R����'Y2�m<��:Í�o���6�ϴ�he�m�ӤFj���;zw�y$���Y��V,�����I�{�����7�7"�ۄ���Y���v #�D�Xk�,�IZ�x�f1�k�/�p�k�1���yH@q�#ĕ�U���O��)62q��KN�CƟi)m��}́�)�-���d����ˌ)g|��d��߫=X,H����� �,�I�3���эb��C>�Gv�	Be��m~(�5
Z�l
2[�I,ɋ@���?\F��u"�Cj�r�=!F�km�.�������ծ���o[F��D�����D���gO���.��q{4���)&\���Z��.�$�A@���2�#�ȁ����,�K}-1iD|��M�S�!!VC���ٚ�&����e5"���z`��Y��_ŉ�}vhIy#�=��]�W�uB�+��&����4�co�vf�Lo-�l�F�yL��e%�{������M���g��ZeTTN���1��_��R��@O1AnC_ҷÍ�A1��2��5)3W!���Ķ�����홃��R"L�o�=�}�&Ƙ[���%`Pw��?6�,p��7�dė��l�h��ꇧ:��5;����eNx��W�H�����o�S��$��P���(����o��c#<Z�����I���i�.����!�6�mX��1���2�<���K�<<���ݩ��Z���v�&������{m��*����w�W� 
��V��J�io���y�L�o�/�~�߹[f�@�ei�ev#&�$U�K��P�'6�{�F�d$W��w|��8G��!�VI.���Ռ�'JT�����[�B�S�e~j/��M!"�rhpQ���R_(e�i"�����F�+��ϽyO�A��u�-W>��}���!GQx�3�e���ـi���;E̠��;H�n�߲�W�>��0��,/� �dg\�_Cr���Q˩�%�������E�8q��P�hQ�adOhj��x�8�'T��,�q�g�s�������H��jv���<p�������ٶNLj��l(����s���7�j���$yW��6��t�,u��$��e��B�@�9�=�������ތ�4����g��uwm>O��Z�i�`1���v����Jڅ��Uь����a�	��4�	�O��]�y�\1���>�:Қn����:�@�V�J��QK�9�P��L\9a�Zh2M����AX�	�5���#�3�Ќ��#U.U��y����K���ȝ�X<P܄�~��Ѭ<��.f�I5_�P��?���أ�A�tih�9Ra/Z�,/������q��-MEQ��umL�m�呎���G�ό� x�|�͚���b�Z��!E(F��}8o��`.��e1<��Wl���"!S������CJ:y`I9�g�P���t���[x��v�T#�8Ɉ�%M�tl)R��8L�����k �}Y�p�/�Ž�-�<	Vȷ�Q"�9b���]��$�'מGT�A��NP�@i�K���ӑ�:r<@B0�>�����,���V��-xLԏoՏEf�}e�\�XW��	s��;�����S�9fW�R�����M/�\l���H� �9���E[抒P��>Ex=xD � �vO�q�G�j�G�j&I{�F�	�!�z2�^Rsͻ=¶�\a��dvz�b �d7��?/�u�L-��D�Z�
�m9��H�c��[��!��*]U��9������RL��"��5���w&7$5�DF� Fp��K2*^'��`��Dt�T�C^8R8���\���§�x;N�r�HTƼ���;�|ƿ�ʡ�K��zs�D������mH1Q^�Qz��/�tp]����|U�Q�������Q�?y\X�)e����X庐]���.CaWZ-��ք�6���~��4�-5p��%�}��x[!��̳�\�8[0�Թ��������o�@����L����Q�}�Ӟ6G �t����jژE|���?ӎ�&��&�����q�{W1S<��LJ�#��.�_��P���o�vU��(�w��*i��E�DS�WX	�] Ε��X,��!�����Qq�A��j����{꾿4�V52i�=6�(�t�����f.1d[�Ĵ�d0�V)/�#]����@��m�$d�e�^�|���5��J	�ћY�آF�¹��4���Y�$i�H�)�K����Q+N{\�#�Z42�]��Id���:��T)�����6S��Wʫ��h�
��ǆ8�<�9+숹���#�L6$�'O.���«(�6H��W��L�!��Q�?�[t�`8��Yx��ul*E<˹#r�ۖD����<�A����kI��v!������}�ՓU^	�h�,r�5��u9@v�6�lk��&	Mކ��t@hߎg7�X^D�^ :����M�����r+Q���[��'���@�s��`'���ż�.r����g�mv/ u=l����CG�}Xȣ,�"��˃�z|5d��kƺv��M��8��az9�z?7��EY5�â�޹<@ť�����ծ
�8"h�����|�{�w���F�/��	�qa&.t�C���52#�4ʎ����o=I��,��H��#>�CӦ����&�Q-�Kx-f����L��4�F�!8S0 �5(�D�=�?|$��i_�������i�:��u��xI�f~c�]&؆�O<�A��x%_Y��f�k9�:P�i0��1�`t,i��Fh���i��M��rMǥ�y]<q�~��G�����ˣZ�!q˟�?�Zv��c�����js�rw�������q�DVR_�U� ��w���ya����3R�M�f��i�k���sC�mh.��F��}���c8��ыQ��E���P�?M�>驿�V�zx=��z�j�� �r�JY/�U���2�m!�����m��V����3��%�(��tW����*����{od;2��Ƞw��Z����d��p�C�����������A��.��U�����؆�; Źr�y�"� �ƞ�G�?�}\l��+�L�-�z][�N�B	ԐĽ�x��_ǘ��AR���3l#X���l�����Ge&(�i�lk�)���}=B�e��q�S��c��r��&�K���@yf�܀����2P�b�O@7y
��/�ܖR�T~�n�1�
��N��2���M$	h��.��)�A�����o���1rT�`?�t���(�Te_+��FbfVcn����}��Vr:}3�QF
���3D��H�-��)J��dS�%���t�x	�D���YZ���;�[uZG��U���E^�>KPm0��M"�J�w���� w��K�8��$�xmSI��x��6,#��&�4㴼�z��h?�[�)��/���q���k����J�[��Na�\���6)���)z4�CB��g��Ju���cN㒚�#�ƛL�ִ]�w���w��"��I�V:��� eߜ4:�q��dv�8*��t�SK�IN7j�(OaZ�RR�a�M��[vI8���S����_���(5"��G2�"7��;�`hx{���o��I�����;0�Z1��C�����h��* ��ך��;���fq''X�a�e8?Ab�fkY�.��{P~���Vek73b9 �}�}3�COh�#����9-��{�KJ2��*c�c���w�k�X�x�N�?��O
�r��G�ņ���h�*����R���=1�B�Ed�<XWh񯔋���E"����!���4�����|oU1_3�[X)�V���Kwҳ#����.n}��G�q��ɈÙdݸ�=���Q$����b������w�V����>@e#�j�,0
g���E���p~E��]A<�_q9��n}M�����"�|ΰ$Ak��΍��B��6�.ے���Ã�tO�j[N����!���uk5p����u �!艄D����=լM[c�0�1���n���vs/�A���x�tj�H���1�y�]�����T���X47"�����7�r�����ˢS}B�Sa<5Ʉ�ݾi��N&�7�,��ϒcCw�4��h�.7ϱ��dq7~"g#W��rWWQF������«�ce� \ �bHH'̈�L��ؕ��Q|�b]�尗YRJ��u�ӻ�z;�צ����M���SO�?0������T�r�ON���� �&dg#D�%�?؇.<m�{�OhV��D�P����@.�7��z�N�\���	��΅f>4_�-3]��}�Wj?��Cd�b�����b�C9`աNb9A�\�^,���.uB���ǹ��Jؽn\�7	t^c�0�<Z���3),
>��@ԧ��
)� ���8G�B����r]?L�)P��-���$�hHM�lkO&MV@�����.g��o��s�AY94đ���H#Uv���
�����`2 ;l`�|&��S1F��'�Is�v��a	M�n�*	�P��lb�,�d���;4Bw roV.b�4y/�t��s�
�ݷ�W�dq�#4�̀K�1vz�=IKm`�C �	�����9���Q������Њ�>���yC���>��g�6���0�����1��%.]�l%�蚑�SWd��4������\q�?@*���y��1?)wj�о��T�0�Ɂ� Bb̓���,�H����qY�)�TE�o�w����a��!�v�\��*F\ ���g���j�ݵ��U��g� w"d�~�ײug&��HI}����⽬���d����[����?����d0��F}��=Kt�rǧ+<��DM��8o�_e��H���Ɛ9>э�d�������m��9�����#�"�t�U5�d�y��I�QԖI^�ZdN��zN��쓦
��P�x�G�'4�=\������ �'^�;���
 p|�hw��p�r�B_�e5�e�����	%s��I��=��RpЅw�$L J(�
i�X���$auӕ��ں�����M�M ���x~p��D���w܂_[M�0 jeX�5h�2N��IQ�
s�6��5����� �&�����t��_���9�5�3:��QwZN�Uk������c4�M�!ۀ��8�T��lð�sSa�7���_�.$^�&>|/hU���~t�ɯ�Q8�N�⏜�R���X����� �/: �N��W��wi��h�Ȕ�(��V��Q�O��-﯋�I��m͋ں��L?L�Bb=�~ޤ^�b%b�� T�n&\qƌ/g�M���_a�v!���\s_HJ1NG�H_��ds]b�in��kjnB%x�,]����z�sR�.b2;�=}�M�j�Y����B��� �Z)x�S��ɶ��_�=�ϗO�;�� n��'���������4����o"V�E�D��ߋ�k��6����S�eH�W����,��wȳ��?D�׆�ÈC��)��n�&
���K���	̔!�{Q�N�*i뿉0j��=�v޸y�AY|���9�ٲ��k��%$Ĭt���o����)�����Ն �
�g�g�;���sL���f�P�Y-u���)&��9��F�y�!�3�.{�g�#�	�� ^���k���?c�q�$5��\)�5>�h�"�u���!�lY������)0T�ׂk�����7w��`C���{�Q����'��̣|������	C+P�Ȃ'im��&L��x���#	=��S��H�7�R]otq���Fxf��F���� �N�	�4%�^âmpʻ'�/�$��z]��R���(5GJ͍�w�:��,7�D ?�� P���_S`���u�O0�@����8"x��.?_n�����[���`�P*���	�Sh�43�bF��6/�l�c[�y��秿�tֻ1�GR�ӥp�H�Sy��&@\l�]a_h/��ʂJ����&�ͬ����~a;B�E��{�;�@vRcх+�[�?l�ƀyS��f�����e�'��k�Â�H;M�|w�M��Ió�I��6)���-A^��2D���E��9D W]R��n��=��+��>��>Z�\<%�j(դ$����\ۚ��@#�g���"Ձ�w{���Z��(�sk
ڗ������["������D�'��\�}Tl�*�1T�T�TB�=δzb=�	�87x�J���A����6�)M��6S0a^^I��%�u�/#�	q����pG�|��/��
OjiA��A/��&@��J@<�{�TM=���O�4x�Ge:��Vß=�a.l�	}�L `�})���@�u`�gn��G{����n�cB��ot�,�XĬӜӭ";c^�3u�����}��L�{�TT;�4���}ա����F����g���\�% P
��80U�N�m�f���f\�.�%D���J�n�G���a��V&}��.��%are��n����#��3�ۖ�\��yFۈh\xA�3�z3���ͽX4>�f~�<�;�L�ġks�Ƈk~H0�{����\������<Cн	w�&L�>��J¿��i]���Z��4'��sH�W��I;6�k;�)QSӤ�Is�Z��<~�ԗ���w�z��c|�x~#�� �1��?~�'?<�� ��;7�(��9[1�t�4"Z�n '�z��1>�� �V{��q���I�ؿ,���l��me�Ŭ�ݑ�.`V���"�`��ۜ ��C�˕
����~����sbh��@
!y~�)�������g
	f,��X.��$q!���[�+p�	Jڽ�Y�<yR�y���6P�󆄋ME�����3����x�zWW�Y�G��4Wm�p����E7O�&������'$R��'��;(�+R�Zr���Fj�=�6�q�SM��艪�>�N�9H.�B@ ���������:�G
���_�w=�^0��(��=B�M%��"�'�3��xڀI;��� oHR���C�+sW��h�[+�Ƕ4cR����9��"�a��]��k��_���eh�\����|�;�q�J1B����x�*��QfY���6��p;�/Y4U�U{��*���X9�+v_Y�����&�v&�V�L�r�2m�j�����X'nbi����A֑(�_}��Fy-�"�����ˆٖ�5��9�X��,������{�o����`��p8��t�=���"c�|iN.b::�p�����ຨ�äϗ��nEY6�-���-�^���J턮S;�G���E�ji$�` �s@�Ӊ��2.Y��~�l�6H �V*S�&&��\����V��I^�cLh?�Klݕm���DX@u��������K_RX�*Ѹ�������u���=�报Z��qYMH����=�����{�����pq��!9	8w�1�>��G���8�'w�gh�	�b����2�^���
�����_�W��L�}xOo_��G�m%�c�bz��/ ����o����hn�
���_�&�uی(T�~w(`�G���&��� ��00w��0Fh:�Ҩ�@�\%_K�q�C�x�:�{�5?�CPЇ/ML�pj�eO�~�ӻN?���+7�z�F3�`��S��:-�:�~J^s���BnQ~�uJ�g:�Ad ����0�y0٤<6���ƗC|.&��l���� ��n8���<H���T����ݽXj�Z����£��)a$��2�['�ܵ�bs�L�0&k?_*�.]$�ۋG�f�&�.{6Z��$�lU�;����p3x��୥��7c_�M#C]�9�*^S/jvW���Gߨ�jG��	$<����ew|q�ߞ����
8�<g��չ�S��-��b��8�mXZW	�O'B	���߂	��g8��O#���ӿ��v	l�8_��TjA�L>�5��-!���E�;Kl-b�1=}�)��nklY� ���_�FO�2>��N��	��g�iz�����B�����kR|;�k3���R��}��1-п�k�S$+[���X,%E��?~��3wِ>�Q��<����^�e[yXq�>�	���O`"X���ڦC��&5ZH�����U醧����\�\��2�e|�aT������G8@I�m�&�����#��L��������"C�c��7������`[�>�Pib�n�=�MC��4@��N8X�8�m�0�;�9����2.9;�"C��6��SLO���db��v����sH�}NB��ͯdv��,"��&FK�;����G��\5�&'�@
��r�A�J�o��]!�O�};��K�Q�7>��vo�>{�����1Ni�g���H�yrZ"\�p��,
x��`@;驫���H�������4h���v%|�.� j����������'�͒� �W�6�&N�V��w�bS���� �@VN�@'qS�Ys�����Ц��-�܋ށnJ��M�"�.�Y\���<Z*�ǋ���\:h�Z�7{�k���'tG���(�y� .ꏛ1`���iL�+6��W��@C]������� ����5�z�2)�\ٸ]zb��ڸ;�E�X���}]� ��+�y�`n�Bi?^�x�$�^�3�a�G=��S1����`kt�T��/s�)7�����$߾QyL_:2�x�����j�	��4��OS�{U���O�u$,PF�9�Pݧg�qZ�
��O&���_���J;<�o�� �7��r��¯�>��g|q#�hq��gk���2�d�/��ጿ�fy�
�5a:9�6�_��7e��r��BzZ(ӊb��Xޑ�L|B��X*J�I��y��
oRt-���#ǙI������3��� U�U�f���7&�ykȒ;Ŧ�o_>�x<(��}T?��k�"�l���Z�y���Q$9?*J'J2ϼx61�xء���W��*�2�9ˊ9�I�!�! �L��n f�'/�"��N�/���/kb�Ҧ��+��M�ۤ	*(^&qW�z��ǰ��ِ��A���g'DT}����3��6x��«og qc�ǟu��dѪ؉/J�-��`?�U���:�˭�EKC4Y�UvCF?��qk�B�$�����j*�嗮(�� �bj��ė�����/�$E>z����{����ʥ)ѓ���D���ek20̌�ڃ+��ێ�C�Y3�Z<F��B���c�[7�R!�bHuRd��@�X+�y�#E�N��4�y�`5ڟ�b6�h2b��Ш�hjk^S��ʎ ��{F:�Ցĸ�7��� $��]�y:��YLI��5�_��Y��W�bhjȬk!�{�G\@�	S�R��%܆,˫E&ߡm�J���L�}8>u�\�I9gOP0[�c4�&Q��=q%�����J��Vs �J�"�V���.����`��W��^m��zuB&��l�P}f��7?%>�|Ĝ�;�����tn�h��;eG$�/92B�������,�����[g��(��`x�lba���sՑ%���F�ξ��k)ץ��b+�a�c����
-
�K]ˤ�#ĝ\ۂ;�K� �� �����f��[�uʯ;�c�i2�#�u'���h�t��ݜ�L��o>\�y�����l����6#�\��2np/���r>�� J��	�̹:�J,��U3��#���\#d��'����3�P@n��ns�s$��o|�rYQ�;�a"��Q@���Y�m�\�
(��;%k��!����\3J��_ڬ�c��i:�-F�m�2�$�N�ۿ�8bb��ߓo:�yzq�y�0K�l��٘�,�]Ng��nP�m
���5gc�ɾf�5���Da0u1��,1��o9�N�k����l�3i�M��.��t>����U#\#\�i���Z�sE�J�v�:f1f��s�m� �T�󔊖��J�>�|oD�>�C�LJ|��x��+�"�jF��z�'�*L���7��A3M�u��m�~/�;��扣�E����P���Wx�=E����3)����5h��/0�9�B��#}H9U�OG�
��:�ov�(%-e�`+n&m��]3�S9�M����ӐL�Ⱦ�`�L�t�O=ƪiw�Y�ǌ[��7�H��[�l=PI�*2&�������TȚzF4�!++,`�W�T�(����H��vihT�W�Hm���S=V@y>�jVH(��.@���oc�w�8�9�pw�.�j�&,8!�̆� �?8��C�g�@'�{$FB�d	�L��rwgȜ9�J4ys��nC���l���(����R�I�l ��z���"��V��7q�Y���.�� ��1���W�]*LW�7�+V��^�P�XT��D�]�W+��ı���45u�Ŧ�x��TW&zgfw��%:3v�c�$<"Oyx)�
]$q����FT�VS��6~��8$�_cY��"�[�'���g�_'f��{@j+	a���d�L��ߌ�ڸ��/��a jȩ(�0Z���71Թ�N�u����������t�M����D��V����!ՇK}�6K��$:�W�6�$�4P� >}��@�_O�x��lG�1�qC�ݞ�W�Z�r�Ҡ{D:F\_��z��,��X|�Mn�J�3#-��(�>�c?�s.nd�>��rK '��C��-fF��ݳ�:�+�y��g;ve�އT�M�ڣ�S�33��)��!�;�F����Tb��T@����-����񤝋��y3[�CAo��jtw�3��g�������E�'��i�"]�I��r%�>f�Kd�>�yƏ�d�b$fza���֪00����d���n"��l���x��x�N��6F��@��7��$���ѝ�+����ǌ�&Խ��L�k�Il���P,:uV&��Ү���i��ѡ��L�I��1�}�S�67�`&�w��o{��s�5hNg[��J�0����ȫ����\
\Kd:yՀDO��q�0��x�9�נo)~�ҖSf:6lDgN�<DT�������r�S���&�ѓ�Z���1vR��C��������M8���Oɼ���T��R~Q$w�cl���������}#��%�P�����wU�3���\Yc�K�9oMS�f8H���Ϳ������}�Ģ�s�>�3C]�����O|6�g�_2kE3qt ��$����g�	g������1�(�͋r����[t���_T'#���E�XwƢ@����-0�O��R՟;֦<GW���9���fɺlv[�" ��E�?���~�A1E�f���}Q��`!c�_���@x!�:��҂DnHשZ��,�ϱuCh��vEŊ�����Q���'���]�?�;��Ps;e�q�+��K�J�;��-�m?DƧU}mt�;#�����3���R�Ը�j|%:�Ӌo{�:�8���ۦ�^l�C�f84)�F
��x���a(�~)lu;��� ��?�p�o�K���G�*��Tau����.+
�D���ס�8�g/�$�%�'ډaN3��n���X�t�R"&mw�gZ��`i�FS���Г9��21aF��a����C�����D�/W����b��)�A�',���F�}����|�(}��4����K&;�[��j�
��m�ԑ`�z��;�����෋e]�ڮ@F
��r��,O�H��������$�r��@��5Q�"���.��d��DH���+��������Txʜ-T8�p�͘�&:-m�X�K�c�Kv7R�٣1����ښ����EuO5���oX��x��_WC�~&c���&�i,FJ��X���:;U��z0���I?������Q���6<�u����h6��d7�Aa�����6�E�6��P�� �(��)��}���8�o�4��f^��hE=�����픯P?�:�O=?�V������W�Ӽ����[[C�T��6������ha��~p�����3���5 �sԒ�0�?�y"Ѷ�T�~K�g����u>7W�8������Y�/{�r��Q�����`±��j����D�ܚ�h���R:�3�y���`'��sM�F�x�	�����s��@��z�$.N�{>�;}��	cX?�ۍuv@�H���O�a
�D�U1��-�ʒ�v����c�K�S��@1?d�_��"ʏ�.z �ő�#�X65x,#+����"��t������gD����*e,�1�:���	Ҳvx?���q�s�@�쨦sW� 2D��c�yY/x�Vq<�|啁eV=���O`SU���;�}Uc��bzĿAm��i��]���CF\bF�d�E�ͬE��\���������Z�8	J߯�� ��2R]�RP��@�F���d����fXתP�b>��e �sXv�	Z^{��	h�!�/s�����M.X�� �Y�Π{Zr���i(��*rG�����ʳ�k�y��1��|y�w/�RaT�7�K���;�/��B��u�x_@@ͧ��w��Е��'���z��;�p�^��T	��XwL�M�^D�,�v����w��ٚh��Xc��������D>D�>�}��k�>!0�#��nu�RC��֤�� ���{�m����_�wl�]�9�r"I�EH���@"�P���85�41Gx�����8��rê.$e�ê��������#��0Ym�2z�� �>�}��WZ����bv��@��(���#"ת�v�ǃ��I5c�qJܾ����~�Z�jr��~�(H^��;�*S*�5��S�@S���<���b{І;��.N?��A��*Kd�����#��0.$
?����g��X���{j�W�~	���a�[��n�,�S�.��R*x���`��u��v۹�7���]O�W�_A�d0(mU5���
D�����T7w�/t����ZcJx��p?C"��4�-���t(p�Q����P��*�G����+�x:8�Hږ���/���V���,)�`�e��sn+!' 5uѣ�d��K.l�?hV��,y.��G�K�
{�I-r�4Z�� :J`<RC4b[餦�j������B:��y�]0���q�":�#�������K��=B̛"?B���[��4_xB޵��Q�w�Zm���Y�����8@d����r�`~g�_[6;\}W��O9�*z�,�-���L�J��-��-~�Y%=����n%G�e�},i���P�3g�=<�Q�F
�j��hm>�{�Dz25��>�?��ٲ72�ʲN�H��S�l��
�K����J>k�$�px�ꘞv�������Ǳ	dy6:�|��T޸�j��=(>7n����!�i����M$n��ӟ'go������%҉����s:�s�Z����.մ�a%M�����-�0��,2�����X�;�􍔢VJcj#�X�Q�[�Z���I�0*�S��a����{VƗ��#�`b鮧p�i�&$ڠ|3���_*?1���}�I�z+��� �_�|5ʇC�QWA��W�Y§���@̃위m���*�s��
J'�K�<r$L~7C]o{�M�D%O�ys��W��:�n�,&��*07�#��?��uJO���-^!��S��-�K��W�(��� ���[Z�d��j)��v��0���#��#J��	�3�αg��K>�ec&v��F���a	���L>��X�{����q��yz�I#��s���f*����}Rk�2)�^�l��{�n5�@o�V�I�qe�e��������og[X�? ҥl�ه�%\@ �*���~Zs�T�C�] ��Pչ��f�Q��ʁz}�^O�'�ߓ�2X1�Ȭ�W��2��QfȖ`_oc����v����2���~���!h�v���ɔi��)�1�D��DS�xn��W�І��*j���ct��!}�&�����'��.����'7�We
�UB��Si�@'�H�'<�!0�fAJs�qp^�HiF�
1R~�(p��mӉ�n�V�7+�i2w�o�t7�0��\p�k�f>AW����S\s��a�ja�џ��Dۮ���֮�-����A�NJ��ϧ-�ϸ�؍'�v�<�\�*��K���q� �RZ��::�:;��򿙊p�B���6O�YTG't�U�Eߗ�>�Y�BG�ir:|J�Ƃ[AINĺ�TV�)ʣ�a���}(��p��ehS��c�Ab?�Kx�h�9��������1{W�(��YP�H�������b�*	o�S2/�M�3k��V7�����YC�kdI�-.�����H=N{W%����ʡ��A�կ[uЪiS]9����&�`#�m���ȁ)�,<��D�6T�^�z&<Y��2�	Mg�`>w^q��!�$�R���o��B��&K�����f8ʡ)�*��\�+��zzl���c�uC��{������7 t�	�Ϻ� 9i�O��ȗыj/݊��c%��n��;~�M�+�}��6��s'�h4�_���1s��  �p}<h����w�:�	HL��H�pJɀ�jK@y����ϣ#G������e2�n��>Rd�Q���X�@��N��umэ��y��f̣���1�rd^����6d�����7Ȇ�P�-L�?E!�M��"0���P����h$�((�WF�H�nڊ�ү�D�,�l��_����u��_%��4���6���Y��K}�#���8�^���S�A�n'�V&��U�-����ʭQ���N�H�X�:<Y���|n1.����"����!���d~U�j�~�2Ң�n���r��v�>�n( �Ǉ�hQ������1��Y����+�@,�����1���ۙi���_����,~�1��3��S`�a��QK��?_���*.��ƨ�(���*ۘ:��PfƤ�t�t�ؗ#w`���Z��܀��Z�T�ǚ��,j��K�JUݷ�w���*��u�{���
��@�x\;8�g��װ�������!�r+���!�6~��&��׹u������Y���'���ߺ�g�8K�����̈́�ՠ`��Ө��r�fJ!r�N'��=�V��r|�.Պh�_�a�cUE8^vbu"����ћm����J�8U�,@!q�I��l���	WW��O|w[��~i0T;�-�K��P�
%�K��<����@��Ap�:�sY;�Ĺ�bL9ch`�������@m;�t4����hz�c�~�s.��5����Ԅn�P��b�n�9�|�ȇj��859��ף�[��q�f��g��U`۩`�y�^���Jշt���A�:�ݾ����P�S&�v�ȶ��M��Љ浞���?�S��Rk����ILa3�UT�����V>�<p�`�"^ߔ��֓\[X|��v�ޝe����H�����V#�ӳ6lyϊy�Ѱ-Ӂv�U�|�	}�p���f�Xl��L��{����0����x��L%����7�IR�w/J���qjI��;���~�x��eg��atz���*8���݂1�O��,�EdEr{I�X�󙿖d��O���*�%�a)��\㲞}���j0�GVyr&t'�I�����\Um=�f��N*0l��W��[zo�:#��}�lo��H�}���S]�'�h����^
�p��[�)�1<�EB��gw?�l�_�
���/6�Ӳ��8$�h���#�����IlkW�k0[L�L�c���{��9�.�&�q]�q�$�*����FUs}��@����ٶ/-Ԉ��~y��V��%��U��D
FP?r�vV�\�� �d����k+�p;/0���n�ދ.���X.# �bTP��%��Z{��=r+k���<u�r��k��6�i��Ӿ�����&���o�)	j�Z�>���uM!�����:݈B㥷�G���Ͻ�w��ζ.��m �0Q��d�A�Z�ؖ��9m�ܐ"ہ3�(f������ْQ�AnP�;��6�وa˚3�$ ������}����u8�����oj�$����k <8ͯ���@.���+�=}���-�C�BB��鸉s��4��k�F�w=q�\�3S�о��\W,�O�O�R?��:A��T~!�]���P��ؿ��wR�&�P,��V����7��&�a^�,~k�4vሎ�?]�/��-��7.�������y}����-u���y�0��4�5`��I5/��,�֏��6H�S�>`��B6x��s���U���H�_v���Q��m��m#��wL~��-ha`�~
pv�l�y`���6���v��V{D�7�Øb4'gTh_�uV�`�u����[6��\�?��w;�؋�����Q�j���b9�$5�iER�B�۪�U��&S�(�r|7w���9n	��Y�0Ė�L���	!П�x2����{}2D@Iu����>ZTD�]��tK+�hp��ȋ���6'W��o�B/�Y�Ð�~�F>�c��+�a0x!�8�jӍ�w,)�	�6z���xժ�͓�e���a�p���q�x�~ț`x�W)_��3џ$��� ��&���r�����Km,Mw�r��n+R}���ϔ�uj�OB2f/��5ix��_f
>m9�2����#W���[�b9��������*�q<�	��1}/	(X�]jȿ�sq�~
@:�GOG�(�eł�ܓ?+(���߸ER5ð�;�5դ�E.�Y{)+ic&p��c̚p6��\W���Ղ'#���'�`|��t]p�]�ƘIu��f%���Ԩ_9\�|n�0@�s��|Q���Qyz'��s�B �A���� �BM��|4<	�Iԗ��7Wco�&Kԛ�r��s@{���M�� ��R�K����~3
�r;�ُ���晚!K��<j���Qw��[�II���ߧ��X�{-��(έ�C���קjw��{rZ-<�O}�M�w���ԃ��P�FwO��v���o�A�ނ�p+���{�1�;fu=[�8�W�ol{��֌�~g�|z�.n�|D�� K���rv["���9ο׹ �������Hz����R���Utz ٍ����1a�#C/U�-��q���l�Q(�q�X]`�`�7J*����Y�"[��'��y:��E&�����Gv�T:�qt_�lȦ�8:����ߟjId���.�� O�Q����9�a�L��g�_��4�Ě3Z����1��=�:��,��԰��&��T�+� ܋6�`
�/��CA�pR��X��O����� DH[26Pj��Hh�љI�?�N�c$μ�#��<C��z�̭�����z�L]t={�?rs�%q����{�|�qxm]�t�Ŋ��t���R  ��2>�#/��M\��	OZ.~YX�4��_R�P�����@G�ibR>���zL)n�'��4�.�Gd֘��N'�6qk7RU��\y0�L���=��\�5F;���Ҫ/�B�!�R9�~�C���TjͭW�C8��O�_a��Lk�]aQB��f��<��b��c!�U�T�����}��gi��R"'M|G5Q�#U�$�!�~����@�nR��>�>�� �kS�������:47*���l�r�/���`f����A�v�����\����Jm��=��rAI����K|P)������Έ�z�z,J�����!&لh�*�4г݋Ǽ���^e�w�o�^���V���e�Lﱃ�jD4n��}�Ѹؓ��S1��d��i4�y1D�W�kE�~�������܎��Nm�,���`nq<@nu�{��A�``lU�ϱZǂ��ru	�*@J,wf�&�E�/�I��/H�Јa���u=VN��3�+��X�af�&�{��I���e��T�N�=T@��Y�增��f��rC%=�y�҄�&ܤ�(6�=����8�!������WO�1I�l@���q��<x��Ԟ���k�����No���UM�2U����I=�MG|�Y!L����!{�}�,��
@w�Q�e����*6&{W3���4�L!�!�S��S�IA8z���
{�?�{��Ь�?wu�(ƗD��-�)�|�u�y�^���D|�m*��<A^��y�߿�42��ԥ7�T�Ag�n�"��X�˚��N��m�!�$q̀������Vg���e�OQ� �VzoS�sd4Ȋ��N7Vh0�ͣU�M� ]�
̟�;��D�ͫxވ|�rҗ�(�v$����3\��T��﹗��9G�����RLv�QRx����U�o�K٣L"�?�P)�5�RKm�䗝k/��a���  �u"�pg����{	�.�z%L`S'U���2�����V����2��}s�Y*b�_�Nһ�=�j%�W[n�C]�3��ddswW�������Ȗ��
r��Yep�ෘ����fu"O�{ȡ-#cI⇚��x��QZ �c{cx�&����r �s��E����h�	�1ث���m@*�p��-$�� �,^���?�����a�aE�{�+�ǹ�
f�#f�-�̰�6����ޮ45|P�D�/a�=���[�a��V'�8�ݰ�+�Υ��{'���v��$��<�WM�T�f��l'G�>��':�<6e��#����v`58�ݲ�%��!f6&��d!
2��b�7�3����IaY�x�G"�2{�5�� ��v(��5����՚���a��Cv_| {W�ڰY?��F��H�v�sbko�%��]}�Œ0lHŧp~ҧ�ُV�T�bx�����wc
�[��G5	��$�E�W�N �*�t�FC *����Q�������/��t(���&�w@�{��W`��]h iE� �� Q}��Oe�I�yxA��G��a��er�o�2(�����f~�^=X�^"�'��`�0�D���%sb��s�SlX-{4J:j��	*q<��5����q�lW�Y�U]�Ԫ	��̝Ң���v�7 #��L�-;��}�����1���������w*���|���1��Έ2�>��RN���!k蘩A����ǚ<S�a���g�A��|Z��Te���ae!ݼ�M����Q i�D��2<? �:P`�������g����$�㟉���~8��F���>�5�g��A+ԣ�J��B��mw�MO;���(�|T
�۔z%S��s��r�$z�#���u��4�xf�fL����利�)��3��5��8�9U1�R@�[�ߘ�!�a�v��<�zp=u�ay[? ��_��pt����<�^2A����}�x;'����j?����"*��'aa;D~!l�4
Dd[K�)	+c/�U�[<Ƞ7�H���R�T-�S���1�J[z~w�R*��}���Ӄ��0l��p��;^�f�<�߽jسp��YE��AD(��KD��M;�7��/�!��/kf?�M�4�}�ȵ8}���uGɟ�̼%KҠ��ؗ���P�sL��� K���������`�.��I(���pԅLVLs:��G��=��K��F��9�^Mþ���U��fΫ�قQa�D�'5��	+!�6C����Z��OJ���kA�цn��bB�X ��Х���^�c.K���V�/��	ן�.��I��o�����U�����}i���6V���V�c7,�o�͊�����p�w$�ħ�^N�Ϝ�� -ysQ:���ȅT�s�v"o"����J pt�K�6��_`��>s�߅�Д�2?4c�o����K���¨�3v�<%7�d�v |4®�b���#�3���4�jC ���u��M8�#��)2�i�D�H�Fu9��cC�I�c�A�o������ڊ�]ڬ��t����̴ܥDQr���)�R&a��4|&��Z�i1��"o�s�ύ�y���!�ģ��'��Q�+wX��M�~��SqDHL�5����}Kfu�ʰ��m�>�L�bL�Q�=��Vi�F02�F��@;��}�&V<���s�Ns���P���X��׌A����z~}�R�	�6��/��y�в�2u܅L��iQ#l%�걨W�!��wQS����D�6CZk����q�G�m��۱+	 50���ԊLI�f�6#�>^�P���SW�0���3r��"c^�Ji�",�u���.������!�����bI��v+R';�����`��#n�H�	��խ��@I�;7@�Hu��W�������}#p]$�+��g��W�S>ʗݽ��5���d�^��(q�Ԥɉ�"�'��z$�?��Ss �*X;��/��%�H�Xړ`�٧R6����M�ZK������q,l �ˬ�?�e>MQ�v��-�`S��b�?�����B?ۊkyS@˓�?^4�\g�<^ި�p���#;1�1q�Dr����#��yN�z�ֆSR�ȹHKr�^�O0�(�nN�X޿�
Wn�����DJ4��)7r���ヅ�YoO���c��XB[�/fB����n����	t�Z�2jD������%�=F��P_\�"���D_��,����*�h���֑�9>�.p��|��ߢn+�xΞ@��}` æ���"x�P��� e�P.���-��X?aX,Ή�E���F���aṆƣ�3�
��|Xl'�U�K�I>H���#w���r�9�~�7��n��3$P �?^������
�\�]���.4!*��g��y˨qB'9�4���AL~tg�\�i��<'�����:��'�T;�p_��e&~����G��Yħ@�ã���`]�Mp1���8i�b�(����n�RWB6�*X|k�uit ��S%
ID�o'��[��i��G�F��x$���f���H>�Jfՙ�]�)~�&�p�E���iI
��>��w[��^)�S-X<s��ʾ�=�lom�v]w��U�T�PФ`9�5���BX�%�b�G�u�������,U"�9�[8��	��F�������Ϩ��|�U��.+�cIeoӣo#��q&�St�b@ў�Pa��/z���'ķ��ӗ��i��n�1��ha�f�X���_�N�^��p�?���*�y�:b4�fs�6⤷���uZ�[$SK��!K�,�P�����t�J��`�x5+��~Sux�I��4m<�Y�5Y��6�������Ɠ������D�k�J�w������H��I���!Ɉ������9��G�#��]�T���x?N���Cy=�Ӱ�^�h�J��c�,Ff+�V� �F��B(5�%R�9��`��~�X��M��Y���R�fZ��z� %!�t�FW�@�7�c���R��U�� �(�NIP](!��jM�R_�Eh��)chtb�L�;��[+���|����:��8��1���Թ�ɳ��o�2�h�O�M�4&��+JB��F��yeP�v,�L�I��N��K�m�l�;�D�{��h�W���}��hZ�lĭe�R����9<���:�U����ɢ�YT�ke�LT��J��G~��է͹\�5���|݅��p��k��M�A��X���۴c������e쫰.M�FŮ熗�~��x��5�&o�_�	'*���2йs �Ub��e&��v�Ѧ���܎y헨,��฽�����Է�c��qݖx�
�7>����=$̨�!?�L���~�&�*�˔GJ����x�e�l�h�p�{��`�|J@ȑ4j����W�(Y>�UQ��Rj\�f�Hݝ|>��f���1�+�X/�����Nr[��� ��ŷ��)"�.+�PWF(C�V�l�i�H9���}��\�2�X�p�ߕ�=@�r�Ӈ-]cIx���4dR�cD����?B�.�´YH,̙N
%���#E�����}֣��RfE �۱K���F���e��S���n��I����n�}QP��u�#���+���ٵ6��?{�y	h��ev�bL��@��P�	Dǫ-���O�RS�ߺr���0��s��u������vj�J�����o+��3�0�/Wg�G�x`�U�_喡��