��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6-g�?)]1H+�歓;��+w�_Y�)-��dn�I��!)#,z{Q}͎��`����yFe�2et�&�����[����V*�����L#�8�ùe�1c֥��<D�޻/��cO;�|Q��aIk?*�j�ZЪ�S9{��ت�
�V��������@��ݥ7�''>���4�r�Δ��וO'�d����� ���$�d�ֶ��&,w�3-яb[��|f�� A��K��W�K��|��1����-I{9��E,�$��tۿ��f�}�;�k�K�ߪ�<�8L2���_(��^�d�����O�5mMþ��(�F�r�G�k��L\��H�\>UNJ���IM�����&�-4�|G�[kѰa�@�ЪW�IfۢN��u��?��q�	{-����mԥp ouǪ���C��Ҋ���)<�����r@����Q�Z�����4�SAT2��hEeMl���v��'9ܿ�dz� ���#Bh�o �5�f�b�cE�H}~3�ܳl����̣��m����߇�B��\�nJ�X�J���Y��<�hz�,d.�z�xz4x��GQ\I��U@=�41�Y���+�9�L@/�`��:�*�(��<��`����}�
&�����)��Z\��I9?R33�Ͷ���!��ۚ9n��2Y�Ld��H� �7�E�
��3�?A��~G�� ߾���7�8�q��z��
l��(�-��x��ٵ�cN�l����$O})�� (������2�9u�m˃(
 ��wЇ	~~��.2��;G��I/Y�z1X+��˩�k@������D~
��w=�a�����$Y ߆CD_��T~��/�����׹�2�[F�CMܖ���1b;��:�Y�a��,o�;6����b����pz\Xʼ��jsW)Yȝ�k���aHg/QOٸ�X2���!�3뼭M�����nqP��P���4p�(�j���*:���� �Kq5�x���H-��b�I	��� N#�昝(	e�ޖ�{ �1^�
�,�8{��<ڋf���	�C(SW�pb�cү"J�|��!��.����WGҩ��mN��(.��D�y�P	\	.�<s0���Y�1̲\�J��Y�x���j�7���;��:$���(d�;r����@���o�EFéI��#bݪt튥�ʀ�� �g4�B�ˆ�ϯ���\��^�Ѱ��Wbo��2-�z���tE�&��E�m޼�(�`�0B��Ս'�UQnǆYH"��?d����k��x���J��H�^�"��T�Dz����	��ٷ���K�r3�������y��H�!`��PB�[���:���UT_B�{PΌ����R�D@�����v�c��s��T*�_p����W?ږ���*�O�x-Do����D��\�.h�L�p�;9B��>�i.�A'��6�U1D����ʴjw�ҵ`���zi����G�� �Ƚ�Bu�,6G)�7�@��J����l�>|y��5o1�_��QX�LfaCHK>�.�d=k3�qGͯ���?�j��R]�.=u(���a����4��`�W
��辅����Fn�WJ"�sʓ�/q؜��V/�@l��?�M����A�cmGD~����S��p7G�v�(+s��P��8&A��T$���Ks�z�?}$}���B��w����3��!#�����g�f��C�9������و{1��Ǉ�$�8� ��+O���1��4( s�"Sȹ�r���w�8CB�E�[D?� �nا2�HǷ9g�9�鬂��QU�6�؝ǂ��� -K�N{l�x��k��tJJKny�c.p�e��ع���>�����@>����`� �$
���ۉ�_.�ۋ��54h����ǣ���	�O�m(��iB�鹫X���o�
	&�sA59F����V"Oeg����z|�����7	�]�w�I�Qޗ� ��Ш��-K^
���k�"{s`�̚e���@��%!@����:�ưчY?��wCݛU��x�K����m���޲�w!�f��h�����pLQ�_,��gwQ�x�C�:�hTqO��r��5�����ˁ���%̶���i�A5(Gb�;��^���D1��{���H�Ax�4�s��YP�|�s��#�����L��G�C�- g�!i(�r��jpJ/9���[�8�fæ��I�v]LX;��*�#W��^��aX���C���&��u�n�KƐ�I]Z��ݹx�H�*��j�'��_k|P��n��T4��;h̖� ���U�K�� YF��:t�P<PАEݤ���i8�jp��~�y^���h]%]k�tәg�]�2��-�f�*py
Q$�O�� ��z<`����Bn&Qr�qQ��^��%��@�/w�y��З���چ�_�-]dДXS���(�U������b �{��p�qxN�YZ�S��|�#-}*��d�5����%P��or���l�[��ږ]Y*}%vZ��}w����}��p���8����\Ĺ���z���,�����"q>2s�X�Ѓ�-L��;b�X^«gcA���H�8>��g��U�8;�
ӹ�K~|�k�IzH#�VJ!"�?�{һ��u��
jŒ��I�EȾ�(�&��50�>i��P��_$k��cY1����M��F>��� �����l�b��ִR�����K�f��Bچ>ђ��1#YثpH,�4��x��d�&��e]�7�ǌ��P�I�W�lkF:���Ӧi	�m�HxBj)���
�<��g��I5�V���=��������ֵ����~z�Jpɫ��A�����������d2��wB��j@���U��C�r�f K2�0S$�-��7U#�z�Kͦxv��~DZ��qөl|գ�"y�	���"q	���`�z�y|@�.��Qkڴ@�ˑ	��.�1 U*��,�)�k�̄�\�l�ٵ�b��!�5�8��v<_�k�
�7����M���7Ɍ`�dXV�,E���y�7���W1��{<���'����#�t��WZQC|i�o�S��Tas���0�B�a�\f,_ ��=�P�
trJ+�"�:��O�i�Frܩ�s�k�*4�Rz^ov�	�$N�ߐK �rC�	�so��_��Qv��=/�Fᤥ�z�FuW�zEG�k�9��
s�N'�3���檄�bz���*w�T-FL�D�1̋�R�n�o���$�H�&n�p� =��=;b�⪾L�ɾAXwk���L���4�*�76!5����(�X���>�%n�{�//���@��Od��_�sp��BT�;m��k���aI3J\�W�גo��ᖲ'�#č"��m.@!��� ���F�� kD�oQ�H�?4:-��Db�~��F�vI�Q����é�����n����,��{���,K5WBӎ[5ds�E��;#raႀ�M�k3�{����5)4�Va�Wh��揕���.����P��j5۸�M��S\>��0�_��ɟ��%�|� qp��p���z�.���0��M@
�i�+��պª�^4��7�\2���ܓ�[5+��`��/��#e�s����surqW���;E�m>AQ�X)�b��y���ݪ4g��ȴ�����4}>V�G���g��� #j��4�i��SP�}���@�f��+��p;�J����(<" �qi����}��D�g���z�i���Z�\	mCB~���K��Ao���h�X��
�HP֑���Th��``�e��_Of�;��zln�I�;++q4T�A~�鶔蹭*��s��\\Ɋ�
"Z�a�N.x�r(l��]V
����n���U�ʻd��}����۠Y����,��N�BV'D��G�trᲮ7(�jM�����4�� [�x��X�f�Z��,�HD?Ԋ��:�v�iB*����,�o�_��5
gB��y޶�<�h�:h��R�1Y�S�-��	_�Q�Y��L{X�#��Q ��?��XmC+S���}+m1�+oF�5_V8��t:b�f�H��w3l�{C��n�����eh������=��Hj�[L,�4�U�d��摪$� �dY����	�(#s6a
����\��8=��T�%P��ri�ɾ�3h:W';UoZ�_���F(�=����R{�嶰�7?�h*�	j	�5EZ��<L��\�`Vi��N�{��|XVI�'Q|�磵����[�U{y����!nE ���/&�75]�ܾ=�l�_�V�+��(�#{��DT�(�RN{uV�"�z�h� ��ہ�#~�dG��8R��oϵ��aM�{�˿��+I�"�9����"�.a8����O �=��Y��Q!��f�(�^�y�lBaB>'DEQ����N\��1+B�=!g�I(�KS6�E���c�� o��`���6��M�7�)��3iE�f�x����>�H'���E��<�\�� ?�̝*D?<�H*1����K�3�{9Is��
"�WcT���"9�	ւ�����%�T�a�FI�E?�gm�����H[��D?аE�����*�$!XJ�|&]
{t���$X�yut��>�?(�ȉ�ʍ��u�Z=�{��WR۞N_(�7N��q�,Zn�*-������y��\��	k \�
��$y�<�`�E���9�c��G��v�n���c2�3���	WΓm:q�B�'����`zTe�ܛ����r��X7J?�#�3�	��s�H�sOk!u3Hx= >��̹��X;�ű���;�bv����p=��!���-�4X��,�(Pa�a�$���J���اUt�bbh�>��f��堂h���eڏv�����
l�4��$��� �vm��W����IO4/��Eď�AD�X��� ��)����9����|H�*�5A�y~��h��U��CY^-��Ck��ٯ�u�����{gq���[��Q�H'� \��3�S���ZA/H��W�Qk�&�j@H�+��8�|�`*�c�ς�x�F"�}�X�gCG��6�c�	�T��^1:���*�9Z�E|�4��[K����N���gv�1)ei�3�������"@�]9���Ux%KbI�Qt\y��%{�B�'�S���yF����J���]ʿT��	KN��,v�MIn!ː������h�)G�C���{i+#��D�%UéG]��;��P^��f��yb(@(�,�q+
�|-�?V���B���~ߕ~�i޶Uh������+��r=�?��ET:`CxuͿ��Wa�ۊ�nӋ ؟������0j{О��{����9��m���v�&�N���m�����g�+��n��F�z��<͔������(;�<��~�E�#��8��b��z��8>J�=�%���"e_DE)���?;���i��V����%P��uϐ���R�3ޯ�ɺ�`��#`��$��,�`Z4�3�5��������q��t�:sǖ�Y�&���ݸ8���+�	��*�c�ݠ}�`�>�,&�]B�֟Qn��P��3���܋n�a�w�~�_�*�OEW�u�� $�D����!~���]�����D��~�D]�:�j@��,�6�ؽ9~�(���1���<ӄ�ʜ�v@xy��/]� 6a�5�u� �����yD�7����L�F��4`ˤQ���A�,3��Ϝ❤]ͧ��8M���V���'mDTt�0nS�3���ʷN�р�!y�ێלʈ�L�
�m��E�E]�ك�8_0�H
�-��1l�[����}$mxqy�ƨ�s�ϗ�y�j�d��nݒӶ�F>�h����<�<�Z1-u��J��^[��14 A����{���Ą]�)��h�Au�E��-j�]p>x��̵�LR7=��{�����t&b6�����0K=����?z��qѮ�Y�zy�\���Y��4) �r i�Ʀ�����*7
\C�"�������4���j���P�"b�� �i��ڧ ��'����p��*�zVVmӁ�ba�O�,eL�����,Ge���]1T���ζ>����h�FX��{B��\��֚0�N�"��>�O�e=����,i��+�c����?�tD��U#���(���=���G|�������⇐�'�w�}��qZ��kDA�-�� z���>�Ֆ%��>����9�"��<�~��08����Ϧ�b��x�p�)!�Յ��Bk8�P���~+�'�x�-{9q�� AD�;%�A�Y�B�㮼��{�dM�-P�K#���t�n�{G��"�lx��]�#O4����H9��<6�k/QM��B *ZPj@Eh,9Xxa���J'�<mad�KXf�qK�v�K�S��*�ͯM<���Kƣ���K}+((��-��RtY2]��K��/U x�Ş�ѠJᙽ!V�'�RD�qG �1s��*>%,�Z�fS)��vb�w�n߯���g�T"� ���5�&��������jʶ�{��5�h�4�:Q���	�L4 +��2p �� a�@�ӿ��^yEΠ�4r�ӗ�4z&�0��(ƪQ(L�� �;y$�x��L*\ඝ��ӱh���~'Q�@�O�y�SΛy��9N�;��7"�(�R�slۊ�uw�r��v�pm��=Ю����Ba���[����#��n��w�X�z���M�p�/!u7W���`#}g�:�/��J*T�Yk�Fbo���f���1�+P;I�e��x!���ඥDK�IqL <�@b�*����Y]1���վ~���
/��);k�c1����W�p��M�����	�J�c���_�3m�f�  !D$�E1�a_k��l��u��+��h��\�~��#p%�[�W4E�;!���1A�`gk�h?�̦��ga�F��U/��e���Fc�U�e���|#�˩X����F_��"~ph �3l�o��~���ud���վ���pE����&���G�E[}��Y����ɵ�� 	�ORӡmT�O����i���~�Z�jw��U�=<���/�Zp;�0�۷���2%τ�܅�Do�A� 8n�l�_��cӼ��$��t|^�i�x��]7d�#p�6ä�ì�慤M�7������sy/7Uɹ�z֮���'݃�s@�,vH�$e�5�6N]	-�G��[*����E�)� =a �����U�� !{&����X�\��c��&��/�{�4ͼ�.����\�]��#��K?{��fv9Ϡ'���}	gM�I6�V�� ���Td�B�B;O�D�O����O��U����q��_hˌ��)��p��!r�	�əzT��@��X7!��MR��n7��&>9�-��n9a��`2�yh3r��KP{!]'X�"�a�
�FTӆ�2`&�����f�ڂ�b ����8S!�jd�Ks����_�I�`&�a����d��l�)� G�K���[=���O"��5|�e�@HF/i��}6b�rH6�߄Hi�jꜯl&2o[w��iV��������V�I1hJ��M�|cW�K��F���]	1�#B������7����S	��x�>3I,�ThRM�H�s��G`Ar�obd��$&���4��ҍP�O��C拓�(&�pNb��x\��j�g߶�<���A'��0\�Q��%��'���;��W����o��plZ��E)����y��)�z���dߘh�Syco���R����+p��ɒ�0O!^ S�·�(��+�n>q>$ 3�N�HϢ�dY�kjc���c?*(�d���������IB�r-R�0�ia3t�	_Y��x�L��F=���\��Bo�M�3$ݥ
)�˝(�&V��@/��i�r�縭���ntޫ���6Ê��_��߽a�Ӄ1ii]_��<���ّ��VV�(���pC�LTp��͖
����e�ǻ�7[�\���FN�T=�����J��(��e8Y��U#Rr�~
#���f\�u�z�Y��h��@�㲖v��t2����	iy��ʸe���h��ٵӆvb��h{9�ۮ��8�$��;��lwZT0_�Hp��l�D����2�`��B1'�-�c��	Oc�	L�K<�c"�~�M����e|㎁˖���5���+si�v�e�̂�~�c�{e������o�w�;��T��YW����\G�_j��Z{�ar�N�V$��r�6p�F�E�|c ~lu~�]�8J2ّ�9�B�Y��x��-����P�%iSl��e������A�m�h�N>�o�;H��B]�k�vҝ��f�Y�\	��V6��w�H?`���3����N�H	�MD;�C`��
=0݅��R+)�^�)�D~�ڀZ	�X�������ˏU�i8訉��R	�_WN$J��~vqH����1����	��c>H?�k��<@+�{:������a�&�y1 �~���u�&&�c�^#�'�*��ÿ���]y]��k�s��>���T���EK��{���jMq>�t��#��A]��Zf�0�}���:�΢G��A�fQ ��΄�Չ�%A����/�L��hQ9�8��)�UN F���Q�sAܡ�,9[��`_�s���G��c�kT��4�H$P�`Ҩ��s�Fs0�"��zCS�;t��u5;�m�'	zW����#Ҹqu,�����/�-ᛥ�Xsn'��Ց�_�%�	��sp�MҾ�r��������4pq͹TӬ܈������U� ʄ���%��-V��R�ə5�rI�3�GW�9D���s��M�"ұ��#@r��㶢ɒ����Ū�z��\�.��F�H�i'Z_(�J�9��/��e4���Z��*H��0�p4�%�{o�.��ņ��Q��[��GЀc7f�'"�������>�]��&����˪�'�@��N�J�%n��
�L���W�qGq�i7�oA"�!��Ҽ����LFZn���P,�x\��C�Zi��\�Wi���PL\:d�s�&oW�#`�.��sXd3^�޽��r����M/f�7c����#/T@U<��FC���1]���d��@��Ah��n��E{ء2�	��� �F|/%0����v>�׳���9�ut�ݿ҆�2|���cnY�6*�DP�9���s`y݉S��R���P�Fop�k8"/ѳ�[��,��l�oӂp|(�L�+΅�e.4��H�iu+�J��2����7�볷&���)Ȅ黡j�a��ڝB�>�ZN@ 9�cW�Ì��2mez2�ңv#�[ݙ��wE|;Hě�$+U$f%�	UQˍ:�Ԛ�V �	=���D�%�^xI��št�"lJw�K�$Z V�D�ǿA��˫&�{2�q��#e�'S�1�<��nu;�
? 3ꭾ*9����j	�@J�<�B�,M�r@��1e[.ij�����A�s�e~��s��@��Ty��!"�H"�g(��v��:%��# �_��[5�����;�����'UȦ��Q^�1�
t��0����,�~w�꽇UKc�n�} 2�2��I��^��g<a����V�PK0ަ�3��,]O�$n;>ܣ���&(~:S��h�O#�����cRF�����*-�#�7�V+�:�};ȓ��V�1�]��1/�w���`_vυ��4�L���ū�A��#p;\�`#����zjڼl�/�ܱ��<��M�'�B�]6Gm+����<�� �Å�:=Q8}�r�9(?��@������YV+�X�B%r�'���mp�H�ϛʹ�V|��� �M]<��x!��%��Z��+͈�i�瓠,U�J;�qeU��P�-6�l�ӱ\d����,6�UGp�v����U
J��`xۀgi��a�~��~�˓����OۻO��@,���HM����ԩE�,YxQj���S,����}۷�Ŏ�������yb���Fq {=ǝ��� Y�8�'(m�
�f�I�I��f�bʶ����U���X�)
'£�s,�4��� ����H���3n&�u��6H�53�gmУh{�k 1��f�3�U���-��Y���P{\!E����~%a�83���j�g���ڊ-p��"���R�̑���4V��٨�:͔)��U�꿘%���DLuʮ�n�1Bv|+eN��W�t���4vK�Ȑ�]�taj�	@o㼐i���˦���k�.���d�MB���A��p9M�� �B� !��i���� �j9���u��R�K
��^��]ӽ���_5�zv�����b�+��u:�:Pt�������*`�T�o�	ƨ��Ρ��i@
��lH}��`��n�_B�ͽ��dMzG8����Y-�د��H��ת�?��Q���5`?K�楫|֮8ejķN_(b�g/�R`�z¿���+�=��ꁐ�m&T���ŧj`kmayh6���m��}CE��a.O���j��}�p|&����Yr��JECr�m��	�)�7�wsۦ~��ul�q�t�2Cy�g��`*�0m�ܿ����@3�%�����毳rj�������3�,=Ő��X�EŜ�=�q�G�Zb:�Ⲱ:�L�B`;��a��`��>K�JG����AW�C�co.�^�rp����]Z���u-1�_��*t2vn&�z�������z�Ξ�G�G^�)���4��MѦf�$�6��q^{<e!�M��N�i0�xz2��9p(wU<�N���R�v.+'�ps�,:&l�şk��K�H�d�%ga�6����s"0���h�&���-Y�����D�"�P�.C��nlys��]k�k��ew�Efr�_�k|���%��Z�;���Ð,IPn�G����n��gXߝ��9�,�����@N���s��|8x"g:RU�9qj�M[���Z��-bRc��]�/`��-��$zþ�(eH��n��Sq-��3�y���*�� ~jZL��TJ��ݍ�(��ްg��L��qFĉ�x7S��>&�d��|H��\(��%���3e5����l��$<��'	^�s �L�_��9P~@=�k�Ԅ�s�=�]���ޭI���ʿ8�1��u]���)]�/fP�Z�4&K�r�j���fRB��
��{���q��G3�	��Q���>@^�V�$�`%H���ؓI�@,�]�H���Ur�<��W�K^�жn˳� ]���^�5�~�9aK9�c1����B2�,A 2̶C�<�����>�3�;Ó�!��͔�`z���bʹ)�+��<�9�EQC�:�q<��#qq}���qO�>�3Y��>�����9�C����ߑ�zB��GjS˶��� ��H\�?S�v����r�C�î�N'��ޯQk��t[���]
	{E����u�z��lj!��83�o���|5@zH��@[=М�y�~�}�_G�j�.�@\xsnU}�;m:-^s�Ş���[�q^�32���8��{q����c#N7��$y�^[^@��:�֟�Z�_b���s��*�I��1CpPٌ����x6�{]E<��"��dV�b�Fq`�����c�H��Tk=�~L��Yr��j�e�zZ��u���U�u���M�r3�H�i�W�5%�[砷��np��W>�N(�4=�L�7���<�7�Xʛ�� R�Xձ'�?�y&q�}��E�Ix��e�C����ls��X�s��y� ��/"���
�������l�f7.F~����I�by���7�*Ę�j��c-Y(�9��US� ��$���L.f~��?��!��(+s�2d�2�*��pO�A���l3��&uc����f�)�/`�'���c��mRO�B!.���?��C	�:?�9=����P*�;��m~|L��ʇd�p���D�4v}<t& �FUy��P�oU�M�ǩ�'e3Ӝ������60�s��P2.oJ�\��u����+jy��]a0���D��of\@��|�@6iF�!׬k5o�$�y[[L����!�P�y��Z,H��ȍ?�� �ZA�~�N�E���8�}l��ߗ��43\�Qǵ�HG�+,��4Ǩ���@�g2	�z¦U6��� �
[Ԁ�Fw��֖t�Nеt����;o�~��Z.Je��:����gۭ���^�`�҅��A'n�o5R��&���L�De$EŁw� ����~l�J<��aT���wu?5w����n4s�W����`� ���l��A�c~$�Z�7r�ڹ��P���p�@�#��(��!�M7+�6_a�懲mY0�,E�-.V���0�o�F,1_� �o��P{U�#b����Ф�Z�I�-aA�K���ƒ멢��B����VXr����D�b���jl8�Ef}������z�w���� 0���4]���t�"�)t�z$"�[Q��{�So�֑~��p3���k�g�
V�y�����9��@��r�y��}�b���m�~,Q3"���|��ze!�ca3�1.T�*�jh�ԝ�z˥���{�ʨ�kR	V�5S�7F׉����6�q6�i�,{�qi��O؀�)M����w�̶�;uGG�!�EJc��vX��l���:�b�̍��v�È;�S}B�i�d&�l�5�^?��h,�TܶdjA�r��j3o�m)(����T�`�"�"�oJ��r�)�	�9>���~~B���/�	l�zv�7��lYǆ��\6Q���nQDw��b�!��Mj��ˊY�|����٥L0�����P0���W���@J]Q��G�1��!�?ƌ�b)�O�sq4��a8q��@{of���!�5�z
	8��S4��C�b�P��A�t,�es0�c
���gÂ��.�`m��]_��w��D-O1)���CKu���7�?���N_
��m�xS^�~�hU*��}J�݅���^���q�N�+&2�Ρ�l̦��}�F���Xv�~Ax����A��H#֛by����ؔ>-
TtNu�=i.A�'$��
�3�ͼr��L�N.VX���̊��NO0A��{�D x[�T���.{ǅr����gn�-���
��1�? ���L���
�?j�A��]t�`U�fܦ(����#��y�D���n���1�L:�^&�)N/���Lk��	�h�mX5���}�.@��v���r+ݴ[9��c�<`�����Bи�^=���CR]'�����v�Q��v>&(/��)�@������Vj/�EW�?��?7}������ST�u�>\�F{̭������z:E�П�wy>�f�̈�5�l�\:��1��g�ʜ�@h�昅/_zҼk�)e�{'�����K�)�8\0��sB\��� S.�A�e�n7�ǳ���|�\�26�-E%�t���U�=ݭp����V������	e§U��cn�?�O�O�����'�:�(�t!dJ�8g��۷U�۱�,��w���H*<����N�C;�qCm��Q	Ty���E�ۀ�#q�j�wX��t](D����F8>g���|RX[��|&
�c���_�
e����|�v��5.	�-����rD��"�j���e;�5�A���ii�Xd��^.��a�ѤT�����;�����fƸ�H8+R���=���x�g哞�{C>/�:��W**�1� /D��)����GƵo�|���Oj���d_��]�:<�S���Jg]�qI � p;��M��$�&���_�E����x�����(Ʋ ���9���~�~5�z�8	-�
����x<9:�N�d��x`AUg�/5~Z����dr�Ϥ��3�A��S��k�ɂ��&��r�>;���̕yFvG�Ƴ�\@=&ƣ�I���x��L'b��s�N��J?��[�s�;��<������5�L1���֣a-���o�������,O��'�X�y#X��ۂ� ��a����z���-��?��̹߳�$\H�k��vT�eU�xVR��p��jIy�+�VRLľ�"f8`@�|�9*��xwɢ1|��sC��H=��س��Hiḙ����R���� �]�OJI�7�E�=MW�q��5D�e������;��涁�i�pB}����s�t�bw�D��+��b9^���V��w�-*����;��.�`z%�v'ă�+��[������U R�mX��Zl�[����R�5G�{ȮQ�������άx��SS�E
$2նz^oǴ�k�E���
�F���W��-�0:"�����3T���s%���1@˱E��|�<�x�>�ЃJt�_F*��Č�����������I�=�խѰ���8 $�dr�z�x��B-'#muxݖdc�e�$�&��d�s�{P�� ��C��(Tdίm�'oah���@g��1�b�(��2�����s�H�:"ak��x�Y��uVI�kcVɭ�[T������p�ӈ�W��3ձ.#�x$P��wC��ҽD�󍴪j�-x�c�J"=�jN�sTCu���;�`Z����˧��G/ Sٵ��I�ϗK���;	*�C��l�]>��Bע�t�vk"�d�_�7���|���0��������K��Ҕn�l(���vѬӰL�qܳyn�Ju�����=v
�Ư�G��W����$v0�g��]f
�t�S��N>��J曊�ګl��S)yw�1�5���V��=�u����2�y9��E���[��j5�3�8�(_w�o�^t�;?y�A��� ,QbBY@M���+$�9چ��G�
�##���8J����v���^co)*컔���w��&.[3=�\טS�a�8iܵ򈄐wu��Щ�f�e�\�'q�v�D�3f�F!Ԇ�==��	LK��r93F
ŗ�6�mJ�ߒ��>��d�U����Rw��z�n�ӱ�`���[@�Y��%_��ct	hU�PV���=Z;�z�Ѯx8�c\ZtiR�J�!Dq�C�����̬��n$��&՗���"��Bb�;q��$~=Q�N�"�㺗~��h�	�����߉��a��F�<���ߖ�[!��N�{�l����T�0q�A�m�VpRuV>��DwF���F�����2��Dx�<3U���J���_�����������g�=�ؗ����M}���i�Y�w��Ԏ�'?�aMm�>\�T2��ۼ�"⾨o�'������0�a�ᣃ_���ph��
����(]����V��oU�*R�V2ƙ֠J:S�^'V���R��6��-��3��aY���.8[Ҵ
������!�:� �?k
pI�<��y]�¥�q@
p`^Sta]6��o��$�\Pr5S
F���9ޕ˨仂I����\;ht'y�H�)�Չ=|{cE�ܜ.��A��DG�
���3���:�>�����	3WBh��24�p��$�$���YIn5;��"l��|t��;[Ȱy�s�.�y�M�\s�*���9�>Am�ٓ_�X��l����UːI���Gc�p�Y��TQ���0=��������ƴ5ÈItsT_%�֏�M$0:���ҝ[Z:�c+��W�Σ�3t���*���Υ�zX��{��VL^�<�U-�
�����د���`D`��$Q�I �<�R�h���j�'l#Qk����Jj��.-�$``�:8F�,�������T����y����z[�f��R���>-#Z��WԀS����.$��Pt��.I#�D��j�AO|��]��x�$�QC��M�bS��o����譎��z�b@�B�
��O|:۲�O�B�js��᳏}?zKW�tz���Z&�Ł�¼�k���[��e���:�����Cs��&?B��?Z
����w.cy"d]خ����
c��j�>�}��j����
eaH��x�-��dY�76�c�,�:CK)rH�6�[� ��V�칃� }=uJ�1$G���4$��$B^8�S<!8WR��b�şi��}����x��H�]��N�����o�2����'�My�>c#ΐ�n������wLa<�!�c.\g&}����ʥ�u'aS��TN�����͹VzJ�EQV��B��?���߯7KN���)	F3��.l��HO����C>QH��gf=���§լ�֬P�������M�?Y��t��.7�VU��gcB��1�\���I>o��/�f#Rweȍ'���-/�b�t����8QQ��3;7O>�g���y�}��է]E.�V[�aJ���$xe!~�����G;�bܑZ���^�Q��Ap�E��/�Ou�O�YBi�czjH�A�
 ��d��kg�%RpL�WMڀ��QX~a�d�O��CY�J�A������7�ҫ���I��<Ҏ�3Э�>]����WY��g�(��J������u�x=�Ҹ�������2���H�M�7X��٦�r�Mg��3@a��%�P��0�AຳA΀Z�����k�qm��ÎitJ3��a$�Z)������ ��Ф\����l�Pa޻�o�!���$��=��/��)��!�(4�|�a���k�����(c-�"]��}
��(����cCI1�q�ۑ.���I�s��H H>{����[�e�����r��L�ǅ5�;����*�4��a�w��^���>C�\�v;$"�s�Qn���pe�U��ՄT�?d�<d��[ybxƙ?�S���̔f�a6=L��u:�qk�g�\�F�+\P7��P#�331c��d ��.Dol�U������[b#�o�G��<���Z�^�����q�s���D�P��qQh��AD��a�ѫ?�f�}W���E� J���Δ�.Ap>�Ր�uyϷ�Ҝ����O��6)�t��W�|c�m�$'a(h��g#f��e_���8a���B_ǆ%5�T��+�$�!qu�nӮ�&"|�Bj��Խ���U�`�E#��k6���R��h�T�@XX^+��1�ASA�3jx5�kXS�G@�:S���
�Ǔ�2&�v7�A�	��9��'
5��2I�M�Zb�s��?��5�����4�W���}��k&#��<69㍸ z�?�i��c���������:��Օ;�uu��=s�q�u�+��6�`� �����{����dݔ��gpO<w}IѶ�T1��r��>z/fS�R�3�R�f"���
�ɏl�3��_*�Ic��ȫ��;�a��B�S'��h*U"��Y������&YC�l5"x¹���
��6��_r�Tᇼ�H�<��(1���D��U���h��:%�f<�:�pYB�s�Y�;���g���:�*m��yxO#��;�,:G  ��G��d�^3�+U��/��������bƐU���K���?s \ �{�uD�J�� �@�Ѝ�59
e�������ʋa���!���x�4E��$ϑvg!{\�m=���X��!���jcH�R��u)�L��&�������Ľ�xޕ� �cF�z�t�G
(S�bē1B���y�i��Sp��~f��b�ϷJ�-��$��3�8�����,Ab"��8<	���[�y3���A
��E�fȧ��V%��_4KK�@>�k�Xe�[x���E%�%��P��>�-RhN�ն'�O����HA���9T3�8���ࠢV|��D�ʟU48��E~��X˙β�PP�`P�3D�vT�6%�N�}��"���t,cL��-��%Hf��?�:�	!�'��JӼ�T���$��r� 5�Q��OI� 3I����K'��*�|����F��:���变�_e��15?���-�)c�l��"]o�����H�B7O�8��>p����#N�KKW=z�j.��X!X���p���.�qn�o�#��?y.z�3k��#��A�,V�aF�>/�̀	���(؉�x��9L��?��YD�>f�%b��b�c� X����j���zVAKu�oZ<����(m�O��3��M7&+�%c�/O�N@8��<+j�7����E�������5���p2A�{�����ĭr��ԅ츧��a|�9QǇ��_x��xT���ĝ�zk��FeR���;K,��b|c�h�\�2=�=��`2�O%O���ei:��F�j��&�؀�L����.�j<�\G���w«E&��jjfe�;|ƌ<.���6�s�6E��7U�p��-����p�Xg�V4T���WΌ,�a���án����7MA_�`�j0��[�H��mA���; �l�q�2|����V�i��9��y~YUL�YI��fi/iAKW( aq;�����E�Ғ�x^I�7񕥃L׊v����P���(�S�ꪜ<���e����Ѐ�g3sNY�r��8~w0ɭ�˹@5�+֚X�JX�?����v���-�҃��T���?g�Wo|�v��K�g4��(�O�Z�to�o���|e�~G�H��:q�������K��F � [Hw�A��!͂)�=���ߣ�ZF�i(����l@�J)���,�	L�g�6Fyp�_lX�q�²�J��^��^���ҕ����)?̸��F�����STp��Q�x`l)SF;����;�V���7�
��C2�P�����j0��2L�/��v�3*D�[k��L�	xJi7w�ȡ��w� ��ͳ�^G�M�hTȵ�g��;��d8i�/A��m���׶`SCP~	SLz�.�fJ�qF9��Y.���Y�R�V��m��V�ntƔ�;l�0�+����X�� _�L
��j�;n�&»�3��0��@7�&MX��˪�ͅЉ1�ʄ�%{Wש�:�W
�l0a�6Ӹ����qP�$�[��*�`)��T�'�
Or�����XI�u��c����$�g�j�Pp�:�"[S-��̉��ht��A� �D����1g�I��s
b�,������#F���ؘ�p�u�������?�~�(�Nz�,&�1�.HNśV}��*���j	2P�X�w�Ӕ�0s�wC�&����+廫n�놘 ����_�f�`z$^HK��������SH
����/��J+$'���ټ��Hj�#�-X@z�W뻅0fo��b9�S�p#t�RG��w����m|n1P�o�ɔ�D�E.<����ؘ�T
D`*~VW�� [�r��z�ja
�֜��v���U�_n;�g��_0�8ri$�i�#���W��(A$��@o\���[{�'���}�D��G��ck�Ll��#n��N2`��I0E��d�H�g�����b��W��t_��h[Z���r���ڝ��,�q�Zp�G���%^���
ixR鱣S�Zyi~��m�Y���o)�VʡɰF��i�u)u�/��=��Wb�(A�U;v��Q���fxC��?;����0}�������t�$���>�����o/�#J5�7;���kM�Π��cI��s���5�q�ԧ<--��j��I���;��=`s�K|R�a��ڊFg;ׄ(A�ȕ#�<.����@�
�E1z��Nn(hi�L���l�6T{�*���Jo���`U������Xg�>4�B׻j�����0
m�c�ƒ�4;��:D$�GLLo��cY��wn�N��U����7�����i�����`�*9��b5�}��)�9g��>@��(�mM��~��� ���@#����!���i�����d������,��X{�xא`~��y����j�?s`���P��*x���3i�%#+��`X��玆��1���ȴ�,�>������E�&�ۡz���Y[e(]�L���y^V��*�p���)2�X&�+�r�d=`�ߩ6�3�a��7	��.[��z�(j�u%=s�%��43Sea�׬v?�����W��S�܂��vڒG5�lV�4#�J��
.x�S�������*��q�.�M��ԯ�N�*$s����7�M�%i����C�.����k�9�Ae�Uכl��	�J����^:5Ǥ�X�B��&�b��Co&�Z��R��KYϠjb�39�K�w�XDj�����T��T.H�^�#���'�XFngpE������s� ӄ�sZ�B4 k�v2��>�@�{��c�v&/ϫ3����V�/�UFw��i��~D�I�8R��$�u�48�Vz=�
�bᒬ��P�e#1��N��:��w�D�=UE1�9�����,Űa̚o5�n�2�$�`�A�$1,��uM�o�狱�1z#i�g^.�eX�OB9�v�b�'nd�L,i.jA�!	ʎ2f.����!�l��o�����u�+xQ�2�2�ܽ6ES�����yGMއgEA����mv�J�X�]��Jĥ�������=�F]��ޅ�	�]��\Q�E|#���:�&W�b��%{�w�'�o�6M�l&��'k�z��G��p�%�*�c��	t�?�5�0Ӏ.����v GS��VP�k��A#�j6�3-�$rt�Gص�?$������?�z�Ao��K ,�CKz��	�����a�7�fn��=�;��%��}-S��S�k�.�g �Tb��R ^HJ̣��������@�X�3�qk�+yKJ�&�|��`}�i#����u<wK�UVn�1;�N(
���R�����#D=���O�6���L�$�{?��V��V5U/�����&�"�UJ�A�-V̟%���.�+F��9��=u��t K����)�-
i�1��I�����2�� �q�ZF�W0�I`���2���1�"��{<|D/�6�`��G������������v|�Ml�+��� ��7�����.��CS־]������뎙�z'���#����y.{�v��4�&p�J*���Q�-gxva?t�e���E��~H��2R
?�:;φ����� ��u��+uk�ޤ�u�_���x8
,�墯L��A���x��;��uǉ6���Y ���xÒ�i
��,!)�~\���.xQwWM��#�-_f���Uz`���")�Kg*����-GC������{�̰�c��vv&W�/�.�_?\�܈h��ƫ��:����r_ C��rZ��A5�&k���r�~����dS'?ZϢk�AI���r�e[I��C�B�8I��v�Xoc���Z�:�ɗ?]�L�R�
�L�K]�QN1�M� `~�l2a�V�-���,m"�V������*��P]�IG��7���	�ۜ�a	|-�Y4Һ�fj�x�U��i�X|UV �c����n���{�G���Z1�5|�'Z�9�:k��*�����?t��>���<i�F� W�dS-�YZ�_v�\�C�g�+ǋqf`�=xO���q�4�l�Ӊd�®�9Eԭ�� u�狫&׃�a7\����3�?˛��W��7�S&�;`[�zH�`�F˥�"$�;�U��.����kߢs�N#P'��JZ���vQ��:�4�����؊��潙n�^d�;\Z��U�n���Ƴ��"���Y~�Fm�G>�!P��G��M)�3"^k��,�-��U,��!�^�a�`rH�78G`z��X�����C��#���yW�p�
����d�TV0٢�d�b�ZG��B�\܇��ߤ�UNt�V��B0`ISb�r�/���D�\�+v��e��Nn�?�6�?^�qk H�l.]Ҍ|6����3�q�<Ӂ.d8�&�^�d�W%=���ȩ0E�~���V���ܣ��/�}+�I�Ū��0
����n.��ۙ�SF2�2����L����A�[�{�3aG[trwQ����Pk��r�a	�]j��wb)�����j4��HQ^O�Z��Ui�0�3�G����_hS�Ѣ�����mz1ZXy��/�xSʚ�A��_���epi6�G��s�Y@gˆ9 ��G�֩�y�v�6f��i\�w'�_�+��e!�`�w��o�<.}��ְ�eV��-�M��'_��깴����?NK�ONO��1����K�<D��}mBNg�aU���^0�)�Z� ���'�xO�X-�K@��O�9L�����m�F}w0��}�DOƎO@�R��5�,?�ޱ�op����^"\D:G(;��AY�H�ab�V1:��4�g�Z4ll�e�U�:��B��U#�pަ�o>Yt��=^�:l�ކ��"�v�.�+s��R�W?��R��jQP�&d�]A�G�145��D�Q�T�C�YNq;��4ՠey��4)��ozlnC_j6��iseߋ:IgC�g��!Pv�c $�a��Ɏ
���z�
�nJ)��ժ���r���ۨ�ٺ�w13えRl��L>��A���e�W[@�|O�^A��C����oN�J����w��g�q*cP�R����'r!h$��>��}:�����	��Yײ%tJ>.2 '�0���M*x8�D*���+�'U㴋2�됒�]3�glGs�e�h�@cX��?�n:v
l@6a4���`?߄s����>�Nb)�=�~�D<m �k�WU��� ��:M)��~ɮ?J���5�?�3"1��{�r��/+���o�r� h�e�]=3vY[U�%II�:��l�*������p=!��1G�ft94��k�2E���,�1C�`�����Q d2�Ù�"~YƘ)��I9�@�y��_��U���zN�^_�˯ķm��YE7��V�be���~_��0: ��������D�m�`QB0��-�