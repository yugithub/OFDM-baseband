��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6߻[^��3�%?5j0�`�Q���֑ﴔ��K�z�����T��Y���69�9��潥����.؍õߢr(�D�e����Tui裆�Q���|z�L��D��{LgH��2z<�v?^T>]���`
�c+��@��t��b$��砆����#�r<���g(F���ƀv)/���� �15��	 P� OL 1%\�d���:aq���uB)���+w���YZ���?7;{���>-*/�f�}�C��t9;��"[Y�A�ͺyǉtFD�˟�m�h�ӟ`q���*�K!���$� 3��Z�:�y�u=u����=,��cy�Kg�m`
@DM��`,�mzi��Aظ��gO֌]mi�
�n���t�p��:t"OZH�c�h�f�H�������d�X��gF�����%�p�����c��Nm'uY�x�B�I�S����C�:)��lu� ��f3x���п��a���i��Pɟ��٠"��ID}dO���7K�:��ot� ��&	�UkpӺ�>qj�w&{����7XǈP.Ov�-Ѧ7�@[Zk�����c��C�p̡��-UGY�o�v��o�}����{}��0�X�L��q�����#��9�֊����������c��8 �˰� qqd%�o$����d?9m��x�C����
�.4l1n9�7�F��~wʳS��"���v4�!���D���9��y����BCR���&�$�-Y��5�a�����9츬�YCj#_���h���OR��̅AE�<�u0��]�c7ZV(�v�p�P���P���ivǰ떁�â�6�N|�J�?&vt�)�:k�$|дS�i�<Q����>���\�^�J����r�zV���{�~��fN!���H1B��ȪX��������T��P�E�X#	fG5o�,u�.�̨:���~	�ډ����4 �B^��WY�i��ю��+w�n�ϩ��^���>��D���z/�w�F�P����X!����E�:���d��¸t��;�1�{��MM��,@��uv鍪� ���P�h�}��Y�a�����ZE����R�L���hj�.��	 �Q�BoZ���ۃg#?2 �w=��_n�$J�K�Ÿ���R�D^��ڌ�)`��]j��U�?��g��o1Y�AAl�s��2��y-$]W����.�:m�/��>��8k��Y�I6��fF6����ZFn+'=��\�5S%�3�}���7R�o	��-�����Zv\�N�R��)����"�����d��]6�@����s�+ت��k��7�c ���w�Fxb4�}6Tk�q��ڎ��{O��,�5J9&:|D�I0_������T̬)F#g�j!������(>�rC5���Y�[2�B�N*>�.�O`,k~*�Ӣ��Y�����A����b�B��9�:v/�?)�V�M<i��ۏ��=0�|�.�~� ��O��
�x�VI��v��-�^�ZM�V�Ӷ"Qv���:-���ya�U)
�@e0���.�M�I��ģ��ʻ��ه跥Y�A)�!�f���f)�
<�+�`�7�E�D3�N��x!�� ��^@�'��T#�Z�1�Uh*G!�!2�C��%65��yL�2�O m4bf��\b?�<�Dm�ܖ+�0��M�}���ʹÝ��98�K+-�����Dj�Y{'Ҵu���c�_��L�e�i5گH��k8�T����o��d4&��j_S����R�P�&^�����ye���JQk���J/ds�vh��A�	�J@ۚ�̠��}����CrGC��A���W���GU����Ϟ����B���Ǯ�H�ҁ�-��,mp�EffOe!�~Fh�W�0�;?S� 	qk�쯸z��x��q,��nn�˰���C�#�b���ڱ.�>�%(����=MP�K(����
;�
�D���w�E7�i����)S�nT=�?��:����ӧ�z�2<�!�]F��aKk��=�Cm��Կ	gF�8�E)�lr`/�#X����;����.��G��e�s6�OH,.��(S�Q���4������c�bV��φ��� g�����{��<������u8m�$�&���KLIErr�7��U���p�T1�tr����1m�cFڭ��H��n�{��H��T'�d�n�c�� أ���5ĺr� �b�z>��2*�z�J�)i��aY>'�Ҳ��9�����	?�*^�5���kd|��?;j�u�O#y����c3��z&y�E�ZsE}A���5TN�޿P�I�'hua��TZ3���1�&��O�pM�2�?؜�o������ͳ���2�mX)��=���\ZqZ8��/��\��a����{��E,Җ&O}���sMl���W����ko�ɵ7>�����Rc�}.�&�bC6�k����d�)�����:��9%��Xx6��9\�s�dSr�
p�jG3�uˤ�����_Bsl_F��D�y�F/�BB"A�s�GM�_p��B���웤�3�$�=I|+�*rZ�ؗ*yҤ��hMi��,~Y�oǐx1�%��h=��p h�q�%%�4"Q6Fҥ#�����Y�s����n��Xq�q�&r5˙;M@����y��fI����xQ�gVLPӁ.X#�A6:U�$@� �{Rr��b ��G1��.�����Ҏz��hT����J`�r)u�^�_��+ob�J�4�!_N�@ޫ&�͑O��ܕ봦��!X�$Io�X��9�y`�:C)�0D�N�_X��?�-Lm�J�_ќ���F�$Ƒ�6f��.��~G
�7��.���\�yL@?M��Z7�HD���@�~�Y�pҬ繬n�������O<HS����!M���^�%�j&��Fx����if�! 2d��.4��Fit��]j������t ��3!.��|�Xi�χup����E`��N�0���.>�G�#<pQ<y<�d����) �BByc����k�&T�&��*���}�S��՟�(�B6&�����'�7t?ehmS��t��r#\/!�&��.$/]���pDU,Q��g�_̎Y?A� �����<�q[�:�'�Zs�g)$� *��Ǧ�D[q��
(��X�9	Ut��g��_꼈8��}�p�_�&�\{��Ր��ޏ�ޞ��Ȼ~��׹e���L \��MR��r�
^V������%b�@��d2�3̚1q����y��4S�{]�k��ó�\��s�>�N���b�>j�.��W#�`�s�VB3N�lhc�n�y�`oVɫ�t!..� �S|C�����e1�[R4�G�0?��L����N��$��6��k	kK�����]`�����.��A����b�X$8����I3���K�<L���06�D��y�*v�~��He�B��r�oV�s8Ӟ�OX�[>�H`�g�>��QE.��ɐ�����J#@�O���ӊ>�����Q�r�����K�ڟ{����	MV>�2�eGJyd*|�o�K��π%����Գmu�}ן6T���!��Tk��j�q�P0:b6y�6����KdN(̵�d<��\^!?uAj��w�B�1��T�w���m�t=#;�Yj%�����/�q���xT������eF��4�02N����AR�ޅ�SR��`��Z/݈Ȟ�<�Uݞ5:�|eHL���Ze�#�����m�'lW9vDw�
���t����v�Ɇ���We�ck/�:"tA�D����s�)0�Ь�!2�V���-�fMtn���DXT�;׺��u� !��y5�ғ�ق�H�	���(�h������D���=�2Z�9�C;6����;�J�q1�;��Y��$\"��&��
�fO���}��w�S��z��Y�F+�fЃJ�#����0��G=w%l%�]��FD����<��#���kYc��nj'Էx,8
��{:��HZZd��J�ضS ���=ƌ�lc;���C9�X�a����@����!�ϊ� j���%�q�x�Ķ�į�����Ǆ�n���9��<�şv��e�T5�i�
'������ru�5�ù ��Ë QI�����y뿻,!��9�z���]�^\=؂z�D&�4?>B�*�����&��P4:�K�"���#s���1@���hљ��z�Tff����n�"����K���Gw��H��z�;��Q^�)�퀔Mrh�ʣ�9ǵ��L�"���H�tr^���;:�{[�~3��E�t�AV�]��:HQX���"�A�8v���&�$�a1�Ft����Z;|��ɢeK��rë6��([&ݮ�f<I�T��d�hy^X^laI'�艗�ƚE�*+>�a��K�TH�J)���Dd��  ���ގ��͔��z�����kH��N�SrQ�4=�J��׎�<	��Ɵ�BPP��1Z}߯͞wxs����UKk���_��*t��a�غ���پ,L�=l�U���e����,*|����o�����RSg-�=�gg��<3� �i���V��pE�+���ix��^U���܊�ј��޷b�(=���Ƨ�1��0j���*��9V����5���7�	F�w��y
K�k,t��93��ݺ�7):���3�dw/�4B���k�W���M���5���lkP�T��#�Q�jtN(^��Eg5o,�.g!K�/��B���Q1̌,�;�Jjh#K�IMP���3�ڨR?���l���@�.�kC��MX�A�l��@�v� C��{�u�ZP:B��}�K����U�ӑ풠Г0Q���X�*R4�[�T���Pv��ƪ���2�1�E�2�A�8�p��1<����&��^��*�8����~�:aE���k�X�C��#�}gĞ'� ����?��"o��.�k̶f6D� ��Q���@��Q�n1 �|ʇ�BQz�n�:�Ĭ���^����{W�L�ܟm�M���܃��<�P�)�k*��f�;)��l]�/q}m,��K\J;��^ڦ��;���Od`�����1"/C]d\	(�=&�݆�-t��c���+H]��%�I����T[m��Rs��o=T+�҉�c�9��?Xǡ�k���	NH��`E*�3��̩1�mF��`r�b��P��� g}�����iR.�6r��g�]�LIb��������卫����`f, �u����g�T��!�7��r��������>�Z��k�@�t�����!�O�y����,��P��P=W��i To-n�m����UW�Y����Ox�h��s+����xV3�߶��B� ,2ߙp  hN�?�7�%�G��}�g�`�!>73^q�	��vZ1GC���=u�}�Z��+�h)Y��<@<(�c�:����&	���4�4�\�b��Q��zi�k��&]xlI�t:,5�k&�~�*��X�O��9<�v����8+�e��={D�rl�-�~�g��$N��Uxjm�G*ן�O?01�{�U���1ix'���B��&H@����������C�[�Y��ŷ���R���A����P���x[ˡ���~�����=*��-�a#i��|%?Gi�K�Fߏ^)	�[��T̉��*~�9�s�v�44�̰c}g��I��ѹ�4.y�,���؞�n9�O�A������lE��s�O5U�ݽ�Z��Y�͑��氱��[:�c��8m�~�y<����m�#���t��WdJ1~�P^��9���H�2K���)tȖa:s�_���"��,��E�;<��S�S(��Q��i�l������@��=T�U����i�m�2d
[ŕ�´,P~$ѵ��G��G�����&�Ü� !��6�5� ���LĮP|������M�$�/�T�%�# Qw�t�i��R6�Q�1	i�z��0sށ�	��*̈=RK2���|�!n)Q�&�U�m|���{�x�干8��&W���*Y%<�a�!q_)>�r�����N2,�
����>Kn�QG�N3���v���6u��y