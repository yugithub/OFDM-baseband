��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|�����F��v-*t���=�O�b�$�Ѕ5郻�q�LJ���PHS�q�d;S�U���6-��^�NN�� ��	�/�5��8�g��k�QC�\�Ԩ��PK�M�� %�X���p�aL%�I}�S�[���*N�s���4�6�?�c:㯼$�j檭�����Q`x*P �?Z�prq\�T\q��|��I�G�v规Η}|��*@+������{�X:S��Y�z�I��0sd��2��V�\��w|��m��-�|�}�?^��2�ԅ}��y߫��3J�-؝tz�VQ����03�wk�2���CF����s��e���Z��4,j)q#AzͶFe:������V�sV��X�&����{9�W`�؋a�o�wmD�Q+�=T�ڮ�e��`g�۩E
�,��EF,��͊�������t����Os�Ӷ������<y��E/�c�'��l���!vr�9رQ����j�i��I
��x^A�m�ʠ��m}H�^��B��}�<�~�R�gj
�@��_� �����emO�%:�B_ʿ��ᄪ����H'`�V~EI5��%NG#ȅ����G�p��x�E&��*;�G�4X�l����oJ�ϳh�P>[4My)��3C"�ޟ'ޛ�f���e&��_f	�n^�Ͻ'�ر_�hd�.��#��4�VS}�$6�u�ûV�w�l�,��V�z�K�������'����c��	vvI�̯�,r���U����u�|ۡ�8��ձ��#���Q���2��� �%���ܴ�^�thT�p��^5_���Lo�g��f�V
����?�J+��o��XB����e!| BF����俲������0m��mx���|��\�UV�/��.�J��hW���d�\�^����ݜ"�p���sHw����O�����a�F,�(��k.l�	9��l�8��bǥ�>�w��2̏��\j���n6q/(�j߉n=��uvu��5 N��	G0+t�ץ��<�]f2�R��*L�Xr_��+�Gɒ6�o|�JV���*v
�7=:5�xϬ�'�Y14-�N���_���ŉ�Fyb�k�����U_T��;ݤR�S���k�N_%�Kj��|lR�������_txR��%'S�{
Q�c*�~�P
��s��%��I���}�|���U��.�!���N��>�x��j\ʖ*�斒�5�����A]R���".ΏNk*��qY�f4MF�1Pb��&?�x��\vt���QP��������e��H�x��Ƽ���3�pV��fKɡ�����U1�DK�%k>��!쯚�^ড়�@)}/^�������u�c�`p�o�=UW)>��1��< U�q��g�u�T����� ����e1p���u�W(|>��_��SW��n���LU`$ʕ�<6���H4ٝ]��k�m�;4�R�\5:G�a�#��� h�R���ؕ�DA�ɔ���~�6f��s����85��Y*P�p�0��Bʇ
���WXᮾ]Dz,�������W6+~�"��ʋ�j�ۋ�?��r$qϯ�[��9���J6�	�~w2�b��@%;�.��!- L��4-f]��\�'�?N+��3`.����6sYd�~�>�O!�Z��k�F�Ɉ*�c�:z��d�d���n%M�
��fađ�.�M��6��:涤`�g���K�\:u��[�m~I"��	އ0��i����ԃY�;?�� �:|&�;kc#��"N�}z�{�kM��?;�3�}�F�� �L�I�#�麈��"i=�"�R&<�v�l�X�b<i@�¬�d�VP�,~%����f]���RN���>�R��)T� H�4a�,
�S�OIm��N��}�ԥ1ͻ���/g&p��?�a;�m�h��GmF��-�c5��B���ه�U��f����2����
d6+���<l3�.��"[,c���}~�4r�9>�[�g :�ͧ \���z0���Z����<�������[���}�	Rw��Bfʺ�ցG����t�1s�v���q&ڥ+���K� �I@~�P�H�>��m��>�G]ϟ*��㭖I�>K�� ۂ�;�6�����H��y��Uj��?p���W�_7�xUq	��I�ֆ��$IKLEO�=M �I�*����#S���1����W6ɽS�ߟZ(3� t��32;m^�]r��DB�K�I�
!�Y��g��c�]+�{��M��B��َ�м��1�%���5�a���t�r�ť����5W����U6 h^#!���~QA�_Q�y�ޖ����8���gTSY؛5F���i�=�yr�^�q�	v	����uy%Ṃq�$5���	оH6p�����6�%���y���ri���؃��B݄����X)x�a��'��U�S�\do�N�L�ìP�jiɾLi��S�y;�^y�_���΅�\9$c��k#�*�u�� rt���.��7��O��Nt�+6�ӂ��~�$kO����;�g�cz)N�oD��3gᏆ~��n3�����#%Է5r*��>C�
��؀�x�-�2�7�߶a%?������7�d��"=����TH��]|�H��� ��	v���B��QJ��[�-�h`�K�_[-��+���2�W�r_\��H"����Ɗ�P�2CDz�cVa�(Aܤ���K�%:%�'��W'�����U�(e}���E|s� �C���"���4rȸ}��	��k����V��;G@H�KۆiU)�י���P٥����D�6�I"�@�.@�c�A엽���luq�����\�DA1�&J^[�+m��8�1W1���y7�3d>���X��gs�F�5
�9v�����1BV��u*��֩��&ej�rd��-����3πc�Tr�;g!��'���������=L8Z����UH�M�x�O�e(X =a��갿���9���U��	��!x3�=��q(�ά�a�v�A�`͌FVp��V�� �@�˵���#����&�(ׅ��@�����sA�Bto�ɩ�=�V>���s�D�Wt�#���38���˴.҅��}kI��0�8q�8͙&W���kh�E���P;�<@����5�k��N���y�
���4vNL���+9�O�T'0
�#w����b�[�J�IX��S�0ކ���q�H����Ϯ���)k���'�%���(��(M$���Ω*���W���@���sWH�4��!�0U��%�j��)��/ډ}�a��ix�.��<��QI�-���V �����;�~���2ٞ�3�v� ^�U�9�Ț;6�Q�C`R�%B�J�8��Z��L&l�q|����9,����:�=��>��Y��	j߳�z��O���f�1��T���'Ӵ����ac��.��_@�=7����z0Q_4�!(P������GS�]�g)�\��V�>��ϏkJGm�i���+˽
ix��'�R�G-�-��U�� \��uCl��I����; ���Em+`Zk��߱�c�V���h
p	n��2N�x�>��`ۇ{/-R�]�SȲ����%�mQ�=���	ci>��d��Ó�%'����G�3���`�h"�Ӷ��R	�?	�:Ń�5�,����5�}�s����#{�RF����~ek������L]��������u|3,�� ���6t��H�;�W���1�d5O�^���0��2�K�r>���63� d�9ޥ�r�Co��32�w���ߟo����Ǐ��&X�O�B����Z?ф5���~��0�nD����,F���T)�B���A��NkJҥI��Uп=h��raf�ڋ{أ�xb�`��ݳ��NC��=���YQ���>0*��*�̥ôEhz}~,\�(��s�r�鉬Z����UR�w�MG{���r�l$)'��=3-��������ZhU��I^ǫ�����9Mf1�y���:���
Q�"��$�.���W7/�:���q����.R�`@\����ᇸk�ch�T�ի��C��˂�R�I&<�,�%@ZI>�^\b��?�T�����1.��Fy�C>Yea|<�j�E��o�	�����)j^	��oݹ�tr
����~J���н�?�~��v �m� zn���&sI%�:�Xlь�d6��?D3a���
�����S"jE6�S���1�"�2�Y{E@��Ͽw���;�wK>;/�P#��C[���qL�AB)~�8T=&��A�LT��)�ֆ�	뀞ƙ�_�4�-������W{�	1�z
��.*nN�����q@'�_΢<�-�0�ci ����Dՠc�M����3��˷�	|ĝIy<�{ZA��B^��^B�m?�iy��M�2dxpGʣ�'�l{�j�?ZN^%Sbv6�Za��>��-7�tb�!Q�{O�j���*]؁����i�"�й��}6$��$�
3�6R����NeȪ�~���{ˎ��n�W㱩���?j ���a4K�y�$K��(���k:���+��ͮѫ�{Ѡ!L�H�k2�3&��'dt�U����2����%���3z+�Z�F���?.�f���|<�혒�[�u�J��_���j�m��VL���M���
���C��4P�*MڼULpޑ��+�{?�TU�g'�Z_�1�ff��OӋ.t`��9����%�dd�*1�K�.��$�k�<���h�z}��Ŏ�G[��)
U��5�9l���Iͩ�/j��ѹPH:���E�%����u0e|�+)L�*��rn���C�6�w�,�P^y��#u�tQ\�N��:�bE=-��!��`��O�|K�xi��"ٟ����>ő~VK��<%�~ �ޡ1���$�Ddtنq{+�@�Mi�� j%�dPż�|���J�<�K|���	��U���,��q94A�L�]S���#�_L��:����5��G�.����<���F�
�-�Xeٞ���pP�no�w,����4t�\q� 
ۇo���K3��FoH�kǮ�x�E�Nod�Z!�^�4�p��N�<TH����`cOvȓ�R��\՝�.Ľ�����G����T�ˬϺw��o�{�i�ڊ���C��h+*$�w[���
�e�_���3*�}�e�U~n�/A �ޖ����Pڢ�?��L;�o�Y�R�ۇxgPX����<z+�T$1;E����)� �C5T���1�.�HY��GO��t;k�J��3ݥ�Ҿ�Fy��K�Z�`����_&.�ԅ!��!h�=7�Z��T1����M�ޡcfe;��w��|��:c�1ƠTu�����|��{���4�d4�?��Q�h����g����ۺ�'C���/�Ӗt��v����	W� L��c���Lig���e��D�<߀��q�ظkTk��0��t��K�h�ôՁ`'�]��%�c�j���������U�ZRAI/X�
&�XˡӮc�5��}A6g���K�uO~+�ŏ�n= �!<���k�{L����� �פ8�~&�do��������Bw��C��`����9	�.��۱����a
Ó+=���2c�g�j��ɐj���XrВ��3"�);g�+7dh���H�\�����4(�m����A��s�Be�`����<}��0 Y�^Q�����+�+�^! ���63��-9I��.��ń_o�_(��7��#�o�z���B"|2s'1ȍ}��B8���%�v5A����C: ��>O@�	��3��+C���Jy��KWWd���'_�IZ�i�Ml*5)II_z�"1tJ⮸_/���W��%�;L��)=Ф�df��#�iq?�Z&Z���a �]>���eV�k��F�lM�{��2�7Ç��w� S�"�v���x\e���ѷ�ԩ�,I5����xwY��1��'88�d����v]=(ҋ-�c�ϜȲ�g��Ev��~hd����ʗ��j� ?���������Qu���%��R	p9�7=X������S���ו����T��\���i��l�/Y�f���Ǻ?�ArQW�����m�D<�{*�;u0�H!D�O�qS�O�h��m����B��b6�&���EX�z�zM�����k�h��G�OR�B�W(�"LB%3qFk�xJ�A���+��g�MHc��jם�fVt8�.r׺���I��4��j�ع����,�iĖ��M��/i��e�]���q��ޛ6-ES�f~��ܛ.��O�*KwT��=�3a�@y�o�	�Wņ-s��d(F����֞�0��]�u��Dz�Y��U8��,�l)�*T� kK���x��lw{�ӹG���y����%�8�ȼ�?�g��X���:��l-޸���O�/�e  ���~0��cc��:�����֦t{,g)�#����d���F��_��l����j��[�l�69;�V;eqki��^~��{�I�N�%L��6��T�l�+��n�o�2\����=(,��X���439J�~����[<IF���l��s�z�/4$Q~?��$u��]����sZc�8��a���[3Cw��E.��Ϲi��8��[p��4�gE-2&v���,s�d�B6ئO<�~���&(��	 ��27�2ȸ���9g��_���6?Ϫ�N�k��=��7⤵�I��q�)DY<)��2:��=$Y��F4�$��J��>��">R���]�����߳!^/`�Όu��?fS�W�mm浟�!�_���Ɲ��r�(���꧚��Z+���C�ܖ�r�2���iQ�5�hO4
c�E��y4��)�-iҪF���� ��eA�yRR��4)�x0=Q��.(�\�6ޝ�|W�>zK~��z|1�Q 2�̎(�ǂ��Z���ý�.�>g�4i^O|f�f��,��s���Y6�y����kѠa�3�A��D���f�'\�,e����.(Z���WFWN��d �EE��B`������y��cރ�,98��DBܓ����g� C����$i:��D���45bY\Vέ�q�V�dġ�ąO��/Y�_��.�����&�V�|�zg��/�9v�P�=��>���ȑ%\��2��4���C}_����-H273�B�Q3Ά��D��LBt����6�6$��^ZVK�XbI��1�NX#��`d�­l.玻%�3�x�R�j��lo�>n.�U/�S�}NG�f{d@E�NDDΊQ��X���ԺH�����jX�hP�[�0UeG#%��mW���zt[`�nrl4�x/�O�%�	�7�o���w��Ma'�D;{�CA�(z�kԆj[Wq�\�Ѕ�ჰ�VF�L��o��2���@���4-�����t�0�x�^˽�z���Ϊ`hY��}v��Zl��{�Rѯ"n܀��=w��w�G���� �*�
it���` ��
���H���&���(M �bE#㖾B�x�1�J��Nѹ�:m�nn�R�2*���1��.O�%0h�('��B2:0�ײ�sύ/�y_�e
�]�;�.ooФ$0D��'�C�2Ԉ��)��5�k�9Ig!}gQ2��D��� �=�4�1���*Ϛ`�N��(:�g�6����G*�yLǼ�><yA�OCf�I!��=L]IY�y"��S�G���<�����t���l�㷒��I|Լ�4��'$_� ����T҃��,&h�+B;�o���$o���ir��k�V���O�Q�
��(�h��1c�ސ�����V���$hv I�s�(nY�m�o�N�磌�p���4��nl�z �~* ��@�� ��tj�\�	 ��r��������������g����d�yBqv�~�b�d:��n��I�\D��u��&��E(j&C�γ,3�.e����j�OI��ӳ�)o��rn���x�B��Ca���и.h��[�u1���W���̈́�e��V1I[k���,�e؅����-���}�!od_4�!@`�'<$nt�/yaS�4���gl.�����0���z��D�_J�V���0o��J�[�!�U�����(oV��:��?���!�@��c���%]�W�;����E���J?�V��	x�ˣ.ǐHg�gbb_T�T4�����>Z��l�\T'ɾqc��>�t��j

B�1fK�$A�188_�����M��h''6�f��n/B��ojKإhhȧ}��My�v����W��	�\{!c:qD��3"��3�:�d0������>�^��� ��P.���G���~Z�@��.��υ�=$Oԕ���F��5�Q>������d0�Ex����[M�}%���SۉT��q�s�D`��P�<7���,E�h��R��rˉ|�n��=�Ȁ�R��ȕ$I�/If���M'�$�����>��I�����.wP��Ľ4��R��44m���_=���7Nq���R��Kv�٪$rN�����}o�A3X�b�<Z�v��bw�]���ւ��,m�NQ��n
�V�j�;�.�$���~��.Os�R���I��dY����B^B�ߖ� ~���-h��\V>�Hɲ��
a����Gi���`1d�d։t������i^�3��Ez�=&��7R��:�����ui�����عf԰a�d���.�(Y�Pi_�CG�`��>��CTtrf!�;*���Zw���GwGO�V���ۏ2��H:.3E�(����n��Ȩz��$�ַ�U郬E��,g�׾:��8D�	f��ֻŊ�	�j�La�I�n���oŊ2�T��tD�QS��q���_;�5�N�g4���C�k]���"���/�)��W�;`g��s6��0����4SUw�qE���J�1 C��݉�/��`E���z �R�ه�!ɨ�y���7V7)-�S��j�X����8����-�HP>�ds���7�sY��3�vg��6p^��G�Yz:��^'��-!�g��}��d���7v�k���f�$se� 1�d���۝�dtGbJH@�k�y�D�1�?K�J�g�xOZ�YUVD�$@���t�L��n���c���9�z����w���]Hq�v^^*���;3[
�vSqy�(_��՜�*��v_�������-�/���3;��N)�&�P''����v-�Y�	�_Ju�3r^�65A7c1m��%Gsn�~,�Y[I�"�3���,=mBn����V��n.�T]`��K��۵����"q��ҳ�r�9�D�$=?�)VȊN�x�S\��V�B��/�Pp�sw�V��a��(XRj��
U�.��o��M��c2�O����d]IT%�e@����k�p�?�T�癔�R�n1/r�!��	cĪ�C'ƆD/ƋtM����n���ӫy����_��?�ZA� ��n|-��Q1ǴEQ�*v!oM�;O�E���2��⍺.���b~^�e}�i���OÞY�]-8�=˔:�k�p]�u&sϒ&]���*�H��<>��>��I9���Վڒȋ�h�P�1�(0�(�wW���W� �����!�;[P��~d�0|2�c%[��L�ȃ���Y֘�4��v�@ߛmu(=-��!�*�]ꐌ�a���|�֖�6\��rW*�L�r�����!����D�S"�g�e(�fuvUJь�#�=�*���⊓��A�J�h���:�ț-���ZX'�Fo3�� ���D�{�֣�M�>;���-W�O&i�1a��)D�+��� e���%O��>>����E���C�pB�TD1�N�v6�S�r��P�Y����C�IG�a�A��&�cwk5�%�""u����<S[.�o�����.sVtz��!�y���;l���ڨ�؉/�p��_�'�6�8���b��5y��qL��h��4���+
s��ɷПH���n�N�Q��b�����F{O1�I�aT|�Io����0Xݿ��p�>]f�>9�-q�����p�Pl����z��9&����>B4��N�WOy�2�}�'��ۄCp��B%�g��G@I�h;Ή����&>7�?"�lȕ���D���N	�Xe��^s�L�I���P���ж%��;b�\��(¥�ݠM)�v]8m�0��kRy(�DC��}�=0Ӧŷ1�w=��o�u�:�,�%:�M'��D�]��,�2ץ_d5ņ	��k��-� ~{�"�"����0k�n���q�	d�S8�����^�w�F�No+��������<�څ�&�@h�#���ރ���d����hR��TѨ:K���1k<�.���.���6!��j�cxZ~�x��57ě}��� �5�b/ˁ-OZ�8S׷�\�Pl�VH��W��j�t6���۫p�6٨�&�>���"�4�! �x� Z��C��!xoP�<��.��9xŋ��*s�D
��p-�W��}��?t�4o����#��*�[|�X��䖶c�&[�Ô��ŨY>�$�g�� ��2U}X�4^y&�)d�}���VW���{�K�X	�q��������v�_V�El���+�͌mIO��?M���G��h��`D}6�E�Rz�s�T۩&��j�h����
�Aj]r�\�\}�Ma9�m�#@�}g�.}L$)��u�j���t��w����%h�)�S�hA�ϥ�>'��5N�\���;/��)^���Y־1��Hլ>U�Х�dr��U��ש�R!0\֏�+!�|�dU����� ���6Y�n
V������6�'����o���^pv����A K�V�X�gN!:���:�H�G�mU���I�޼�e45F����'������r7�����:ʲ��%$��~�;�E.ו蒦�sd�_�M�t�x=4Ke$�㨢���踀���P�W�s�"!hF.L�K5��4{���3��{d'�г�U��ʏ���w�}�?j��3c�,��@T6�'�ǻ��LP�������;�D!iK� [H�)\��3G��n��2������IR���g�O��
?=��2!P�A^�Kz&࿓�any؞h�i�j�"�̢��Og:/�qlr���[_�u��D��������S��k�6pk�"Ln�v��[��|�Mgk󼓗�\�:��:C����!����V%(t���X�'ʪlPE�9rQ�vh#0\%�{ʀO<��3�C����<��蜂����z�<)<3E���?�����~���_��ZT�p[{��\���L.������-uH?��0b�#<���`���*GT��O�,����Ѭ�Y�V(��N��\��A���AG����O-SK�!����'��fC�2-3^-�`�Kƹ�51�%�%kИ(b�x�؊R�3+&yЄ�.h��2�Ēz@�@F���S�d���*	�4�.�����ek���@��7YV*R��3�̄����\E(���k�&(Bc;�D��T�R�`Д1Q��&�h>�?/~���;�Ƈ_fYX�N�'���0@�E�rX{�9�_�e&Օ.�3!g��Q�G�X���۫?�&E�����%|�!��Y�~;VI��W���@�{?��=��A�*��=��Zذ�ȭےC�X�?V�l�C�,ors@�402B�����9����t��l�G�1�Gv�L����(2@��<�ۻ[ ��X�p��Ǩ��JKc���L�ּ9|?��!�}ou�&O��cΏ0�Yϋ�qoI&��2��͹E����X�}�2�����ܨ�B�����MV�^4��b���|&��e��P�wSg|^��_�Y`�$�f��I�!c+#���e��{� �(Hm���u��wC�أt��qD��.*`�:5p˩�X�"���=�!�Pz����E&���b�ì��<h��B ��LE�!S��D#��`�/�[_�+�~Mz#�V��i�.�6fJtf��
z9<�,4�γ-eQ��3&�b�zf=�z�
��I�I�H�?VQ�F�
S�ǧ�{_���d��#?/�+�y���)���0�.��P�K�]}<�2X�l��W�Z�H��u���_9M�?�g���Ap"gh��y�/����`��.����[��fުl�cMJ׭j�t	 4�NKDɏEbf^@{���گ���v�jp��>6��y�֕3xJsGDky�5��[�Hϒ,-5_��1l�:�?}�V!d�K����'	!��]��1/��}�@+�^���o7�ܣ+ue�SZ۪�!�l�$��b��A��2A0�`�n�������g�E��|�S-#����X�X�3n�ӌ�����7y?4�8�D-Z�a}���$K������ S,�l�5�3�B�9�+�15I!�g��Mm�h�u�&�#�\��� �d�lzW=��g�o�K:�~�]�
��7���ʤ�YĚ_����B��S���2I�;�1��
���@oYR($��L:�ޯ�%l����|���b!��J|��Ki$��rrO�D�Ф��ǛT�W��}`E3B;J�<r��غ���њ�@��7��e��ւ����-��_Ĉ�P�="
@�8��*, ��+,?Gk�Cu�9��h(���|1����M�VTyH$isSo�D�r�|4��l ���?�A�sN��l�fl����O��<ZB���r��l�Y��G�T ��T
�w�3��Q�e�=-}�?������g�`x��_!��#��=H�+3d/u6�Q�D�r|���1Pٚ��sٗ��V�N����W<=`]�M頦�$��D2���.�����Ҡ�l
n^tv>����\":�B�G����N��:_R�R���n~r���M2��:���LN���X��-�n��	3�z8_�����)���&���(���E�n����sДv|�B_"%���4fBG��X΋ܫ�z��Κ�iЦ��旡;����ܣ�L��HM�')i���?WY,�J�ȁh:�����]�EDg <FP�
9RX�� ~�Z����F
Y?��jchLpp��o���Ps'*���N�D@T�ݛ��,o���ΒmI�~뿬�g�V��4�܀��ӻ.���M~���E�|ڳ}�r�N x@
E�M�V��X�gA�P&�*m���T��_�ZA�ȷ~�Ϲ�$��F&���X�Y� �. z/[ J�ص�[��U�%�Z��{�7���{iA�`����{�`^{�g[/�����4�cʰe��R��4��
n#"�NK#�QM�!ƏINU�]���
I��OgFK��9�K�6˗"�k�u�c#M`۬�&���X�kߦ@�ӁSƩ:Wd-�5P&l+_�S�Q`+��a�!���okKmF��&,[���F���̓��fǖʌ�9�||QE���������U�M'8е(���x��I�x\�V;�����N�*I\�z�O&q�ҚmcV�r<�om}���[(7v�G:������)�)
k�dv��9�5�6�E�r�]����=ȥ��F0�m��+�ja,ԝ��>���yv�άt����� OE�验��\����EӋ���/�/� đB����$������I��`9ɱ:{��bD�w@�y�]ɧY���Knǚ�\X�)���Sgi�5��ǟ��p��X&a_�m��KFg���1�����xOΟ����)����LAɕc�,_&�!����|[J�wھA��Љ�I@YĄ9�e����O�ϩR7M���E/�X�d�%��ç�����,�L���H�}+.�����W/�����،Ŏ���͗�
�r<ӳS .�ډ��\M�`�FAĘ����� 0�q��;�� �I��ɋ~�	s��������pc�(�������(p�9��Y�!u��N�Ӧ��J)R��z�w>��R���`q� P��O�A�3��OanB�ZY��[,�=��Kw�"�9�W�ȸ醰�_ֱ�l3A���)-y!$Q�g���Lo���.4׽n�5Fp��ZS)�6���\�6G�~ft���roߑ���y�m]��a�L1�o���xeR���;��>����9?���dС	u�0|	1L]����1�h]����r%�����	[�z�у��'��u�\��_ć��=u�Q�q��������j�f�K����4tͭjY3n����S�B���wMw��0�b�*��\LOt�����փ�Ӎ*�^m�s�o:�_ψ
�Dd���7��B23=7�i<�Ob݁�:�����,X��1�Fx���l�=X���� ~U׵X�V��͋��U�{Ճ�׀�j���d'#R� �{�*w"w	o;ʋ����It��N���d ��a=;��!�#��_���q'Ė&0"��>ć)�exp�bڿ^k���>��D�Ĩ߹���{�����8@�RhY��7���Υ��@��U,!C�:ef%����Bev�izkiB8(/���M��IPv�]}*������vl�t2�T��7��M�5����G�3Ƿ��{�b17yM�+���dӶ���}/�fH,�ӎ8�Qr®)����SB2.���yƹ�+��O9�`��e�"���̊1�d�a���	���"�����/͒Suw����v�BY	�E�������vv�
>��ͻ�-�I�e��\����gb�(�3?_�aH�I����!W;n�w�a<���S�FƌmZT~�����ވ�r��^H���a�?��y��<�&���䮪���z��i+c��x��3�%E٢�!
��N���w4�Λ����^udp�ʳ�a
��˹��zɪ�����U8�F$pwUa���z�O�!���:d�$�8t�)QU�$���hE��I�^� s1�x�+���f83�\����X��*��G���Ӱ!Y?��j���X��s=[ʫtak�����5��!"�G�\�-�'��l���Ѫz8ȗq���Y��ē��S�*;dE��DJsR��NJ}hvHd�@}%�}�2ϧP�3�25���'�Gqڃ��~��a�?3�C�!q�b%G��ZՅ0�[K=�\���ԓ�B۩���"��Z�����|Yܻ���^?�}��	�i8xŁ���[MR�P!��EP�]bi�Z�v�uMI�ʱ��@�j��c���퓫"��>�8�&P~��r�c���?V2r��~Ǌ�����'�A�^\�E[Ɵ�V>U���7HMj���>�&�b�+q���;�K�ݕ�E�i���rP[;P�f���j�"�7��h�.˿k�]d�Kw�x��~g�D�^����s��b�5�I�#��ފ:�򃘶�i��Niء�S��������=64S|���|��*՞����ʇ�y�IbI����u!e��.;O����j��ui�Oއå�	�u�ݮ��>�aXc H�_���_�z���t$���Q���,���bn8�T���$E-���ܬ.]{TO�r
���U�^-�j�Iٟ���}"����0) ���D�3��N��1M#��qPdZj��၇��SR�E��:�Z�%�Tb�T�~k�`ԠpIHu�l����TA�֟v��bd�l��!��^�`g_��F��_߯���a:lO���
�N���':&κ��Vc�k�]���,5&��Z*OK��,&��ui�(2Ӎ��J��٬Y�HX}C�U�RO]]tW��5�)��9��k@9�Iϗ��q��ɇ}���������}<�#>�wx��Ǚ�]%�c;Y6��)�l��EtD��>?F��9H=!k�*�Lu�r6�!J&�n��gb�U}=	��B}R05����β�����gp���Bn��r}C��z�s6�|Ds@�]fKV%nW�hM�t�@���0� ��);y'�zN��61��OPQAg�,�ЬWQ	�߀V�ҝ=��a�p��g4�e�D�O��L�/M���j5��bĴک�!���T99rv�y�;��I��.�L�n�HF�Ng+<v=��z*9���M�:i��!7�e~ب����_�L�@��΂�M�ڿ����b�M��}#j��>(�Ę-(��.�V	G^Ṉ̌Mb
UZ։T�{��⭞�cHĕ���*��������E���\�Q��1	�)���Sє|!�?�������L%�:M���ewc)Z���QfПߝ+��Q��'16�}�����-�G���Z�CL�Hz}��b�pF�0(��w-f 9�Cn���f���P(,�{�z0��͙�3��.&��-k�UV�;X��fDq[�j%�{l��̵�/TO�@��QJ'Tg`o�Ԍ�WCm 1���A������B�N�����T�+5�Ɨ鎾ll����\�Z���6�J%���$�5�B�1��3�Q��a� �>0) t��loy��G�{�N��)�D�K/�L3Iß�����=d��'���߂:��(��m��wb���%��]3H+â���U-��/4�C�j�$0'(B)5����2�;�1���Q1��le�(�t 1fe[�kU�#O������+�ʯÝٵx�����Ii���1���*I�|�\-��5�b�a����f����ѥ����~y��0],�a����9@�>d!�:�^p���ʧk��/��"L��a�H{�J�h�}�%���D�J����Ķct9\��t��DZ[�)�z�E'I��AJ�p��~�ѻ�SW'|�f�G�Eѝa�4�@e~m��og�'0�3����1���6зw�j,�v4	� /�P��!��xy1�hY�j}�骗+R�k�����ĸ�N����|��n%�m]�y��n�^�� �LJ�%!`��R.�@�I�C�j�H�qGU�2��6�g3ߏ<���,8N���Y.!lCq
Vµ)د������76�����A����љ6���J�Ud�C��[������t���LS䞧�{rK�ωa���ÿQ+�x�T:
o�}�Mj��;��� ,��(�Ŀd:��I	!w:i�Vd��[����>Ųm;��w���?zuI�zqhUC���7β�%�����;I"4lY�od�	��b��HodEqW�E�i�<�-0]�]N��a	�r��1�P�BE�R��؅����j�"4!z� �����^!������D'�ʱ�h�K�A@q:�N�ס�g�[���9$��((����ꋼ�6�A&	޿���Qh	P��C_� ��d�5*�-��Vh��	,�� �A�U�r���=��#�*X�(N�/(`\;���;�����ѡ���xY3�Gd}���M�������������Q㨍J�x��ׁ�J��y�͑��kl����D�K�q�~q_�·�����O���Ջ}nc�*�b��(�e�S�_����rIs����~�o�ޢW"�m��
��3ې��QZ�����*6W�.�E����aVY)�j��+���BBH��N�S��C&��6q��r4,�D��< qkFP~n�.>�d}dg�'�?g��ԟ��GȬ�'����6��|olY���l���>��ʭR�F<�W��$z��{=l� �/��DW�w�ԑ���D���l5���緖�da*��@��1z�ǽ*�b*�"��f�|ӓ�i�y��=e����9�cPohG�߈��;��6�����q��+c�P1�?��󷍔\�g��}|9���eH&��v���,���ׯ���<Ft������ՌcvQ��QA0%]��~�x��Em~�8��j�˲p����#��,?�9����@�]YkS��ˊ^��}��{�	}���%f=�R��g��h����$3pcd�)�ҌhQ�*����������<V憧�95�j`����7t�g���L^��5I�WXih2������@z?��}��^KYM�H�[7�O��o¯b��*�ɲ���A!���p��0K�L���S%��V���q��[58y�>���S)�U�R�u��<1��VJ{(���eh ���E��5��%l�S�+�lѤ���LHet�%��x��X�s.y$5�>��Ž�5$���J
�A�e���罓L�=s�ĩL�� Ri2�f�2��s��v��{V������}4��D�Ī��v��=O7�I�o�I;<(>e����這ZFI�*�D̓z}�4��Q��9����>"�F/���5P�ml� ��%F�r'�1o�:fZ1\�.���	��k�z6��-3���e��-=@u0>���og8?�G��(�5��L��۷�n v�ȴCb�gJ߄A�ng9=gj�nC�X�VV��D���\s�+
�$�T�K7<FO��<ҫ*���Y�Q7�>>�'��8��X;$k�l�0C�ɼ:@��]+�'6^wu&�+*u�t�@<�d���5��PnCTw�`��'}h�!�*�<4/tL�u����㧕���񏹥.(��hPrܢ|Ui�p@8\9?�P3�_σ<H�į ��db���L�����2�D^�n �t���KlL�OQ��z�8cu�TKKl�oάR�I_j��SH�P�4�ݖ=��8�Β<ǲxd�by<��g�H��Z�<���_'��*���b�j��M��e|ץ��<A%؅���-ց2,PN?�F�\з��h�[���fB����0�M�tp5��R|��&Q!���m_ET����c��&-U9�A�B��G��W�A�FH=O�j��MIq��@Coiz�ty���%�wx�9a'�:�0Օ"�k�1IuɂH@��l�%'ك�����/��͹P�H��]�wkWqCǏ 9��ߘ)}-D�����6���.��T"��X*GH�<^���t�o�aE��c�6HJ��D;䆻�r)	98�<��v0��1�T��0y��9w}�)b0
�%�;HI+��R���Ե^W|ݕ��9��%S�⿬k�"�+C��F3T��ۃ�;7쨃4�d�
�V[�6'-�i���Kyw����Qc�[`��E��aKF��1��#�\��i�N�>I��i�����)!'�4֩����\o�o�9T�K]!_�����\7�ʅ�;L�A�l���cx��=f��Ʊ���t$w�r��j�^�W ���/fņޮ*VB/����\6#�s�ʝ�q��F���=}�'U@��%`�]7��ax������c���5��}*;�ָ���5�R	ɔ^[j�Y�����=
/±>nͿ�g��ۉ�GVF��yup�B�Q�3�(�	�<�������Ph L/��FofC>u״;�4O.�e�,���ף.��ʙ�AI�j+�vB�+�K�՚Ή����<���� ��W���� az����Z���L8�pLZtNŢi�Ǝ�t�P����C0jSE���Aß�e%4t�z���B!���T���LzPO�a�؆���pC�6ȗ����}�n/�h��;8���R�5w �������y)����S�4�C��������oA-�X���?<�S�]
z1r�ZxH@��������t�8�m^1�����4�#���X���������B��L��?e%�.��W�ѧ�-%"��n*�VF=�j�
E�d�O˛[��"s��#S�d�F�+��T������.��}�p%���'ئT?~ν�RR�$!G��X$@��V�#����;��h�QF�縳�e�bʷ��Rp���cuQ����؎����� ]��`��m�ރ��?x0Eۂ��Z�,���,�3�����8��qI��Nã��I�.�lY��߾��A4�ram�g���e�v���@Q�o�#��J�S��">�y.� 6�^y`�񻔛�F#и��S*�ʴ&�s�H�2��ݍ'�Q��A^���U�4�E��|��=��J��*I<�V�"�r_��qpYg?��ص�� �1���;�7�?D��;����⯯g&̓q9.c�(����7�(�O�S��v;g�
b�Jۨ�mtu	�)F@J`�$rw i��.�Ci�4�����}ӛts�)����^'�S���r:,�/3g)��S�8̎W����X�V����p|G:+��%!�K�n�-�D��\S)��"�(���&g�T�6ߛK���\�ʢ���SBD`��_{�-�ӄ(R��Iy�[?�#��?��G�$4Q �A{tՕ>�� �lx��q�(r I�<�4W���_�X��e:g�H�pGk��q9~��\����(*C���sA��_���P�gj/�(&/��U�f��J�CT�;to2\ �*Z��Ja�/!@4S:��뀜�L,�H.pXdm(3jz��ˋ\�]
�9��c4:ڞ�.���Iߧ����1국+uU�1��$����Fk�Qn��HC�c5��@�쯴G�{VPI��s�
fydT)Q�0M/1jo
��ݗ��rPe�Z�&�'��Xګi�������pws����g�g�g�_@�����W@eH�߰�Vj����Ai��]�;x�� ����7Z��@歊%��5~M�����7}9��4_,m�Ȳ��g{���ftk@�D�o��5<�y��
�/���E�(�E?��6_i*�!#)��!��U�L���_֋i�SߕS|�݇p���`�UR�	�|����U�����3�9�)u�<\�o�t�Sn��szGPN�L�Cl<�b)�6���r��'y�cX�ng� �Ee�k�\���p����u�{`e��H��&�} M��#ɏ���d���(����!�Ts�J���U�=D�^X��"S�H��i�`d�/	���3m�"+�m��!/S��Ӡ���H�1�ߒ`� .e��/r[�mБ�KCe���C��U��t�{���OP	#�y��v���M�Uv��6R$�Uv��5b� ;U���4=R��FNE�f(��Y��k)'@���|�|<V��Ή&)��4�D$FG@4:��ǹ?���M$�c
RWE\��咅1tժ���Å*�s�w���3^�@
����	�!�c�r�Iѱ2g�����8H伾��|5�u�o�``3�`�U
[��<�Q`���<ڝ���r����A���]AxP�g�[�d���m�b���]���K�uI����5g+�ZV�m�=Rb�rͥ�p���~�䫷����sƅ��_-	s����n!Z)�vZ�	�?⡉�b�U`QM��Cg��bu�ϱ̀][�!h�+ 	�n|�V�ŏ�x4��� �/��\�A�Xd����\�A�&˨������*�n��-�s	��ii�nđ�g�p%��)W:+�zQ�̱�Z���k $����a-d�f����e9�J�N�ݡ�K�5K[sK4+>s��g�)M��i���;�����=v�������b��XH}���ʟ�g��H�����<�I�;3P
�7�7�0���WQE�zv�$A�%�����+-���@�ƨ�����Y��@�;�5}-�[D#fE�w�#�w>�y��3G:��������=b�$�~�ˁw���1o/������$��uֹ�U��M2�s�٘�RDv-
7����W�=x�� L�oU���Hy����Ki�����r���#{նֱ��l��cĴ7�D����7e��@on�<���H��u������gXUKg�"/����;Ȭ�F��I��qO|��l@���Ŵ�W�΍�8t �뷊�r$�v�.�Hė��q��_L���ώ���v����zT��0�m7�����b-*���hvc�y ��Ö 4�3���w5�4㚆z�"�s�T����qy�|=�eG��&q^:�v��"��w=�G��H�ĵ�^�)�'���V,	7U�r�Ľ��͡��N_������<��=l������K��F˹
:�YtV���|a�8�0T���W~�%%�F��k�\��2 ��}���3�3X�f�U�S6/�D�R����y���#���������0b��q1����e>����PF��c���ހj����������������/�����{0X�^EՖ��v�$.��˛��b��/�
���Xs�!���A�#�<�:�Ik�ힼ����p�ձ�!���1Y�n}��#]�iE�j���q_��B� @m�ѴUd�����z�5��Nj�vQy�X�8V)հ��e��^�n��K���7I�c}G�*�񊾪��V�_^%9�d���0�s1[�B�폑XR׻�K�Z�B���
m�WI�~�)D���٘&.l1-�,I�W����pp�K�u�s|� �I0��b:Լ����С:���/-"&p��!�v_�v�Rޢn;D����0ʮjj���\
kGW��#yMտHa��D�ѣ)���)A\|(�5�#_��C�E�Xls*���:S�K�o��n���.�w,�iߧ�i�XZ��:��ʃ���Dt��K�� �T j*��;�$��TX
�Cf������?��O�I�~җ]�3E �W��ݹ���ր����������rv.M�瀻ݘt�I�ں.X��	S��Yz�3�تO���s�6���#���$��O[�"�-�S����O%�2c��e_���P� `�z'��!q��	�p�F��@�
��n�8eS�+ ��N��m�W�3�V���x[֒i)>�J壇�w�!5u����&0\)I��q�k�	L=k	e<�ΆiZ
��Ts��>�W�������v���CL3������s�θ%P��� ���@�"W��2�-�ʇ�<��`�[��)�U�~��b����;ݧ��Eb]�3D��,�S��H41�8�Q�'m�~��?���Z���1��rr��<yh�4w5|�Tu�	�S�!����IA�|q[�?�=1/���}EH33�G�7���,n���8" ��áң��\��Z���OCu��m˺{T�~
U��x���p��rD��2��u�s�!`R�<ҷ��Yaڄ�O��u�����9.��g07)4<��؇SRg�Ɖ�raS����2��~ȋ��؍b�I����ģ&�T YXRw^l4c&�q+1�ka�,���w�g������L�7{d�4�%��A
ޖ�5"��yc���	��\l֎���������nk�W�R�F�SE���l
�׹',ɫ�-`!����1-meu���*6�Υ&�CԌ����)b�'#��o8�.LR���C�A�yV�w}\j��Ŵ.������D}3�X𾰝��sC�3�$ߘ>�A�{v_+feHEw��p�&ojY��!#Pqݚ��to��e�Q̸��A	L�}v��� `Ut�q����E#����X`����P40��P}ek��ɍ�O������+Z���~ָEK�(��D�Lg����[�KQ��ֺ_�{f�F4�H�n��FTt��6D-߰�g���9�;�l�X#=�8���p��L	��7أ��cݽ��v�&�A�4_���X1Rr��!��%�SK�����T[y�;���x�W��PM>� ����@��6��%2��/8�f �F���l6F�;g��e�8WP���ɏX�#<d�HnS'TvP�,�՟X.@X�F��a�����Rk�I��G�igc|l݀��oy�\4�9Ӓ)>��6�O�U��9!�׻��F�[�!}����@��9h-vn%��i@��J�E�BN~��g���4%uO��x0D.;�U�K��ې�8��8:�p�U�,�|��ܨ�oSKX�*)s4q ��r�m��Il�x R
x����v���
e�j-��9�OP���k����kJ��gI�21���,D��Qg�Qx\�&2`�I���q�
��'�TZp>ڜo�:(4H8���n��L�B�Bd�7���9�D3H��m/��vjgl����A2f��c�� ~q�����B.�U��k�o������@.M���0���t��mmh���0�}�׵?a	v3SA��r��^ Q�U�ۨ��T!h�X�Tf\�nj Gs,_3�ϟIufy��z=qdep_Db�nn��9��K�}��Z��F�*�؇�c8g�	f��"����V��q���Z�ΚW9lr+1��C���S��9p��ҧ�4~&?�-��G�t�M��N%/Cv�#�YKiRH���,C�$�������5@��Hϸ���>�)BF�Z��\�����a	�-ݱ�s��6�T�Â���
�	W�e�m�lkJ%`	�	�����<Ew	eB�0$N�K��I8���i�d9Q[��x:�m��u@0�����~$=�5+�{����Krf��T�b,��'{����'T�_s,������p�Of�s�a��"bC�;h�/���gVw����a���d[��� ���]���Ku����X"�f��~IV��>�.�d��:0�<�I|HEdxS
.��q�3K2V%~��FF�$�~�����2�H)M�����EE.����qli��I�	
Ѭ���
f�9�<�-���+.7��H6���{�i�jx��V\���
`y�,�7L��Y�K|�$��N�,:ijmvr���u#��>v�i`MT��	������`0�M��1�2�<��/��Tt`�̔���2�E�a��Y�]-��{!e,b���=3�j3�dG�P��Mu��� ��$,��F@����	
N��Ԑ�i�����+���>Ho�8<pS���!u	���8�4vX���UF�Ol8�V�_�>���h��-�Vh���z}#v�!�|�i�QQy���N͌y�`	.��o�c�Ö-�R����y���Z�n꿔:�cĤ��H��E?�	&p����f ����`��P�2os�� <�-�W���t��˚w̻Hx��! �@��18���Ǜ��";ښ��`Hy��Q�1��}m��(�$%�)�[ɀ�S�\��>�ZI��V���6z�X��0�<���������kŐj�c+5�,.�_�U�5��I��`O}̄�e}�-��PG4�׏^ -F�,�N�9�������m�������#;th���<*�&Y������o�����@@svgJo���	Z�}�Y��Ɵ�b���Nl{��i����X�g��HV@�@�W|H&U�|��A��X]��nA�w�u	����i�
�<1̣?=�j�:λ�n�L ��W�C
e]������ͣ�x�����*�t��~0
���#��g��� �;�e�/�ټ+C��_� r�R��!�ee�q�q%r�9���;ԡTz��	ױ��B�'��Y$^s�Q+?�7��y���E"po��9��~��tڬ�v`3��6�zM���ip��D={���t[^󠓺��4��IU���F������Gek{o�X�o��?%��eU*]Ԙ�#��.lm�.�#���C���\z�l�������X'����Q �O�0EU`*��es��.7��Y+�~���Q�f�����i�o�G3� �����GW����$���N���r;&��VN�U~�5ҔF�u��o1(y��c��5Wt-��C]���g29��b��0��U���rQ��f�er�-^z��v���Ԁ�0�*3a��/^+�_J�%�P�+_�5�-��� �v5�%�\'zO6�1X{L�3�n��HAc�I	���zg�?�*�:7��֦�,��ͦJ,h������? q�`|"����(���>��NE�5����!���	�8	�ĥ:<��t�[�����9V+�]B=�hL��h�*�c�n��[��'��f3~�����\'�����/�?R~|�`q����u@o��`�)v"�\#�G�l���	��%�u�,g�c����?�`�m~|�A��)]d���}K�s�}�Y^^���6}B)P"�!w��ehP���ʡ��	�6�"����`+qz�k�j
[�~Y�]A1F�>g�=���;/Β^�)���?&����)Y�T�q%���G�"0V�8��wc�!��^�t���u�4썇���ߗ��^ܜ~��ȖSV��#F���x>�~L�EI��t���+��T�:�WFP�Wu�+E+��ˍ�jՠ6�-<C�H+��� ]�=����$h��>m��#\@c��f����ϊ����ק���F�7��U�@�Rxk��J��c�19��o8���=mt�%rDU�f�?���Ʀ]�r"���dO:^�#[�̈́�}�*v��:���y����\�<��Ђ^،p�m��9B� @�w+�Y6��khJ���J����I=|L�ƫ���+��+����hb���Z��qٯ<IN[ �tL�����r�9�^¸���T���cN �MG?����a��ԯYu���6�{բ����_"����$�������t��[�QLv��\dyh�	�0��ԓr�,z8@?-7���T���q{xNݮ7�B���j�bid
���c�������G����%T�<�w�s�1��:�®p\�yOk��)��I~���?B��������"����AiŒ5�j�,U�`�	��:�&=�e���M:�'�mz��7��>Ҟ&�Ɖ6�0?�$�������M����c�9�Ύh!sSB�w�W��&�Vj=�-�X����]tt���k� �;�es���^O��1Hx���ӂ���PhӖΗdC��r�hFm�g��4�A�ֺ��ha�J`܉G1�ß��ă۠w���N2Tw^I˰Q�ﻬ:��g��O��g��ɲ���r���xG���TK��rHNG���4����b���L(s��Q��l�I�`a�� ���*`��U��*n<@TB;�
2J��ID�2$��)�;^ɰ�,)�v	�.���҅���Ղ���ڽ�)\��`2L �^:��dY"��l�;dO{�R݅�߶pi��8�I����Y�J��k�7CLVF�G���ϒ6Ƚd�P�|��<ha��<u��u7X��hǐ�����_��:Kf�n��^�.}9�P:/�|�no��������nU/��=~��R:��,�d+��$H���i�+�0���C��zp$�nu�$����QG����}��������O�Y���\wo���j�x����j�u�6 V|/���������$�h��`�5�%��NT*��U��Y�G@�a|X��J�E=�u�sb��}���]�{;6����ȧ���b �`Fe^3«�TC*���Q���p��#l4��e-��S��E������m,~���!DR9����n2�ˢ�F|z���4>[~#�.��P��N�Z����Za*�BGݢ��y���L���z�n,�k_�D�	S�*n��8�K�׵U �W��a����Q�h7�*��U�ML;H����ȟ�g�����tb
��܁�[<��l&����E��#z���)�����N"H΁Vu��7|1:\��ҹ�v��^����F��U�ǐb����|�v~XZ
�Z�ড়�,Sf0	lnv��.�3�O}CC^2<wh��.�#�F6tItP��,��:�k �~t���8��jb&�������W�m���^ɪ�	h��d�^9�L�F׍U��ɓ�7�K�{)���6D�:P�>�l��'�گRP
7|��2p�(t�2�lc�b��&ɲ�>�s����Aٙ�Ha\xCȊ�����lz�H�Ę9�M�V;���x���t����e�4����8e��/��b�N��Lv��53~;�|�x�8b��=(u��O� ���w����T�{�d+��T9����0���x�;�����T��-��̝Q�GLjo\��v,=I�⟤B�$�G�<إ1Eb�rWI7���6��=
�s`6V���6ӤC�D��[���p�������F7�s���W�4*I�5�s��x1�����Jƥ�,Fx���0��9q��#���&�(�v�ȣ��o|�c��j�J
E��Fr��7�C��x	���{�vP$�u���wj;����/eC^B�o%�{�R��XĤ7*�Dg�+�/@���\n�4��Q��J����1�񊗴/*s�M��֬�#���d4�X�� �o<vw���c��tV[;��sg�q|�:����f+�Ml\��'ls ^�sq�'<eM���\�~��N��3jâ���{����~�a��eh��Ǽ�2�xja-�ʢSV��b�m�d,�m���c!*��<�ҁ�$X�W��E�ϟObGxP�K�3R�V�pӘ%P4��H�WאL�_ҏ����yن��a���u�-%Z~�t�*�q.�
����孖S�6�s�-�8J���T^T��;cN�Ϟ�����;����c媋�iz��D�.���|3fu$��P�?	aX����=��3�ۏm�r I�	JNf&u)���ʡ���� �1�6s�`1��D����� 7y����[ O��񓍨%�}�������*��y}��J����e��f`bz($��>W{?�I�ڞ,����W��A��Ǫ�d&S:�9�}�Z0;�����&��7y��?@��N��ju5��D2�&H���EB!R�ԧ�+~5�-+n'G|��<3oJ��a8-C*���Ҧ��R�	��I�!�s�X:.z�B��.d�)��$"��/���>������0`�ڒ�r�r���G�sW�zV��n�/,T��A��&�{O`�͌�P���[��[{o��*6���ɶj��Rl�ˢ�?�[.��b��-�t��"�޽P]7p�$ zz���y�y����P&�$N��CK8o{*�NF�,�<5���n���:C���GFh_B�PY=�m���":��6V+�
0��	>V��_�?�?w �yª�kH'��οI,�Ɩ�n<�����Y2���ejpPޒg�s�p$~.d#��	�qS�T45	��α��&����sC��x��*tћ�v9�f��x��ǝho(���mK�P���|�e�`��*ֵZbq�K���n��_b�L��2_�:�,,�d��`t��9Fd�w���)��U��5(r���2{?�	�.��i�[cke���� ��b���)��ϵ�Kqe��d멍�]�}�n�LK�x��T���χ`?B�$���<�%$q)pKwk���8�3]?n�z�q��U[��kz��A)�~XY9�S����%\�=<��>�*(v��cNX�*��9�)�
y �o�*P�"�B�p�"@	2���4Qh��������q�O�_�l݈DJ(�-���:����;�P��Ay�^+�=|���U79����-a�b��w�k�����y3���̈Eո�Xگ�ZD�s#u�̦t`��Փ���'�PZ(�H'�K��1�'�%�>`7�^�N�&�p�����72h��r�Fn�gJH�ց��O<����u�b�r.wG�y#�;����q���z��r&ݑ-��U�ͩt���s)xk��ǉ��I�:��t���l����k��5�
�v�Fj{���T�vv`Z?��E�'3
��[\�zL����C�ɞ��Y)L�k�������	��
A��ى��{1��6Bx �\̑x0]��x[	a=��=)�A&RX�S�4���V'���c?�q'q�􏛔[`1��?����=U%�7A�Iu���t�x���n
��u�Et�f�p���h�zaX=uKߔ��X{�\0�4����-SGZ��G��J<��ϧM�O��\�'Q)�^�AU����F@�?@&I�c���&SՁ�HN��:��8���s*�����:Ŗ�Kת�g-wh�rbf?�J��_��XZm!��ӆ�Cز�N��e��U�U��9��}�F:Y�fH���4/2!%Ŕ����V�	�=�Q�
_���<k��k�|Ȍ�Me���U��T�tc����2E�,�)��ӱ��[&>��W��ʸ,�ϑ�J���C�/*��k�	��GT�}|������9w�E�f_�^
��u��[M��C�`+�.λ�1%�$&��i�h�8�F�',��C�䃺õ7��[��~�=WE��V���E�� @}���n~��1�4�URA1�j5��ƝP�kou"vK�{�]mn��8O�^D���U�����Iݘ4����~�;N���h���d�o��e�~�qQ+X']�v��P�5(w�O�Є�~���@LŞ�<m��(����j���qMgl�'�J����%gU��!�\�\�jdP�a��v(v��{�Ze]�Tͅ�dy'A�c�,i-.��R�*�n����`�����IgL.���C1��5�Զ2��YwP�8��p��)�?`{+L�Ʀ:��U�+B�Gz,�[�yNu�B�������&���-��C�}�?y3�F^:��a���Dj���hdoJ�Ǐ��}�יí0�k:$�ޚ+�QVډ�U
��⌌Qʑ�gJ"�5j@u��!�Ot���Y#��+�ւ[�"2h7��U��E7	���W���f���P[�k%R���~:��W�"��	-P�¢.��U����ro�}@�$�dh,AN�x9s�c#�{��w�o����gi���ى�5��8��µ��1D��]��
��I�T�Gi�O�KQ����~ �i�!��9�##oU�J��T;$ƔH����m�j����hR��FT�"\�G	�!7�r�6�DWH���ŉ��4�hP{?0"QX �%����N� �jnv�n�ގ"��`�̟ѸlǾ�3����B��	�}Zٓ�`���B���C�_
C���j��<9�U�T_��	��o�]·/��j����nq|><|����`=��	f������e�Ue��<�MV��P�KN6�N��Y�4qiXnO���֌R�Z��fX.��>��*�,S��_��*}(�U�N�V'�E�~v'�]*�����\{sJ���l�l��6F�Ŕ�G��~Ӯ�wЊ�Z�ٱ�S���{q,�u�}��o[�`5i��>M+ t��gK�Y��D��v0S�B�{w�¿iQ��Z��_q;Σ	�P�ƽHX[U~���=v�ՅĴR���z�O $/����f7��@�\T�5�v_�Sg���S�L-G)W�h?�.zk{�Vg�T��@1��̞��ڼ'���hX�J��D�R0��L_���j��AP��Z����Ì P�3�o��JˑiY E�c��Z=��9xt���7�e�"�ٲ�� ;���.��W5�`�1F�/������[S��`�W-*Rw>��զ+�X���=���E�o@@� �H������_B>��y=�.$���淿E�q��s�B�K|J������ ϫ��W�\���ߧɽX�bf�і��!����C�;C���ʵ����r���z;G��3˓T�90�
�^7q��ADVNv�YQkg	�	�B7-p�^�B86=Pe��������G�;���lȀM.�yz׶�J]DN}��P~��q�ĪͰ�����x�#$��r�=�듣2_ -\�`Q�V���P��;,!�!���N���;�xx��{ѕ�;n,�{_���n��������~��c���|^���'A��'�m/4�ԥ㹊3t�J���*�����5����r�b� ���B:Ob]R�n��>��Y����Aa
�.Ti�*�,�"�Vhӳ�����x������A~g�!�@;2�NP�.��"m!Y��&���G�����'�Z��0������|��'�	���3w�-�'L��H��}4Jk��sҩ7��}�VG�ۭV8:0��2���d��������+��DRZmZ"/e�\$X1$`	���V�A����?�<��3�:�̠�9��-��~�ĭF����d�4����E�M �)���G�iw��lE0&k�Q�)����K����6��$P���ρO�ȧbX*:X�ú(&�y��>�&�'>���h��(��ԕsE�����o:	}e��Z�_�:�������-=;j�����|���0<0��h(�fұ�1��ktϪ,%�u+j>�5�����xUvn��2�S1M�������	H^5��B��Sb�< G�E{ s�,Kr!��N��%�+!����1+=5;��E�q�=C�� "��z���3a�^F�vX��SX2:��69XA�`�t�cʑ���,��D�a���M��EZ��s�:Y�$W�Hp��촔�h��؎�޻Y��ƽ��(�� �p�����}�+�+e.OF�ZDS�.������L2E���a_�T~��8�iN������8W'���!*�_��
� iޔU��n2�	��R,��"ת	Q6���2�~������P,p�N�2 �}��ؚM���}�(�v�P�������9( �,^볃p������ӯD�T�TdC<�S������������r�|��ϫ� �{�����z�ʛ�$\�>ه�Ɯ5����e�����"��@v)~��܀�3�s�r|
�|�2F�L⛀�q�@�tӼ�F���/���������l6���"4_f��4�.��j�u������qR~�B$��b=����31��������"E�Uf��6���@���q����5.~Qz�žT�-l���b)'�� ����a��S�:�$�5�	��r(H*��1不���(�w� ��=���/Z�4.%}].��w�ґ�ô�73:���@#C�; �������}�i [��悙c���Q�3�������_S�ai��V���Tn�wXx��оzA���L��/2"��TDe�09�ݏ�ti���R�Ę1q�[�ȭ�����*��Ea�J����¶���� (}*S�G��f�����ؿ7���Ĩ-b� ���?��&2p؜|O�2H�
p\%�_���A�1g�LX��n�RM޷�ǛD�$N�Q��,���ۯ9�N{�"ȝ��u�k�\����������
cQ��l��/�o���Zf[�`��CN�Y������c�C� h�#�&!:�Cw�\}t��M̔�D��5^#
$c�'����]�8�`\��������l��~���,�G�F�E��[�?�7�.C0'5^��Ĥ��k��+�E�?FH������TS������hhh�Ͳ�
�w)z�Y�|��<�<n�3D����&�=`ڂ��A�6���-��MQ��B�W�-���)�a%w����_����Uʚޫ� ��RJzc�|�.L�_[+:�S�<t@T2>��f�Du�pz?د仾�1P��R`���,��=�{֪���D�8@b�E�*����lDՑ5@���i�C��`|p.n�q�l6������?��b�B����p�ͤ��n��̈��.�8�,���)���~� ��)L���j�Tc\͕�����[&Ꮍ�{�	ײc�U��%X~��ۊ�3v!w9f	Тb��p����Y��J�2��җv4��ֈ��9|hH�u��~H��x�멷��Y;HH�|�����.��!�@J�e"�`L&�澲M�!Q@IՉ�Ӵ\2�ػ�����CO�s�.)�����<��H��$���]��mܛ��n}ݚ�NK
9O<�a{�);OF�����ss�+��Q��=��ť�5�"O�s�A�W�t����:�[}�|2�߶� g���bU9��%q�7ځ2 �}�����L4�))S1T��t�����~%۬�G�}GȪ�w�t�������U�4I����7>/j'������� �?��%��s�3�����߀�HE��%���9P���GqJ�7G��������݀��/�H�}��W��(�FS��k�aw���ȸ�7TfT�'A ⦑`�u$�[i�NoH���:K�nb�j��\>�=�s���N�$���#j�9~
�`�O����yb}rǋ�>����`&:���`;�u��f�1̂�eb�*�EY6 Ҏf/2�����fX�M(/"?�@�F�&(�$�!f���4-~lc�FI��P�_�k���w�� ����h�0�Q������J�s���H��F����N�F�[j�)��k��aÁ�+���Z���8�B�γ��ܯ�!���B��Y��ӈ������j�P��ϽRN�fv"ɍe��I������G�e�){�?J#��dZ���KJD�wF�����J��m��w��ܤv-"����w%a �mJ�r�Okd�R�~�ҶXd���wc���j��foE%��I|�l�z}�D�{�
aA�|����Ͱ�5�Œ��[~�ü�qa��\���L��D��_S�zħ͌wi(B|�Io�4����Ox30G�u��+�����ȇf-����Һ՗��f�	>�
(�]�[���`q�SG�]�NK���d��:ƆP����gC��U��(�o!��R����F�����@A ȫgC�TSX��G46�Z ��fA?�?U�%z��L8-�;����e>#�mz�Mf�(&�7P���W�{D��;|54~���;�pGpϬ�\��>Kk`��{l��Z�k��0�n��\�zj�ڋ��^�^���r���l��x&�m ���`�#C�$�N뒇N.{w��]7����OԻ�j�.��Єx�0Щ����v U��s�LIHY}3l�l[̠o0+t�/�_򽄈��:W��6
Ƕg`���H�e�*!
�;6���]�j����<�����t�6�k➩��6�i�
�م`� 9��(/�B(��ꨝ�`WGS:r�/O��ﵢC�c®jo7BvN�|!z�Vwϟx��R����́�(feD�� &oP���0�@���5V����%��6�lI�HpFw�X)ݕH�J�Z��Ѿ�H�_7�a"��|�ihM/�)Q��EƷgT؞�I�LJ���S�浻���z�sl�x?Q��;�;���f&v�4�-@��,�3BN�GM�[?Cڤ3�O7�HK�
\[�����z{p�8)*�ޏ%l���xSùW��"˔fE�ˡ�v`�vs�@����0F�>�,gN�B/�J&��leTi�ci�V>������^�Q�8f9"eSh1�Ԁ6�������'CI����#!ƽ��)6
��{Z-�l�;�`w<̻�B��w�:�"^g�xsU]4�70|��*K$�?�g�Z�;�uF��Έ�sb"���s(�х���ҽ�������YVo������!��*Iف~��m��[����Ng��P˨~�&?�G_VW|P�(���.��l��H
"�I�0e=?��uQ��o�G�`y@}�cwFz��n�r����������S
܅�y{1l���VߤP��B(^��B� �P�?�Ğ��iw����!IӋ�7c�Q<61E���U����9�#���,q����1@M�oV���I�U%����>1�x�	q.tX�}������]�Z-��ĥ�%T����.8Jx����Q�Թ�Cj[�&��#a�M~.[���w�K�Lr6�Cy9��=�.�
Ө�.3�A*��� ���:�n[]�?;ҡ�m�=u9 ��%���8-�6�z���^W�����������+���7C˵�ר4��b�S��kI���]��}|�20fw�.�)�L��T���DsX4�����#
jX�걼��-�L��|K`�_�ҧO�Vڕ8��A�n���}iF^%H���P	������7(�Bŭ��r� ��Y��3GfA���LE��jߓ���J[��WF�X�,��7C���%@�'7���}뻻��b7F�X/qW�,�V+�0�\`7��(X�o�&����ێFQ)�8�����p�/��� M�F"���{����MFѢ�x��4�	˵cz.�<P���5y��$+��jם� ���� ?����7f�l��s��Eu!M�i���Sޏ���l�l%�;����w��#*�ٛS��C�/c�x�u���Y�9h�G_�^}�"`��F��a%~<�J��� �����m��\G!��o#��1�dJIK�< �}�\�I�����
��/�&�=|m&�J��%ټg��Ha��
�nק��O�/��4�KT`W��|c���b�Hg�c����0�ne�1��r�n=�6��L��hW���b�8z�#���ˋ5g�n�UǸ�+a-;��t෵��f��4a��'Q�����25 �ɿ���Q+M�����Á���z[L S�<t� �㚥u`�e���[mc�U�M�h���{����ū'��C��s�z��=S�Q�d�)*mgKS9�.�}���CM���c��^ =��/:T|*�I�~�X�dy�����z��.>d��_�l�&����9���4�Ζ��L�Q�޻��m�{ϭW$@�]"�K���{���� �YV���us� �(�7��qnD��q N���J�J���]i����Y#
�$�������"����~������q�թ���֪Y���3�2-�d���/�#(�n��5�������889�3!0v�Z�9�O��Yt�����8
�P�nu��]�'���B��=�ߗ�������'C�E���x�Q:7�c$:W�pq�cI?���nc����S�q��|�)=�w<���)��2�Bp͛=W0,�`����a)�|:� �uҚ�ێq���U��]�:�ܙ:���]�4�@�ż�%1�0�G���4���{</ϼ��1'3'�JgF�NV�]ޏuV�a��b>�);vG�������*��� �o�&�vf�
���F��>�>�ӻ����y��^Ю�\�7V3����d�0d��Q�pyդ���2O���!SWݢ��G�/O�X�g��1,��TΒ��b�3��x��X���4 1��髝9zC��,�h������6��('���I�@@
6".�Tk��:�Q��cB= �\v�d�/͕qI��@	Ao�����J�;��a��",td�d��N^i�a�_��^����T_���H(��F��{Z(O�"=y�@u�m��k!��:�
[����ߢ����0��"p���h��`ʉ�e��BVƈ��='wOn�ڶ�5���?
�6��x�W*�>j1t��-��-բ�����,k��w�-�\T��f�v����M`M�/�u�M�����> \�N*����l�[~CW�a���s��}��F.��M���'�V����{�S���1�zG��m<�D�Sl�
��]�<?�4*��d"���8m_'MT��=��������g�1t�M�a�����d�*6mq,Ʈ��x���zm�f�7j��;����}�Y3�����
�;�i8����t�h�F��o	T1`<C�UK]2� ��/!�	)�*����Y'��8238�<���=��/��p&<���ĺ�<P��ܮm�Оg��8n@Q�O|
{B�o��&Յ��GF�T0�El�X��*��j�#��˰o��Q��b������ʁ�x/���i���;uS=��EY����2�[�ҡTn�������l8�	��^VAw�?JI�n'6�S�/N!,4�;�U�����昀2n�ެ�{����೸�,�6&Sw�w�<�:R`0,Y��|��̴�g�'o�`y (�Tޟ)����Vn����Q���Y��X�Qo;�烔��r�&?Zƿ�"m[1���&�˲�n�GX5)D��)Po�����2A2���K�.B�ױ�0�rl�M��&�:��1�H�+kS�:�f��"���h��x���Y�-P���g� ��X�P��
�s��堻
_w�0��ik5�I�3�z���B��ꯅ�#��Q�\+be�*y��ևG �T�:���o�^y!�b��|*�f�J[���L��J�:䑈���:�0Ka�@�&K"�>�qt�a�m���Gŗѳ�q��c4wLAW��Z<���� ���5�)����4��u2=( {��cO4s'�c�qtKx揄����3�c�щ�m�+�7�7�̫���+�}S>�� ���.�r˥�ă��!U�ܿh��,c���
���P��:2λ�46N΁3�-v(�@�k"�xq�
O�;��X�8��MSBi����c˒���q:V�S�!T���X�б2f�a��.�<��h��������췔lh+V�������m�ϵ�*�l�4T���/� �(w��A����iM��{�o��' '�iJ���TN���R�skUW���2q�Ml�}�x�+jT��T����#���aF%���c�H,f��-C�m���|
�].�ꤓ*��ąՖ���z������L_��(��~ެա��A���qg9.UDz������o.I|xj��C��qZH�*��!�]T������8����q�KO1�Bg�3G�-'@��E���^g� �v�[�[�q�Mg�ɼ�'D]������6"MN.�п /����߹!\��i�F���Yl����F�]���gu~.�pq�P�� �����,2����|�����*yڏP�����V6��C3dp��X�0��%�1�FC(����L����z����p�^p�+a�d�o?���t�̭RJ�	A�������Q�`���H�t�N���uz/Gד�a�d�9S+�3C���nf����6�D���F�͐�9_
k��o�b���n�������_�<:���e@��
 j�zHn�?�/��n��Y��=�v�&�DFpIV}��E�ro%�ǣ���zipr6���pW�XH5���_/�!&��d�f��O[�����ʖm�����	�e�x�1�=%�ݞ��wd�k�y����W�E��Db
��L� q���p�*Ѝ(oe��v-�����Of�^������|���Mb!Z:ڈyQ!
����x�ːa�(K8��v�g���݅��w������!��ƒRӸ�%d�C�8�,�_�j^E�����"�L��5��R���=�k/�Q������L��J	��� �ᨂV�/�Z�kG&􎒤D�9�`_�����p���=:�� X��;p��N�4�+���O�r|��a���Z���������0�s���S�]�>��P	��M>�&ʭ�]��ŉ|)u�'������Q��a��p��L�қ`�xcF;eW�a�Ի��0h�v55�7�9�}U��x�:��a�\���0zj74ތ7X�ud8h�L���~m/��~@��w�k['��2�!���d��.W1�$�\�)�If]�ֹCK�d���ò�|�Uj�@	Kd���懄��U��� 
L@M�9ᙤN�B�{H�t�ؒ$�����|���BIʧb��κA0(fR�R,�k� �Y�:C!3=����
�D�ߢ��k������v!k���l�^�d��a�$�M]2� D�tv�ƺ�Ά΄Q���غ��2�K?Ɵ< �s��Lp��r*��/\Y��
E@o��gd{�ņ�`<���	�3��I��AV����G�A��"�P�j��i�f����Kh��K��]�t��>޵�Met�u�{%�L��f��\�^y«�]ʌfC4x>�oI!9iTT3�������*5�_&���W��5����r#�8�T�!������� l.���M:]Q�C�ݱazB�i���ͅ[�� ���<4�D|���'8�y�k��Q� zHm�D�}�)g.4	mTa@S��`ŠS���%���D�ݏ�>7�FT�X٬���}ug�"`��]ZŇ{�.�L{�;�cA��C��{Ų؈�3H�G|����4?�M煍��2��lr
1r��[Kf�z�@��ɒHLd�j�k.C�2�+� ��#�`�\�+�ֵ�!��Hf��s4>��c�;�T[����O�~k��x�f�r�G�� �z����MG���oW�(��l> _p�N��f�	p�8�_1y�la:���H�Z�D�|�D�i0I&��#���#�Krv�ۈ�Eg��C�C�g��Nk�ê����Ip��kX��%ڦ�NbT&[�с��k��d(�t�'���"1�2AH]�� ���pTba�N��)'_����ktǪ�o��]c��NS�;�S�gzۧ@��(k��χ=��m_O/}�aJ����"�d��n�3��MU��!�}(����nZB(<��T��Ɇ���,�
 ��r~����h��+�-R�5�ZWz�E���W��:^ߣ�T�ܠLk���ՐN�AG��Mj��)?r��2(��'��,��2�1{p/��y;j���!�Jp���0p`�u]t�3�������K��z����B��H�&K��i��<.M9܄i��Ħ\��=�lE��2'��]�qـ6�+�F�����ƽ�v��"�P-i�W${�I��>吜>����]#�Do|��c8|�������i�|)z����dx���8���vV꤁�:h�/����-*E6�x@��wU��ǈ�>��jeX1���4�p�'�UsTOY]�Q*=]Юf[�0/�~�.�:���x�'�������Ԗ���4��K��@���Ҝh�(<>����Ј3�/��7 D
�_�JB%pN��>�g�|K���r-�e����G����טʴy뻉���P?PQF6��NNdvL����
��	�Y�'���Y���=�A�}+!�-,��-���J/>^���CS�����O-m�Bx�o�4c����u��!G����tz���z���=D�a�������m����eı�1ADH��\;m��Khm;�p���QV������J&MQ |yS�Y�`�|��ډ��h�0Z�wS�p��|�#�\�d���7��|�(Vv#zb�������'W�ް=b�\�ǐp]w c��H�-���@x"^��\�d��>��k�~ �_88�=�p��\�w��7K�@
DG$�������a���-O4ƆcE�s:�Ի�3�N��4�I�9s����%>%�~�a�:>-��;�j�2�'�4���fSBɬ'�Eb8 �pϹAJ/����8�v��tt�k�L4K��0{e�ZӰ0*41�d&� ��N�Sg�2�D�KDǩpZǤ��V�#鰼J]�����b5�7�D�QO���C�����8r�J�d���f��h ތ��X��G;���7��n�e\!�����gu�bEϫ?��'Pe/�[TC[L�����}�e�����Z#�׋[���4*�PӬ!� ��Fߒ��"�w��hkV�)_M����yc�{��8z������[����0"�gC�j���$Pr����kenۄV��62e��6����p��U<�F���6�^Z8���g��d0��_="&KN"�٫өn����W��Z�$��H���r~|N�?׹u���<������(���<���>�̢����$�Y��3�z]/��A8w�z���꾋�Bn^"�'~��4/E��rx��T�Λ�+�����7���Sќ�.޳�CS^E.�e�:kR�=N�5[$�
,�%>b�X�'*�ia鱢=_8���N�����Ê-E���������*oT���l��-��Z�F:=y&�Dt9�$�B����Z�l����Z샨�O�j��坈>7!���+O,x���i��]����=3�o�y��1���7����I^��y�	�k���=%[R�Q���H��!�x|�$[�W0��)�����\�ZOmL3W�.�Kn���I�	�,,U�����/GY7��f��
Յ������?��<X�\�]��#|7'�w��T���J&TҲ�*�?C?���	HhUB��G"��@�c�#1H�"�d*��!�e��ㇺpg��-o��`��U[��fl)��&J��0^���T��o&�s/X��s��gIt�C�֘�q��u��q2j*:u��J�ĭ�3�VH�`�~���U<�l���_yi	d��o��z�C���*����U (�ڊ�jY+���z_���6��n��^�ҡ�.0 c*9v������RE!a̫)�ZC�7v��F~[�H$�BC�Jۓ���el���U�W�$�B���XSr_���J_��m �Z��m��e�L��U0�T�;�}�u��]�� Q�$���-F�*LJ�*��$�XL��J(^����k��h*ɰ$��N�؈<f�bǫ�PV�7�f�������#ڝLp7`X"���\��esș>�Mh8�P�̂5���)�U�,)uO�R}C�#}�:�y�R�*	'�wZ��$,v�C���
_��{�N`f��}�滄���Ф���C�Z�
�W[͛:߯�JT��]����ݴ��+�yf02N*���	ݾ��FWiy蟑��=c����͸:Pt�5��" ���x�)�M_��9�'�����Bi@/� dqgX��6�w*��=�o���~��h �|MKO�`9��qL�'������Ru�..h������;�b̘_�^ՃXJ��b�t��(_b�8&��S����Ol��XŪ�}�)��cA\?�����ʍ���W�^�u�����ɿ�D� �)L(��4b�S٥^fJ��"B�ǆ������g����<4��R����o�OH��]csTu;�[o�1�y�8����LI��6���!p�\�W��9X	X�����-Zs���R��(%��C&�~Kam:���kv��wq�4�z��W��= =������G��䀹�J?�ms�u^�Ϥ�3�?���o��%�b]��,��#*�������886ݠZ9����0@)W����z�=@���1�J��W�ו�`:^��fJ&B1c�N#9GC⋝���@���Smqwc<.c� #N+�5�_6����H}��t"o6�}/�%�Po���_�P�e��)L�2�&t�������u���:�d�?��k[��Vz7�Qr}�JSE5A�3X�.��[��8��Z{v��FP#�ܗ���۝�&�,�Nvj����Y3� ����Z8�1	��B�"�� 0l��d�	�@��]q�s����3bWd�����k~�q�������T%`�`��p��D[�5G��F8�@ֳ��t�EΟ7��:6��Qz�������[�u�E~��Y�S~����$��7�O=q�B6d�+��	.��"��-*�!;�cr�Dg�;#"yL�(���x-S	���fn��ϩ�9����B��`��� j�5�Q�&-\j�{`��%3�~4�P�pI���H=h%
���B�*����	/�u�<-Ć݂�o��<�1ó��#Yʵ���VE>R���#�����,D׷K�ڏ2�̟"wqD*�9Zt]�5�7.O�=�v(�b:v��TfS�/�4`�p-�!v�Zf�5ܗ)p��xNi��M��������;��v
�Ȏ�b*�&�#A(r�"y*�_9���i��U�b��Y�M�\���x��j:�ɏ�ʵ�ǙX
���\匢��-��a��x�-��(�h&v����J���k��p�'���g�����A`I\�<�z�x��u�WHGhOZ���80?��1K!�4K��p�|6��bqf�BK%��%��p�^��~O>�S+��7�c����mosl���\1�ĎU�[z+���oE��݋�h ��Ԥ��s�l"F���p0%1~t��]��ؗ*�9��p��-�"Mp*�a��4�.q���oXT��ch��,m�ܚc�v����f�%o�ϱ'��gM�Ȏh���TYo�VC+/�Mj3:�qNsfE��?
6G��,�X��z����^�5:��QMs~#I�5�����ؖzF̋ok3(!�VzMAW�iDV��Zo��4�N�D���Z�t�W���%b���E���8�X��HA�y3�+�;�ޜ9@�gX�'5D)-�AԎ��vI1p��tұ����*�#H��]�t��H��w(N��)1�.k!"�Bx�F�H�pje0��ޖu��-��;@L_���Gan7(9b�����y�.Z 5pQ˞e(9q�^�d�-�B7��C�y��1r{���7!��Tzh��	�3���;�Z��z���i��CXnk�)6?0�?nx�����6Y���g�08��hi����ˀ���;�,���F�t��)I�����(�U6��o���&���-��?��9G{L����6� *��_�=�8�{u{	�st03a�Ts�݄�����͌�����c�7�۴���oq|*��5hy��e��N+�Dּ��$���;WFG��d��TvE6�c;.3R��ڧ��l�E2�|;�.B1�f�����9�8m�����5 �$�Y�8����:�9ǃ�.�ZԷ]��y삮��nh̀4#�\�H}��W�蟱k��1F�dQ�C0��,*��R	N̫��!۪/�Tp��r4��A=|���k����!�Y��ZuŇ������+B�p?�ٙ-��)�!5*���C�	V ��������	֚M"iLܞ�����i����L�nVuO��m�?(��b�r�KY���_GS�3UՒ��~S�z�ճ^Ng���a����q�qH���S�a�GƯ��N8��|�(�9-1�KB�Ł����4>T�_�m�8$e\��.c�Ň0P��?��PǑ� �}�Rw���c��t �R�5��c�x<G��ύ�s��:��y׳�s��	VZ��~V�\��3S�[$���Y;_��l��a_͜���}��N'�h�Q��>�#��]�g���b7�m���jJ�s���I�_�~��A��F�q$Ő�fR}�b�If�1<"x��T~d�9��ȵU�<��d���	�y?kS��z�4в���ʜ����=r�s�c�j��^�ӛ�4�@���|3��K��}NV%�k�u-�5�&Rс;`��:��E�>�@~��n�к���R�N�^��4�N<�~�W~�$ ����hH`����a���b$_*T�G��:�0��Î��������K���\�|.�>v@6��Z����3��qj�P0@쨦�Don�6��U�}�	9&��D��?�틧M��qG��<�̬�g�I��ٿ�5X��R(a"�yG��\$�>^��@Ê��Mb�9M��ϱ�>�ꄹ�О����܈�ȭ��C ���S�"�����՚�����h �����!��3�e�z�`CP��g�D2Gb&.���-��7�53τN�fX"|o�F-��=��=��mQD;�){��w<H	wj�j��_fT���T���SQ#T<-.D�d�k��]���)l�Vw�Q1p��֩���W��aox� �A���C�k������%^��.CQ����L:^z-�nI{Jw�hyi�5Ak�`��|k��7�m���ϔ�)�s2k7�)��Qz��8��N@B-<p� ��j�zv$e��-�P5�ξ.�.�N~c+��I1Wh[�B��)�מL�r�g�ʗ�`(s�EyF�|�	���Z56�V& 8�=M�c�:Q-�{L�1gU`)6��mNp:�Wi��ͣBp�\tm8�S�dI�L0�֪w!W��ܞ־۽�Z2�����W�0��� 
=�Z�j#V2`���M������hIn�p���r�:��Rř���5M!M�_����*��p�j�ؠ����R�puεRv������=,ڼ^�R������"�/���&��aqh�} ����$0�H1�ȪV���<�*�-j�;.$���3�1-2�?����NjN (��y;�E���U��?U�(C�|��8���dM+%���FP�j@�W��xa�\	�\�f��`0j	�Ӣ,@����S��B��?2Y��l��g�����Lt��#��߶����\j�����v�\2b���T�»�����g������
M⊙8C5qJ�bk�s��F��";E��.���x�{Cј��)[����I����׫��es��%����s�V�~���W^m"�}�_7O�;0����s���^�v�s��n\��9���e���X��0.�$W^�x�uoE������ܨ�2��*Tt����=q���-M�U�}e��i�ɛ<}���|�ؒ�l�I��ҤG� ��\z�3��Oۢ{����/����h�P�h}�z����o����&�B�Di/1͑DND�˺Ѕ�_@�ܰ�z�k��jt���2�(�����i#�=G؜��,H�G9�ꇿ�Y؁��������?s��d�WMt]�#�S�)(�)�;�>3��u���9֊#� $`�UWz�t����;�Ң�B�� �2��p�
K�9��A���s��>��.%�ռ�G6�D ɚ����tz�Z���c��~o��51g�� 99UeaxG=��\�"X�S��J���=�D���d��*�hgp��Ӱ���l�]ܕj���Lt<iW�ɧ�ũ�M�_#�L�l�V�#��i1��]u��3��S��n��{=Ssə���Ϯݯu�j[e�W��3aY��`�6�w��H�B�5�D��\vI�Ud淔�� ە���V��h�>Aj��Z�(�㎢.��e���?]�Pr���O(������� �Ic\B��-vJij�4�J���	�J}:�?ɊRq��n�_�'g5ږ���2��H}��:P��'�!u�Ӻ@H��>���y� ����L���҉!��A�Nڭ���6��au����E�%��̮��6��D�Ϟ�|��*��G�ʏ���s.�HWɸ?W~�v�];��i�D����煫���<����/�??)��= 7��r�E�#��h�+��G�N�����5�=������W�ήN�}[�9H9/A���V�Cӂ<Ƨ-Ѝ�h]�T977p���{�*.��r77��v<3S{��N�J�2ب)�
�ѡ��H/+&��)�I�3����I��i;`��}r� �V|f��G1��|�@[42�}�S��e辛�q���N%��~m�>s�k4���	P	�4HV��^ȗoZ��v��ڿ�m-�&/A���j^F�O��8M�F"�2�@�	�6\�գM�a���=+�2%�)�h��}�"���}w��Z�J�0�����g3W�I�ÑԺS;fm�ר�y4
�O�W~	��� A�Jѕ[CF��ڡ�|��5H��}��]��y�)˟k`�� ��dߙy�s�$,�՗�%0E�*�B{����_vǍ�Je���5�p�+�ʝ��{Ku��7�	@)���_p�3�8�`�{��Q,n~�xVObXG<�Q7��)�H��i�Z��m>{jp�`�>�7��L��!����X}�	��4+an_�ZNw����8���[d����A�&ˣ���JY�� ����'7Y�xq6Ɲ�V4r	g�E�]۹:�$���TY��0z\\�{���2��䬨@݌mإ���(��,�p5-�Q?ڷ�v���=vט��	ź�=~A��.>,�D[?�N���S-�B���� ���>�*���­��p��E��/������ho:`�ߙ���fy�H]Wݻ�y=��2�r�e���
�=({]�5�'B�y�z�� IV#^�>��\�#йr�m�����Q~�nw"�����A�F+L�m�HQJOE����ӣ9l�Gz+��f\�0-U�[�S#k�h鴦�r��"��C��#�P�|:�C$}/ߥ���)w��!���bs.%;ßf��mf�*OP�H^���k흪�NN|#� r`CY�CJ]�İ%�c�r5=ۙj�[��x
ǳgL�C�5���z�$,n�#���M�ժ�[���R9E�����[�k�]=Z8�.�Gq忰�L!L���
����I��f�\Xߪ��Z�wG'2��b����ӿ��9�WR�|��`Ϡ3������6�����b������2Q��ۤ�ן�ƤC�<Q.P?�����P�֎LE���^�]��d��(��dc��5�hV�K�w{�xЈ���p:1] �A�W�3����FxM�x .��g����STD�sV��l�h$�'��n�m�Gz�j��1�G��qFe����ù�=���)p�$��v�����esR*ҵ�rj �F{݁��,��G<aEՓ�m�:���׆$F�ZR�f>�u�S��`Ҫ�<��>�����Q�����i~g$1�p�%��^%��df崒������o�Ǒ�s��M\5�J�<Hpm�`#��%U�\h���lE��#�yX90�W<<�7ȥ�ZQeΉ
*U�WŐ�������yo؟;q����=VؚC�2����&�!�Ơ�0�����"�"�,�xuObU��Н�ݲ��)lh��$|���h��f�"�N/2+fπ���s�f�uUJ�#q3�?���;�����ـQ�k��3����K�U�p��Kf�@��`nz:��;�Ez(���܈���ȡ�|�a]O&2�ċ��]�B�)g$��`t�eRx�Y��G�
JJ2|�	�'���^�D��x�=%i�;~����]�B9|�5 +'���\����ڵ�5@`R�s \�&]A�4���/� ��,����#9<�(�8j���Q��}�)�����1找�5���py�bwv�ñp],�:�P�I�_g�i� c�,cl�M
��'��b��k&�Y.r�������%l3�rP\�	(�#U@���5����c��҈�)�3�F[f+R\u��%��.)�� ��Cyx9���m��3L�|~��V|�O4 �l\<$� ��z�2��?-��6��H�e�z��P�*-�	�L�rj�65���)m���u쎂:ۉ�?�����v(]���$2��lʴ�Ȝ,��X;��~=�Q�ehA�^w6���� �7���dO�W�hVA������ zJ�g�\�� ���1�=w��6��yF��ɶ��f���G1��BRQ��R�����R��5L���J��tg�������Т�9=Z��%�a�D�&�3��x��	��A�LD�_7�F~�ػ�IORdw�i)�Ci�o�K�����	���Šb}̨  ܋|�w��}����gעM�5�JD̮��F͚�\�%�	l)�&��s�P�x\	(-O���/xW����9:8�}��!Z!~�h��	1�2�2��q����N�[Җ�*��9�p'�y[U�,^^β�v���͕�� jm��O�L_7�,��"�9�8�R\��m�K�~�H2�3/��N�F;�6Vҿ��X��9)�}׳}�&�.�����Ϗ�w5��&
�^û9�v�����ח��%� d� ��3�9�'���dF��S�=dX�B都�ĺ�感���^�STn'����|�_��ē�-�en�[<��]��!OşW0lv��u]��(��t�ׄR�DG�̦9Lw�X�S��V�M悗U��#��'��9��N!��Y����L?�mR��n?������Lq��e+	י`v��1w:g�*�k(�1�ᇩ�sλ@�1��}C��6j��`��
�5*���fl��I��,�S�E����{yK`��b��e:�9��a�lAY�HU��;7O8z.3�tc"?AR���C��HC�]�kf�
$���N^k��T���3�nʣ&#����G��Յ�xu�@�*1�f���9%A�L������7M�'FF�)�ZpR�}��<;dvx��_����_κ�ߦz�|7t��5[�?�Vݻ2q�f0ӱcL9K�}%��&�f&x9~�];��uo�������j��p1^�G�p�7������<򎧨t:��G�j<1����[|#3E�ef���;�SXo2D̵�wG<D��������	��[�PY�T�U�7�tX�]�a	�ɂST�	N�����玜�oJ����^�OgBWg�p��i ��S6:]u3��O��/�s�p�(�s����%��}�� v:@���D����YgG��m��;�F���	t�n�f�o?bf�t�*-a������bkQ�$�p�o(�"å�4�"��؝`�����f�B�G��6mt�Ї����!�Pxe3���hjqS�fY�N���t]p���;��>���;�1q�~��u U��ۢCPev��ɱ}+��U=�"1��`җ̉)�c��=�[nA{F���t����55\�dق�����I��V��'�~�����V��~��Z�#�SQw�׮��Qw�7���H�%9V��)�5���A#�*�ϰI����[�*�c,,=g��~�&)'od��i���K*A�`?D
��b1�&�n����9���譤n �����`��]#S��Ɣ*�Q���ƐQ�&~9C�n~RWM������,&wHt#s�t�J���B�'>����g�Na�N�9$��mm�{bK?ueȄ�s^(�5U3���e����kV~Z��
��ʂ"�veB���j}:|���l�	�:�N�37	*�^�E��d�$��I�5Ǚ��2��B�X������2�j}<;Ä��B|M�3��[��+�����<lbb|6{-)N_Y/V����h�0b����Г���.n���$��-�6�}��cQ����z�[�9�����e���>��B]	��:En8����;8� ��9��A6���ݧ��HD���w;�ܖ�J�����:k�S����0i^��l����HfB ��|�?a�p?<7$#ɮ ^?���,�O7�<�AC�Z�������Of���v�(�bN����`Ym}�?U:/۪��DO�1���Se��j�������j+ɴh���Ӟ
W��멅���@��]T�ҹ�4n�}���ò���4@N�/#E��j7���:����T��B���ի�Z{}�f뻖��q�����XG�����Hqɝ����@Y�ΓӿS�<���_K<,� 3�	�	p Ιg꼍�	|)���gX9��	ީz4�1А���a莌��*`��đ�?��b��mK��v��xj���S|R���PP��t�������j��� ��>�~�YTV$=V΅v0�!y�,~
��Tn�_����͘�[�c$oBT��`�؀�uĎ�y�c=gU��\W*�=�P�~�:����u��%���'T@xp�V�:�(���i���Ϙ?=&��7FI�:�.�
��j�O����$��E����,���Y�H{;d�~5
�1�hc:�s\6Z<�H�)"�k�����ݓ|JC�!�L������K:xF�YNz=s}��&\U�;~sk��9�ۘB_���p��x��8�|K�=�r_�����94a)�C�s>|&t+i�}Ӈi����bI�H���=�
Q9i��n���h8����l�T^�#Y5�	���ڟ'X���7�h�p8?(��S\F`TZ�!5������h��kٞ�m
��qw���=&i��V�J�5K��u�&�yD�-�V�k�z��{��O�k2uP8՘z��~+ ����6�?<��!���!���!t^����"C�6El��s���J�&z��Dl�n�D�'�[���s@�M׮Lt(fv�7����T2��]�����35�jH�P�UxU�p���O��<@�~���(A,F.�������:DFܹ�P���]��z�(��Bi��ag�����l�����l��|�� ���m(u×�r � ���`{�c�I��B���U�t�G�X�����򱽮��%��g��2�PE��T�v�
a������{��;䮹pu7�ED���H�*;�aO$�!0��ƾ!��_��X��>	������/��W�1-����{���~D#��+��2�]_v4#��y�� ȑ���R�"���h�R���S1�=�B�t�}�Ȝ�I
;��+#iQ]�W)kޖ����Di[SU���� ���Gɪ/2�rp���U�͠,��C�[�����g_�I��`��G�;�]�Ǿ)���g�m���U>YAsX�ȁ� Gx��{����䮂_[������a\�����p>va}�~��|9:Tb�'�������Qze���dDdf�\�t<�aWR/�֚�?�������F�N�9�M��5�?SS���E@ �T�x���mR�Bg��1�RQҳt�	��YX��7�(���GTT����ƣ5�	�k)K��$U_�˰�K^	�:}S�g��e����ļ+�p>����8M�F-q��P"h�������7��9�}��"yY�1��Mz��!v�* ��?�m�T��O��;�"V�aL\'4!`x���O��6L�3?	�+�0�3N��Z���N�4��ןZPI�߁�{��8���Ȩ=���S�����,�j)C=ɮ��w�A�kB~����
�}�B�GY� ³��%?ۻ�q����+M���?�X��ۀjU����{�[X� �@u$F����1��)�T��U��yʰU�Y��s���r�J���)$E��ch�os��՗N�۶�+��@�U¥��aťF���&�7�u�5N���L���?��qV�����UOF
��*�B�z|N�ud�^���:�s�9,EJ��0��{7���O��D4O�>.� sk*�q���>�N��g<o����K�ֿPN�>1��J�<��r����c�@��ߐUm� ��%-T�`{wC/�~`]�|�2G���L�T���@
� Z�~�`�����+�/�Q:!曔I�r?yzR��\�蘹)�_�cfj�W���X��i��W0�Z��������W-�0�PK�yά&4PTB*�~ָ*�"��,C#��k�����Rn�|�ua�Dm�i��Y����8���+��;����(�B�&:�s�hnӖ-ŧ02`T��.{ߐ�����W1��ԅ\ա.6��"�xPFe�"Ԏ+�s9{�,c�Ɏ��i��n>��.��Kp��5Z��vn���$��[�����Rwv%�ݨ�7�"�A�b�Sf2�m�wSJ���4%�S�`��6���,m���5�o�G$�fI��$%�/�Q����`���]�@O󬜧�{��kƐ(

&a~�2��mj�	0]ćq�b!�
z{��WA(��ۙ�����{@&��ˣ�Ν��WI�@���<|f�7�Iǆ�O�"��0~���N��#7*Ȭ��Ro��y"���� ���RX���1bX�U�UQ\Es.J���߰f�d����^Q{�|���r��YC���x��Bj
,`!��E�㾎-ew>�[�^����ML곗�� ��$���\#k�<������1���VҦ�� 8C���/�[&�����s�	��
]�%�x%.�z�����I2�c��0j	�	(���.{��V���5��ܷ^込��.� `��i1ބ��TTy��@��a>�:�*6o��D+8�)��X;	��B.��哊L�]$��k��_X8%	�*Ņ��؇�1F�	�ԟ�^",��l ��i����"[��'�4��U���>-�$:� �'�w9�O\ń�y��E$)���X���Z��ڭ%��������`v�3�!�"ϖOm>"9b#+ט+t H��4@ݺR���^�����Q�_z�1�Yy�^ɹ9�*,�0U�L�y�am�FS��˗{X��Ss)yI����|�����CJY�����{�jj��m&7ە#���Б��l,_|(\�ux���|=��;����-9Oy�vk#�y���H=ڄ��v�sG�W���Ц.h���rGR;,y8įq+�t
]D�5��e�^ <��Z�vM!�S�=(%N�P��~�bl�C:�7�}��eE��Ʀെi�f�S�ƒa��C݊��f��{̣��b���OC��-ު�~�GLR<�F��T���S0��.Ngl�oCsb.��k|��_��BO�f�x��͑�AL��k��̔6�0�w�"��4J�7���`�N�"b	D�}ZD��Gۍ�����x�ƒn�*�Z���>S"�h`��A]tYIUS�~�N��DH�Q����B�*�S-=�=�
����(i~v���N�me��:��G3K!E�6n&�ps���Sp��0U�*8@��|�Qq���w��5�xF�h���PW�$��E�߾Y^����|�K[1�02%;�����~m�-t��$�s����9u���T��GC�g�#�<0�ie�;;�n��m/�c-��If����� }�5
��\�ܵ<$i�v\S�p�\��������c�ӽu��9>L��]��ae����D�2k���+�c��4s�������ܡ��^p�ɳ��~}B��yf�����&.Cm��6:]�>8d|�[��j��:3�����Ʀ�V��d�����?G�%I@YX�����(˰�'�D�����|�`~��I
���:���'�8�V���)c#̫[����	(N�3��A�*�\��?�R���H�MQ�U�Wa7lH��~�ԟ���?pd>[h�W?��v�&���8{@�A�O�?�ЋqtX��Si�\Z��������"1+����}�6����2-��4n��Ն���Ć�N�H�!vҢr�&I�'k�uq�1ݤ|2�:�2��+���5�`����mR�N��z�8�������x%��RУ�������S�:V�����]��|�� �$�:�@
X�k�̀�[����V	�tw��_e��×�gp�ވ�<�E/>����/T���_d�[�OS�V�#*����%��:zg��] �Yχ[�]�:��u*��5 �9�N�B��m\ܛ�ɚ�⨡xz;��1_�h:�{5��A���!���Ml'�[;F_jw6���zTA�B���������}E"�S��6j|W��X�i�o�B�|�k&�@QcX'2d^h\�u�q��/4^~~�ʃ��.�������7��*7k��~ z���X��)L�	���=���BA�����v�?��ʯv�'x�x:@P\�cN�׾��B`�9b��G.�*�R=y�΃�I�O%E��D�a%}�2�T���w������:aqK�kBaSG���m���?���+L��B�M?C,:���+��s�ɩ!VxQ ����a�c&�4L�lȟ���Vy�߱\S��" �����@YaJ�*�/x��e�*5�	�_瀧�#c�/6(uce�7S߳�_4ˍ�=�˯��V�H�QJ� �
l�K�gt��~ɴ4Z��,5�����G�L����0]_n�j���(5�00Y�z?#����g��f����=��=[��n��$+|axԯ��i��s�!ɚ�f���5�����UF-�SB)�[Iw$D�a2�kW��s��� �+���E�ϻ�}��V�u���nQ�}Ļ��O2���B��xr|^�V1�`���~b:;�����iI*��C�*��fsPKD��@cs+[K��T�k(Da�ݑ';b�CgO���,Br=��)p@��?גȍ�nr���/�I�|� ��U�+
2�>Nf�ιrC�5��-E�ÖAX��\{ٮ[���� V���I%�'�\1�hEDh��0c~�~�dȒG�3&���U�J��tє��N�[c��˾_�h�}��T*T���Ǩe5[�ԡ�-^�Y���'0���/�?��R���v�и�a��e�-�>v�q%	"���>\_I�_�twcG�h���v	�~����Yo�a�90�%�tw`d���?���ې���(����c��!In�]7��AR�!aǟk�E�q6��R�VM-vVZǳc�=��h/`�siq��p�����$�4N��Tft��3C慌��Bb׀����ũ���(mL��UHhs�������ey���?�O��	��\!]�����Vo@��#.��w�E��)��TK��rP���uu|�r�̆�G�t�-S�x����k"-��*b�\�K'��bUL̏ՓyC��[U�G���(o��~��'>3G�-��̸1�=D������ۚ J��(C
,�UDs�IE����x����;*΀bF����	 W������� pV��TP�(�僬�=0�K��]��Hf�[�f"��T/��J`r�A��ړ�����=A�q�`�p��eY���֜��_ѡ:l�/,9��!�ٜw���j|'X�PT��g����y�8wD�	x�
��쀣k�;ff��&�?�t,�r.MG���
\k��2��Xi�y�2�/�q��+����n��!�B�F	���/�����{���Nq;[�oA� ����������A֔�3��K���/�X�x���cvЦ�~�
9E)�M���:��z�t���-�Fe��o�\��ߩ��_��������>�����a[�J0�Lq�:�GxX���p�BS Obޭ��an>d�$1d��I*��USYr��rs�#ſ�%�̍w�5�y[�̀e�#83y�4ȃ��Q��cq!���Δ�T��a�3���
��8,^�3��39sx�Lxy�^[���Y�T�����g')%�%��
�K7'�߅��z�u������@X�L��y�_H����H��ʟ�h�C��_6|w'��'Q��u�͓��w����@q���|GN�
���x���ϣ1N�V�L�4~������Np����i{����^Y\�V�Xe�=���O��G�9t~B��!�]�>�t�G4�UK;�S��0�X��K�ҳ���H9ڪhw2k<,�.���Ň�-=�u�}�����k��[i[������tKs�}t�v���~r����N�����6�q��K)�����J��Q0��^c��mßk��E^��{T���R��
���]c�T�<�0�S���S��Tt��k_��=@$���LGCi�T(�	�4�]���9W���Ґ���p۷�~��WMf���
�@�����-_.��oc�SOǑ[҆�=�Xh1`��h��J��=�p�Fg,4(����!�?��j��0���6�*�+$�?����0]�Y<����?����b`�g$�%�#�G��1���ԥ5��@u"+�ك�,iIu�����/����d��t_�~;���e7�)n$�	v�tj��Z:�l��ː�W��b�"���½�lZ�`����L�)���Z4њ8�s�i��Ёq��br���u%P+��3�j��u��Գ^u��f�n'�.������A+O��|²g���z�s���������S�̻Gh�u*p�։Hż_��c2 5N�������������_$:�Q��j��6�a<��2�����rtd��"E/�Pǎ��f�[48l�|������>�2Y���Pp%�T����^��Q+�1����Ͷ3��٩�Z�Iy�/ k�4\�r֠�ƙG�YgD�̔�aS������T�Wj����G6�%H���4���g����3ja[���J}��v��K���*i�vxy5�aًV-�'CG�[��9!-�Z��l�@�v�.��Q��2	��W�Y^.��Q7��:�R�bw�3D.�K����}0�0����+�����,��֜������[f�|+��(��7�.9nt1�<EB�W�&����V�x�2Į���gIz���*ڰ�[������3c�$&'��J�N(2M�xW��#�h��X�-
�Ս2_�C)��;�:�!��m�*A�V@�ᑈ���CvD�<�gM��a�	�*�yf�l)��J1`#�GWq����i�R�q�R%�(B��"	F��
1�

(w`�d������:-���8蝠
!�=�����"��u+H�CIg���*b�/{ą%����卅T�F��e|ʪ�$n�#��e'0�C��z����G�i(3��Y
���Vݽ��_�yE���1:gz/���C��+q��ث�W/ٟ1�d��y��Ǎ$��PF*^��M��B�lo�d��>��<=T̰�a�����i�����%(2f�U��e�ӖMދ��x�Mk����F^�c4p�!�O�V0/�Ԓ�!�UK�)�nw�ǋB��g�G���onF0�x��,97zٵ4�/sO�z�a�j�t�2��(2�?�N���YlmG�n��G�JQ�X<n7���m���X��n�ӡ�;�b�l��}��fk}9�% ���~�=c3<��ܷuj@۬@cO�`�^�v7�����H2��	J���e��>c�gS��JB�~�5Q}Y��ɪ�H]�%��"�s�a�&.�-�a��R!�h?��4h:[ �s�Q�D��R����n��rڔ�=ژ2A��{΃��;"�?~�>C���<�T�z|�ȇ��n)�Os��:�8���3A�K���N߭�k� L0���'��娫,�'�xDj�9m��,����h9c[G��>�vVϗ����+׉��:��e`�5Y��4['~;�?CF�q�Q/� ��X6�R�>*Mq�`�O���3��}Ք[~�]8����E������*GN2�[|W��Pn�"�:��R�Y�`��0 ۯ��֕�I��aA��m�Q:�����Tj��7u�BP�U�S�E�.����#�F,l���M앣Gop�}G�J�)Zө�o��4;�V����1�	��I_$ǚ�5�����&�V�k(aY,�@�jq�BI�H��Cۯ��1il��]�NE��,J-�S:ڌ Op�ρ��g�T���%X�
q�R�� <C��xt�'b$� $f�dڱ���?�Ѯ����;XYY��'6�El�J@�1c��LtM��$�:sǬ?]��cIˢ��a�3�+Y[�Z��7�!��I�n�e���X�֗u�?�L/}���(r�}m�u_����z� ��������\�8M��ݢ�kc�˚ b�<�&xZǧ:�J�ߚM-��Y��h����+�iķ�s$&�mt�^nR6���J0	���~yؿ��8L��f���� �L�#�"�o*�wዜ��$�T�1Ȗ���(����لD�9�9}�~��	t%����3x�E+C���d�����# �H?�Vr�TণH�/+.f'C�;�#N�
���佾v.Q&AҚߌ�TYSoS!��2�� ���a�-V�:Pe���M�����)K��a]JN�xQk���:El��)���y�а3�AL�@�GȀւݖ��C�+�j����s?J����R��y|�d�]��;���ם�V2B�#[���o�q�L}�V�N#)��=��U4�u��$.�����i����j�Ti5�dh���T�<~.��Wg�<��8��s���eg)�4ٿG��F��f�8�D�B�F��T)�ڊ �!f՚p��s>u<�W���As����{w�o]�$[��>�./�H�
�Mc�ի�K���o��|9m[�p�7�Q�k�P.%Gu`�����U�%�^��!��K�~��p�E}�W��.���K�%� �]���=r�}��zj�}L+ҵ����������@G�q�Q�7�eNJW���$��r�����l���).GV��e@���!>��{�%c��x`�X�P�V[��UR��m:p�C" ��`E-r�QnI#)G�eg��.��ͯ[�FI��Pڦ���)L��٨�q����ȡ���*�������3�*{C�ZRng$ʣ��h� ���n"�B�3���3_"���ֹ��g=_Rvs��d�!���v�]E��'|n�g
�]a��?���<R[���q˹��m���.yK8��H���ZY�>F�o�����.�^�g�=B^���N=��λp��k�_�U�y�0��X��^�>����u��BE�0�_.�p`�\YʀF�:P�Nĵ�509�s�r��]gX����%<H����2U����G��｜�	9�Zf�Q
J[rI�_�n�莳��Լz'�;�!����B,�}�O5�Xٿ$��o��Z���=B=+�?��2�E��0Z^��20+)s���M��3Q��D�,�fT�.� �2Xr�-�������!��3B�Z�oT�-룤�C'g�"Ni.U��3�4U<�3�,5�I�f��%�rA���q#�6~4��&��`,����m�\Ԫ�{�S�{�~&�{h~D�E� +	��Il������2������6K�tQ�G��+�:�c�{� �-'��?N��W����eT�|�>�3���I�����j�
_{&��pQ)b�s�F�mQ*<2��u�.��¯�Q��y�.&A.J�_d0�L��=�<��b�~ w
/ɠן�����-s��ӸD����g$蛲����̺�y	;�fq�+I��!e��ˬC���ި����t&1�R�����!��d�����!�&�$.����
���Cgѻq.�U��is}���X8������L?>2M$ N��-=�Z��ȳ�J���g�RHL�'<�m&���D�$���
���c���D<�V,�Z�zb���c#<I�L=ӉHcQxq�k@�h�T�[�ی����ϖo�ʫ7娃Ie��|����lzC)��W�Jq�/��zn���W�zE�ӷ�d���u�Q�/ު�;���0E�\g����N.%cT�C�� [��$��'_�޿(�_) 1�p��>��N���md�T�D�K�m��靓�BG�ЙBd��:�?%��0s���(���q��i88�D,� ��w�]�FI��VR�l�^�p/�߮�4�i�ߓa�JOyw5���h��M\X�-��y��c�$ڭ�2�n�B�_'�vw�$�sQ�����b/_Fl���d͋��$r��i ^�v�ID����<��u1z�=������H�:΁I��l]'�ǹzx�l0��E|��W֟,�NC����[QtG\{�p#��ŷPB9���&�Ã��J�ٞ	�
~��T�b$Ҫ6��Rz�����������t�լ�r!����kz%�HT6_P<�Jۧ�V����?*�̠g"S��3�ԃ��3��B�s7�KK�r���
�w�?�fT�ATR`�/s��v	��-�w{!�-��ӝ���yЎ���B"<	�_麯�{�V����[��z����S1���N�5�E�EWzT�I�V,Ce-�m~�SN��S�>\B4X�H�p=N�.w��at�ױ��~ui��/�-9ՋnV�㐑9	s����@��	=%�/6��B�:�4�Q��HMG�L�����ǞLM�����Mbr����|S XM�1����2 ^K��^z�6�H� zC�,��գs�[�&#8�)��^�g9+�������
�Ր��C���^��K��6j�^�g���c�k��b�K�������k�2�Џ�|\f��Z�E��`V�������hP����A�pS��|�LK[�TCf���f?�D\�U�|M����n�Z�!��/7��9D*���/�
�t�^�a��
���͕S���Xn���^1�+o>�R�!F���;��E��3��%���=�.�-������,��=�?;�RI9w�iM��c�� �:d���o�E=�'ɨÍJD$V`tj<�	e�>J�\�<�A�LSe�i_7����<+�_�*���U������ �@77J��B�#f>׻�z��3\�jv����Z�惜��(5�u�ޏ�h���*Y�ֹp�3� �H܈�	�X�4�5܀��C��u%]g5k��6����o�-�N�w`V*�<��BN�^9���d�"1J6��K�$㄂�M򮙩��OX�]���������i�wF�	Ij��6�S��,�%IiG����
�vr���j�F[��_��u�up ��W~ �0�������Ջg5�
i�ۖR����'`f�V��U\Ơ��Ơ�S�~��UQ��',���f�̅c
pMf��Į�|9�1o�9����љ2�9��GQ����w*�p��*�TW�F0�7�����Ng�D"K�C����ƺ^c����V^Ս��..vDs�Ձ��ȏ��zK�6/d3���/��c��{����2A�p�}4.og16�J�j�T*�T�|%��_��fY6O�:@��s��O_���F=k�(�-��ۆ���D�s��J�e�14�}�cpo��\�z�_��ӳڢ2�©��pr�P��f�(�Oӥpɫ�@��݌4 9e�'�7�5�pU��:�ڬÆ1][#�6� ��0�Y`��'c燓��g8��1RT��
�ZvI�>O���=�%�"EiJ6el�
WOS:�X��� tw�q���I�{��l��*�-�5��t([>h���*�l�3�N��w�;!�M���4܇�Ԟ����1��)��B(a��C�g�,Y��0���� Ur��d\���n�6�3�0 }�_Q�G���������R��ey+�6����o�E[�D��&+�|����	v��Q��B=�c�����\�-�	��iz�N�Eɨy2sit�q�U[wp?z��+`~-��p_�x����:[��򗱫����_��w~d�����jUoo<ԷH���Ĭ��/����-���o����"!PTl<&�d*�6�߶��)�B3�{�U# 5I�WL��釆�A�7s|��qͅ}*���H�_E�{��K�f��~G��������=��i�9�`nS�A� xq fc}5�D_��z0{Ⱥ#�B�߾N#�9[-����a�u+Rc�3�/��ff-c�dz�����P�����gH��ш��ܻ�	Ev<@�	%v���!�q;{���Do�w�e.Ǫ�#A�D�a
�Ҙ)�t�=�ݼ;fɣ�eU�&ԭ@��̙�4�A$��t�;QJz�Fa+Q{&yo�-���=)=�+x�%���q��-�m�lr�(./o��S,K�L��f�6kv��x(�r��I������� ��Q��"�Co-t"�"��Q�C٢^�7�jK��ъy�w�(]-�[O���R��il+��G�Ა�8�_@�Gm�����N^X�j�yK�/���:�FI������QT�N��
�}]��VS,|ajqEU�3�xgڃ�s�l�*����l�{�<0E467��wZ�����~/�V��]b|�f��T���+:2�u3�]=/,�)m����o�U�����b�Ϥb�-T�N����Ia!�A��F�5;a��u�F���M`W�d:HB���$�6�NM΅�_�D��Ȼ*�[R>�[�:D������C×2$N�fꔛ��1SB����y��b�B�S'� }�N�4�R���q%�ո���C=Y��~�4��6M�K���um��S$�m�t����/��9*d�n�	���o[v�X�[�|�bu��"�g�Z-hB��\M�sS���z��9љ4���J���qkӸ���5�;B_F"\5�K7'Z��t���!��d����Q����"ǐ*m�P���X+�ӥ4g�Q =x1�N��|,��������9��N������Djy=tg�NO��:���&T1���7��n�J��7�"w{.LX��چ���)BP)��FU y���`�!l^C-ּT���/mTV���)�?�͛q���i��ª�cz��g��GX�o�x�W�������!�q-��q���85'�O�����Oz,��uu�9#kLcd����>�sr��%��Hp0kׄ�zꎭ�]Eog£�8������2>��,\ݸ׸�Bq���� ��	K4�}a�%�)��J"*2�F��ܻ��d1oT��p����	H7!����U	(�'<J@����!�D���:�kTQ[����SsnW��b�O�w%�/��>F�i���>�o�#��\n��f�O�0���c� +�~<���G�r��]��P��
7��Y�')��N�z�p��k�O�q^�
gj�2mG4���͛��vN�z�\y�>b�@�x����b/�c:	e�g�8�ќǂ�ƞHgZr��F9"IPZ��%�1�Z���j��/�.�"$��)��NR�����9�7�_?._�
&H�����|~�e�.^pB;1�D��T�No�K������1)Ra(:G�\���%gP��
�e-.Bm���>N��:C���?��Tew?��� �0��( �a+?(��9����ΒKT�K��,�t&�D�#� g�鉗�9�6�C��0�m���G��:�",.n#a'������ �!)s8�{�lf���6S��KSm#+D��4j{��))ϯ����\F�0&1T��"b�y>�}�7�$;��-�0/�+�汗9�|]�&��ޟ�ts���׽5S�����[�LQ��_?z��^�;o̧���s��g}�0g��D�]�����;�Ro1@|US�o������<j�pD�B��k�z4�{�[���$�������O���F}�JM�/��]9��?3L��eP�<�����CY�d-�����, A=�U�m	>A��e	�3Y�hbJ��m���'�5a,�j�=MƗ%���3Wl��O�x�v���Dd>�F���p�ϫva��ŉ߂hSY����m����� ���� #���J�����K�ӡ�Հ�)�F$E��b�����*B�]�K���?]$��/ ޘa����A9G�~�\��K�.
"�aM�#�J�Aann\�q�NY{���.HC�<���� 1�g=،2�H��C��V�� ��� �?�}�eW"�x�vR�l�7�-RD�և����u�< <���	r��Ni�7���$��þ��1+�"f���f̝��ga@'��e
u����v��q��3��ZtWHy�S���B�Vb+S�tמ��e��ʂ��Y��St�QiY�u��R��U��N��r�ϑ<��4�PsoT��I���!�����H!Tb�ar �eG���W@�\Wj��B6���L:��Ӷ͵�_w-:�!ɻe���p�s�Ņ���-_렦�|�)�-�(��g>U�-J�ٶ�`�.�Y)�{Ϛ��o�H���� ds�w��
cP|؇;~N/�y:����Ӷ��$�e�eXG$�<%�CѠ4I_�~�`��L�s+M�#׀���l�����]2�Q�%ڢ�����H�~���(&�T��6%z�C~� �� t�[���85�t�LZ]�a�\F[y�����]�I�PH�C� �F6���͐[�e�?���Y��@�R�G=��:��މ�T ��h�Dp��̆�M4�#�w������c�U��e�[(5 ).=����K�ic��~)�@e9Hc�f�1IT�.?f���K�@����E�2�;b������NF'*�(�w�<��z�؎�A�](� ��8�z���F�A�z�pK����|�X ���/rBA���lg��ZA����{��������%x:,F�y�z�&K�Z��7i����$rks��f����X�ٱ��H�A�u��=`����I ��[S%��F�O%�/�h׵�������z:;{�A��?_6�1Ip)�:o��_k�r�@ M#�����*���n�������,V�b��g�R�����|���b����cr�47����ReI��7�g�YW��Y��1�:����oF;� R�z�䎘��&4���h$� �
D�C��=�m��qZ��;`�fg����r����3�W^�(�Y���	Q��+���=�2�~8��|&Ut�bӰP�~��[������Gth��'�5�\���������a6<��z�W�����n)m�C}Z:��bWQͨШ�Q���I���f<WV�27��/�H��n����MʞY�Z�6�	��
����20���?��Bl�p�oj~���*�\��Ӽ�/^�KqԮ�2��:D�K��E��E��3����� �2x^FL�-�^%m���8}C$ҪBk����"3�F������Pu��U쿨����c�2sSeG��8h����T��]���T�K���l.���VƋ}�I��L�`�U�d2����Uu��z&e�������`�kpv��/
=�d���ϬC��{A,B�e�ֈ��M1%�	3,�S D�mf����n��ԕ�&��\����fhy҈ك7�w��-�%d�|M��b�c��/K�9�d����&�_+�T�X�۾M$���o����"����+�	�?|��/���4)���@��К���!F�ɽ{�P�V�CN��`��D�9����9��{�:��6�,����;c��5���|M�&���_UX��B�nM{ѐ�Ŭ�Z ����w�7G�{��W�\fhv�U�c�hǰ�n��Ն"\�*O���L�t��ѭ!|�>i��c̓�=�c�X��z��z�_��Π�,ȱ�TGa���,W�!e��!Gz2�뜽����G��ff(8N�/�p�/�*�._��������<�s�����w���b^��|��5�*��d�%%ʸ��Y����)��p��06�B�l� ��gdW֜�ZY:ʅwőX�q�zi�������0k,*^��;�2TC�u#k�*e�\ծ��2��/�9)��S�E�|9n��>$ْU�\�9��e�ص��~�E��
�5���]���N�	�)��ӽnq��̟��&�1s������_a�iP���OX�8�Ѝ5�y$D�/��9�w]�YJ|=��r\4R�^�M�G%Ҟ�ϱ��i��X�A�C�td�ڵ��k�[11}��2�#�۫hⶭӕ�)�:ٞ��Ja] �,tQa��'�h��kRC��c � nQ���_[j�l���r�ϼW��'�������`�$��P���xg]��Kvu�d'�ױ&z�����8�ʘ��ƿU"�C�TĖ�hF~�����<�%nd%�K���&�2{r�dƴkI`cM8��9b5�0[���� f�c8jb�ٚ�m��v�"�6?���vM2숫�5�j���M
\���Dy�����H�����@�&�&2�B��u� n���q/#Q�ᑥ�Êv`TcX��K���� lel��;�N��v��t�N K�"/Xч���iB���{,���^�.�F�ka�Ri���Dp5�ƫ1�L@%�
�z���µ�j4;b�Y��Л=����x��F���l��L����=!��W��ث�
�
�	|@�� p��g�1 lJ��ʨȨ ڥ0�	JT����H�m���
��J#������ü������쭨Kf��w&�C{q>k(:d|������譔�ם��l��|�U��p#5JA�9A�O�S-�]K��Oz1w�9	m�U��=i���4ӑ�
�������5���pe!mVH����4[���ؽ4�p�B�
yn��f�cn��S��vdE&X	���P!��Z)����}Jt��P&�/L�E�<K��`~�]���_"ĶG�f �$���&�!K��q�6��7��.��|MŘ�ig�(υ7�ƱjɜvR?V�������$�G�A�͔�N;�5M�z�����|!��n��z���O6d2 �OG�cC�m#̬x��<�T ��ۉWt�|H��L�����}���m^�뮖���jX���
:�啉�|�E|��3����{����-5����-��o�J���Ұ�R���(����W�Sh������!Y�k]���,-�V�il*��$�.\��Ƭ�)�_�4[��`���T����Z��V�f������^0����$���d�q<G$�(�&\��VO��m}�e�w�"�3�`�O}h�}o�~���>IO%^�܏(�T.a�s'��A󳊯y�M�'o����W���,����-��D5��byC�r�b��QM%i�]0�V2} �$��m���bo�����?T��W�9�P���1���g�]&`��Q�}ܠ�#ٷQ�8Kș�h�
�
ά�2r��hT���ާ�������[�HS\����r9̐U/�ά���䢱������^�=���%2y��P?���}ѣ�q��Zo�:YyAM�6�_�~�+��Q�Q6��j��^��U�l%)^y{���"l�
LBAKF�g�Ǻ���O�z��q���!�\�)ب�(Fɤ:s�(O�n�,C�f�G<?i~���t�=*��na{~�kV!b"�a�	�j�0��`�ė?\��g<N�r�y�Pf�4���QP��1m�x�uU����knw�/��4�U^(xW=@0��tq,�8?z�ٷ#7uֈ��� �nj�/�Q��Ű[8`��%n8�E���f�a%�c��wۄUY[@q�N}ݬP}6cL&�)�,e|�`8�¾C��a?ˌ�|�S�� [�y�<�u��pB����l����V�S��9�"jp4�x�J8'?\�b�HW�&�N&G�.�#C�v6���x�,u�j~�UŠ���divb5ޱ�j� ��a>BpE��.�}����E>���u#%�|�?��|,� n�x�j�rQ��A�hY�]M��a�3�M�@[��V���Isg�xkL?����~��{`_�q��P��K����{�m^bq����c�K�&@pc<+��ݻYqR�������環�F�Ϯ#u���X#~�#�I�C�o:Զ{�hk���}��h��L�gdY�m����Q�
-���S�T10!k%e�H�MT��o���YT���B�e9؀��TrP�k;()C�\#��/�-s��_yȟ��VS!�%�O��ȋ7���hz~4`��E��P�h[�%mK�)?`J�vl�af�f�h�p��&���V�u#�:Z^�p����M'��C�T����h�JIb�ׄ�c�����cL'8��(��I���aQ�g�u@�j'�~5��6�{��56;'k����ڲK'�ғ�n�BF
�"[��~QYk,z����e��y�K�~����+k���̌����»ms�����bx�81|�`�Yb����I
���S����z��c��?у4;el�Q��Q%&�Bd��܍���%?�<Mo�:�b�q`DD+,�f/e;5������ oܰ�-ׯ"WN�������?n1:�3<��M�M�6R��b������\�gų�ױ��'Q*�ƎŅ����YC�U�&��D,I���u����!����~ո����Gd�z����?|�����~�X�����߇l��pR�������
8�k����
;s2rF7!L�J~?:���/�:I*C;P)��}���ߌ�v�~���0_�����#@��u}�(��������E?'Ю�*1��;�"�
��ڜL<�o�iϺ>����y���n�����IJ�}'z���>Ɣ*��h��Q=���/2�@�͟ǝ�� '�W���vSYJN�l:�j�� p��V�	֨���B5?y���"w�Y�٤�®�-C�FN� bf,)n`���m�])ǻn���Gt�K��lہ8h�p�hz(�˧7n�p���uS���B�gPg�p�����K]���˨
��N�g)d�����A����P��G�LjJ��0���r4Vd��������Μ����\P��e����j��6�3�d�Bc�v�p�H�� w��`M�o�ڥpG����@���jH	�\��1y:�B��TP�T���z��k�v��G��^�I*U��ϴ�n�(�!	{ӯ�j�g'�GxA��KTA����OI�ӕM���@Cai��D�$��F�ȧo߼V� /�9k��j�щj���Е�ks��݀���b>1}_X�~;Ջ�=r�h#E9.0ֆ�M.�d�.���d�FaF����A[��R��W�U؊%$ll��qƉD�u!��;)����d��wd�5�y��%��K!�'Դ �fJ�����K4/˘k�Å�������6Κ���e6�G��UM4�i��h���APk�x3.��D�>a	����A�6�M��!�q���z��D<.����5zc48I�(3�>?L�4:�Z��o�X��.�1����7TJh$�?� Wʐ܃O(��e>��du�tf ��9-��h��i+	H�oв1�eM,6�7���rK:$	���Uz1�|wfh��m*Q�=䙜�l6�e�lz�X���0�F��ap?l�ّ*�e��@���0����Z�J�7���~�A�^�@��vwc4�����#��/i�n�T\�����������d� 
ALs��50��qɻ<��їYOý�'\�E���<j;���[��]�C��	:�����V2oqxs���]^9����Ę����4J�������(ߘ�R�X�x=|�����ˋkڞ�,e�]r*�qACJ-6s���%��S��� X�J}���@���:��#��{Ƙ�;� {�A�s���k�7��Їf3IFY@�?o����ݺ�%r�����PF���Ԓ��+澷�`�&�?������(�Dö"9$!�,�@��G�u�.�^�q���U\���{q)�����<A� q� ���CD|pVc@��J+�c`�ߜW�)kR%;�M	��qC�d�)�6za�ڀ�a�<�)�q�?�+���2~!x�u1<|�3���d��������9�G^+Jh�%�n;ʧ���8���k����5�x��mxŷct�����">��\u[�4��	씾:�l��@�RԴ=<uf)����/�5�Ve�}["���uN�!E�Ҽ�q-����{.q̤iy�����)�C����m��:�ba�a)rz�.� �8��M�
�V�(�s�DU=���_p0t��ĥ� ͦ��t��3X�
�G�����%
VD��*Lh�7������w�,+Η
�8jՉ��������E��,[�F�N뭕�����@���k�$�\�nU/
Qm��e�m��b�>	C�h��,����t�����BIT>%���f��݉u�ްc���/��⏣F�Z��,->2�7�H� j��/�;��Kݷ�^b��d�]e���X�q)&�ϷY�&N�G1\3��$�����a�v�O�
y�'��8o_�ޞ����.�+��3���'�՘�L����^�\��2vi�#ʰ�c'1X�%�F#l�O�� �җ�������#�mBc��'���ds��<tS��b�~\��8�R�Ƴ��2�;�VEQ7��*{�����~�O
���)S�H�� ET���x�c�W/���V�sp�>�u:�U���(N�������� AO ��,�"x�W`䭡Z�Q�4��*����6/��*I9���uj����-�+���ql��$}�ܠ,Ji0!'g�$uSxש��h�?�y���o��H�e��T�����_Q�;�/�5��3��H��X��Q[n�i�	�{g��b0_�x�S~:	+���&�[<���!��v2��Î������_2b?���H��T �2�͓�~��F���3�k��:#��*�@��b�IA�c(O�C���54*;}�ݕ���q�#�]�.��q�M�c�z��� 	��,�>��Q������Ps%�2B�u�F��Q���T�0j�<�@ޣ¹�W�U����FD�cl��_y)_��༔[-��y�Q�#)XwXY��|��.�ޝ������m9��\|QE �=W�w�6��E����[Ĳ��e���ͨ������n1|�Cy�o:�ƪ+�<ױ��9dk��t7p��gvT5z�.����/�'u"au��x`ʹ��������'�7�iA�CUmWՕ�e��e�l�y�F"2xF�����5��Px �6?�����R-n,ZSt&i\�J�� �h��m��A3É�8@��KiS�gX���ˍ��?�?V���\5�_�Йv�|�\@[��x@����tVI��ɟJ}E�@dL@��۷�3+��_Cf�8�����D�Mo�\5CY��Lx՝�¼��V��ⓚ.�ض=���Z���0������k�/[E&�$B��v��η?j��#<��7(:�w�̦Ȥ����ѧձKͶ\hS������do�I��w��
�p��c�>�l�P
�<�$��{�L��R�k]��&"�0��	�#s�qi���\`Y@Q,�M�5�o�}�7�%�����G�t8aˑ�p��2��E�p���4	Y�l�ho�!yk��l�#xtS9��̬f~��m�,֫%n�"�4��yl���B��� F>�?3���C�&�Ō��OP
+��@�}���kT�!F�=V�fE�Zt��Q&����a���W�E�_m{����BO;/�u�a����\�/���?P04�Q��󴭩��������:�m\��^%����c'�`p(��d�㗭���s������f(�1ঌ?���\+��-�YO~���?~����`B�K9�jd����!���{zW|��ǳ�A~���N8l��`w[�c�I)���#�4R�z��<b�/$�89�m7��Pc�F�c-@�ȵ��f���m��a�w1i�ط/7�"s,]~]ѧ�@��uC��(yl�8
j.���t��)�N�@ ��<�����營��~|�;�=3�F�x�G�$����tF�����c�+B4|���sQ8�Y���$Kpn�s�F&����L�����1�d!��+~� �,�%�ZAѮa�+�@��h�� u�,�����u�8>v��dF�W��D��]aܾ;�hn=��IE'�<>��]�e�MĎ�e�=^�C�7Z��NC���\�pi�&��&$S��|��Rn(��<gQ�}iDv�d�h��Eg�=�� ��}6�5�_"v���w>y��q��^)�ew���ě���ZUқ,�>��y���q��L�ڷA@��|����������q�q���I��TAQ���c�=�)�ڐ8W� <���H&�2<]<�|.��)ψ��]*_��(S����j������L��4dw%-�
v廭�H��+b��iA��͖�` I듰���|G�������ꉑb��Ϭ���4
�n��p��X4d�� 	�.����ۋ�ͫ,����[]�\~~t �A@��_�=O�%��Jq,�P�N�i�U4�*���Jm���i�To�b`�f�<M9���oSc�o콆El��7d������6�dO������	�om	���g�u�}��D�߮��߻�k�Z%� `���%�z��.t��aI�t#��~p0I�<G�+üZ�X,"��
A�g)z�pZ���~O+�¿��$*��$�>�2�M�qż6�{���Se�^����|�Q9��v��5}��F�·V����.k��^��4�0h��i��K�^���T�,~痄�.l�L������E������]^/A+��w.@��8�QN�+Y+!�'��0A� =��b�Ty�T�3$�'rw�;%�!�j���0x+=]�|�`�Lm\������MF����(��[j\�=����`	R<vI�8�3���F��x��&�����=�3�q*��o�͌N$���[���y��-�C7ʮU0L�/�rH�t?��������W����hU�B��b+w�)_�M̫����(�j����{E@����o��Mh�d�ѓ@RvC��o�b�i����֬%\o�}wz�XԤ�y,e;�Э�b�����NZf�<���c�����3��N���%b���.��pw3E�-�+U�0V�	*5e����j�%,@pG���<�Fp����q���R�ƆX���^���Jq�lo�I�66��n.����$�UG��/���&B��k��f�;q��I����1�ˑ��gx�S4��������9����6)���۵<�������{�RN�����eO��%����ـ����n�}'�����f�$�yJ�t �G������C#���v�r�Ph���o� �<~8�����Y2=�:��L�HL-�KS���zl% �Ƽ�cfvdK��n�l-G��׳��œ�-�z��氞��*�Nx�O�p��pu	�^Q�P|U���1�H��c�S�V��]�O��b�7��cjوJl����\z�Rg�����QĢ��B,dUo�ofx�؟)>H�*�6G��k�*:�	FH��V��f��Y!����K}��4�Bd��`\���&DNJ;4���c���J��[M��oM�P�0��p�Jn�,��)��3�qs�\-u�[��ϠfݞM���O1�y$�Њ�1Z���@ŤQe%�9nRq�Í��B��҂���)k�S����;'�����Ǟ+�MW
�c�m�D�"�ɔ��, �ח�X�k��T����"�w�EYF�ŋN�����!��ӄ\G����m7��+�ϯ���#���f�ۅ�;�
��d�y��jWW���~�I��\��t�D�v^~��s.�+�g�TGx#��j��HĶC|-$�hQ��t�ͯ#=ξ����J����ݑJ*�Z1�[h�Qh_Zazͪ�M������M%9x] �C;t���wQ: ��d�U�<��*U��o��I�Uf���5�dK��a�������Yw�W�X:�:1=��x� Q��w#=�3*oO��p��C��rA}���T=��I,*UsO.�DP��bj��f9"o�ٺ���ۯc�aU(hY',���8���cF�-�o�r޻H:X���@+N�T�c�뽱��a��
�	�����5�l�- �[$܊�}5�~��Os�4N�Ss�Z�(`₶�(����f�M�"�yߟ�7�|X�0`��k��VB��Ƞa�H���2^�0��U�No�NMLaޞ������=칷�$XkF�o�j�2���E3�B��y�Ӻ�q��Xw��z��h�\�l;�8�xjdՆX.vΖ���e&���R��,	~���!Zk�ڝ�ב��{
ו�����K�UYc�SK���q�l5�>Fq�8D]�!~�RB�}$�im�Ru�V�a*isQ���:6��e��B�B���zr ]�A�{k��O���J��F?�4����w��O�"�\δ�w���C$�5��n�<�ζՁR��Doi��4UM|@����4�,1˟��%H�yQ�a�I�b0�J�s��/�_##w`&Z^ԁ�����9�x��\h)�:���5�MoT� ���R�	�%9�=��Lr��Z����c�6�w�W�4S��^�)��\�4w�PZ�� ��*�3|�'x��d;����t�Uj��f�dtd�P1��	���H_w��+�9�TK7T^\��oOe�p	�1���L�=�t�M�=ڝ/��/~��6cL=l����d�� 5�z۱nK&��^�W;}���]�I U
0	��W��z��/5G� �˙�8�����o�b�vJ�%3�������)kv��=`4�����d@��V:��r+�"�5�������DCL����9��E{�P|ӓ�+�'#�*��G��WZnV����w@�T�.5���z":�l��Rh�X횗j'J����(oI@tV�w�)Kq>�kr�y�y���E;T�vrs�^���R�`���A��7����?é�w��Ӈ��;&>�yy=��[Ts2����[x VN�̞��$�kʸ�z���Dg�t��F���\W��VlvJ@�^���B1�Rm�63򘣧W����p��_�)bI�O�>-���������e���ϊ9QQ�[Kfؑ{��@bC�٭�ʣ�ij���G��Vu�nL�H����3fH:dc��\S�RZ4��~w�7���J0D'���,R�!�n���4��/ZSu�q���d�Q
�F�2�tcH�,�sPȐ�2�w<���K�怟����g4K���9̿�0{�P�s5��l���wjfK���c���1ȼ�������綵��m{ȯX{N>�Pjt��C��KI�����_�h@.�8Xѳ� �:��r^5g��f�ҵQ�Z�ڐ��2�}�[�q���T�ړ��A,X{)z͑�����5yA%ːaPm��P���GM`��ݻ��a^�P���P)f�4VOU1���ϥ�>��k�-������~#ӵAt`c���v^)��P�w��l���M=�5JYRО�K�=�L<P �v-������;�sq��d�M�FJx��S�X
�ـ���eOt�@-e
��2zvq}t�6V�x��
Zy_���gV�(u�5���;�5�t��l�@�,(� "Ռ7���S>� ۹Rpo�a�&���>�����U���)�����eL�c#��^8(|�7DQ���xġ��W&��D��=�'^v�qV��{N�,ۮ�߬��dIc*���<M��逫�ߖ*�	_G�6�)�xE�pm�y.�.{��y��r+�r�_�]�F�m�U:�B!ꑟ�2x]��N��9��yb��7��jw���E���v3�cԭ����yq�k���l� �q�h��1��O���i�GL��l�N΢�]����"����YTyۥ8��jh���Ѵ0q%f��/��2�	��Wzm�m^J��ݫ�~�n��C����:82˖Ų��̛	A�@ҵ ���ї�{��L}�_3q��A��ݭ{_�~�Ĳ6f��8
��L���bM+�`	�7���7
HbWb�>�I�$�i�)�5�2A#��cӦO;�ו�AzQ������h���S�(�lS���T#�x2��@q�r��M�~�T(�����f��T&jMm�a˾nܐ#�:�Zh 8e���+���
�(���"�e�o�ʚ���]8[p2��o�W&��(������BG ��>n�������H�f��n/�8�GvW�O]��-�a��r2���~֬Q�d}�=�u?��y����L�v�Q��~�<���wB�LC���E�ڜK쒛T���\�e#������&;g<P=�\�@�ei"�e�Z�O�>(���y�(��˗��d*c������>5b�~~iC���f;����G�*���ʁ��	Y�XJ�a��4���M�(���*�u��ؼ���ތ�����U�yTWׯ��P
t�CQDj���G(��(k�P��q�'������Ёx	
�D�D/@1A��hl�_�#/[��{dD���3)!�ݹw����#�2$d���az�%�7��}5ddml�:��sGj9+&�v�d:���<r����e��������3)ϑ��х�
�j�ɀ	����˟5H�<�/QՏ�s1�0Y��O6�S���E
�|7�#3g��F7��9>��K��J�:Q7�~vܜ�Qr�ʏn6j�C���?�u�g]���{��7[��*���^}�8Oz�Q7;�~]�+FK�"	����6_�6}=�sQ�<�!�b�&�����ݺ:` n�t�|��ѱR�eҭ����cc���}�W��ajY�:Lr���2�E�| ݼUI��.mP"�X�^�u�`��
�m��y�sV���l�W�7�;�5u�.䧋���ҖK0ł��=���%���ۅ�� ��;u�5ns���)%��>���[d`]�!�G�ԩ�,�zCT�vԮ#uQ��]G#��!��r�s�u�gM)�zH2��B�tr�&K��k� �BD,�������������}����D�C��M�]�w6NcE�@@EN�Z��nZ}e�����iރbN��!٣fH�ѷ5>5^9�_����|�=Y���_���M��`lq��ˣ�Ph�U`>(��@�g揣�� �͉��t���Di���eQg
@�yR��@m�s j,/�!	(�uP�A� M�����zIV�	vɬ���O=�|�2$��;]C\��T���=Q�ji�9�i�T�"��	"��~ �߷�e+_���G�zW4�^�&숝�-\z��b�9���"��X��\ؚ������~���A��둸�=N����-�B:n2�����]|��x��s3�, גE{�I����{�M��ݒ�n����`���Z��z��q���_[.�6�䆴k#��n�n_�V��@�=����<n,E��W]�`!.��>3�t)s����b�`GZď���[�nʞ,�y�e4]I�Z��]~�L�6�2�W�9�{�<E�t8��[�:}-���XGgK=����r�8���o���>��l�3?�<Rt	�o�{������l_`����ƚ"T����^��|'\N�.Q�n�5 �Y�`�Σ>%��n��g?YFX\�RXc�A�]�n�IAW�����:����VHC.����ę��m�8fr?�NW�W�_�UE�v���z�H�q��F�9"�YK��ɜ�ը�Ͷ7��*_�"j�}[����k8'!��{�I�1K�O��¯X��/�+�!3#a��.�s/'�	�p�N�� �*(ӥN8�:l�8��5����Bw�%��,H�[3?,BL��z�;)�ճ�?��LK�3^�n��e���\C:'G�G�`�~��1�
����`���$K�t��eV1��\W�O�E�Vv�w��A����l=狿F#azQ������btA3��$ ��ޗL��KG���7�C��*Ɩ$�z"FZ[��^����tjy���X/O����G�z���sr�e����������A��c,J����)�q�u}�i��V����p'�Lh|�.�htnҲ��p��`0�/;�+�Q�ߞ_����]p���.0��a�K�1��X�;<ٳ�y������o��h�.�<����-&0m{�(M��с[��V��K9��z�3<��O�Xrf9�{�Ehȶ%���O͆�ZI�K�@�:H������Q�DŴ��>�h%���Cd?�˰U�����{�E�8���Ր���/�z��e9a��Phw��{�Kn:��P�䏽Lp���{g����D�Z�A�YTg�XD	\�/�������<�_�9u���_�F}���os?̓�u�bVK�ǖ^�|�8����Z��v���\�F�����j��E�@9����2	yt���a��݈pG9�ΗJg����;�� ���J]/A^.���?��W�0��Tm�p�������O�A�ƚ�K:$_�e�\	N�O�Ś����<:Lw�=m%��X��n��)/T�0�as�@s�\3c�u]���l�xt��W,��P@�^L$>v�p��;�[�?�u�汫���O�H��ʸC���t,�g�n��j����)\�M���z���3�!�W,��ؙ�\YH�e��g���A4��3(,iC�5Ƭ��{��ȘV7�;#�Yz�r�+��<v�Pܙ!mSVr$�(Y���nl�y �w��"�S�0��\����Ҿ]�4��~`e5mW���#?��5�Ae��E'_��boj��mY;"a�sNGGP���\)>�G�j{�"7����k|��og�3'p@�3q�(x�������%>,��#0J���EH���Ln�%.�)yc�X�_v|S�ef#�WQ���b|\�a��M���m�٘i>���{��0�):mJ�S���ʂ�$jU�
��:��8X���"��0��|�}�V�~(n���*ZԼ�8u�9m��3��� h�D� <�G8|Y�p}�[�i�����9t^��'���2�K>ײ�D�QLz�Ā�墂�j�K�� ���i��s�8 �5��n���E� �:���S$��-#���z+�܃�c�1[���li#���S��QA�?��Q/�/�����V�g����+��{w�%���'P\6�sƃ�h��G��U�3~�'���2�c�_Qy�D�������lϘ�Y�8!�U�zK{b贽	�[�E�Q�Y���>� o������V�q�@9a��߾:1Hp�%*�ή�����;�櫩�'�~����2�':���͞P8��W��Z��g$��rM��N������{Y������h
��?+ �����Zϵ�i�jV�i��c�g4�3�[S�,�w܀�V�N6�ʏ's�ar�E�ë�\�G\#���a�FJt(�ep�ջ.�b� xH9�7�m�>��Y�U�[��y��^�/��'���}���R�"Z��8�k1�V3
�{?ʬ�{j�-Lv���	�?-�Ȃ��I�>'{�S����}R쮘�Q<�`���w
�\mI+M����J�����������@��c*'s�VXS�M�x����s�v�F-�r�p^�t�Б�Q�v)����{~P�2����i
����q��d	���2�f���!����xzK ʺ�,U%|�+7��s�e�--�t�myh�����5ZR�M���N�P�˰Hf��i�f�YV�e�h~�BI1P^=^'��'<�`g��F�a#��G�Ɍ٥��%R�܉���u���#&Y?�!a}9^�2�9�{�R� ��!������i3z��W%��%I�.Ղ<T���F�bp���Hܞf]��������Ls�V�Qj�}�H¬`lfX�J	U0B��Y�dz5��p\��0p���_|����o�)�Ln��3I[�(��Q�4d��� �Й �@��c�7I�6W'H0��2��1��I&B�B��G$1Y��Y�4�k7�S��D�똜2Y��D�U�;FS5Ǌ�����.{�q��y�$���}MrٴYW��sUreN<��3[�%��ާ,T���$X۩�d�����z�۹4)�(UR����ɪPll�9J��4�o�:y�����E�P��?[���?�[%���|���n��i�6�jh���N��i&nҖ*�(�f�Fx_���Z[5��b&K�����2R>�G���.(UZ�=|�
e_��yh$:_�O�Oh�v����`ˇ���0�y��s�C�j�t��m!ږ!5_�gh���i�� Ԧ")"���/nk+�\��'��?s�?��3y�D���al���?�Z�o6�B���� \_��a��^D7K(�NB0H�Ģ]��/?�>����v�x��^:oS�R��=7a���C�w�<F2.3�$+S�7�7�OM���Z`�녺q��b.�=|:��K�
�*;[�U����;O@D��x�Þ|3t�����<�u��<F��ꉋ"ƻ��N��E���\�ҩ�;�Y.�L����4����{��W.1(p���&��_�p�s�V3�+��ǉ�'fy씲L����#��YoE聖TD0��.n�d-�h%*�7!�5#��.!�tr.ø<"�Q]� H�vs������}��t^	bJ�)�=*V�>�R�@n%���'X����o�Y�67*��+� p��%Y�����U������/'��qf-Bi����칛�1v�̯MW6N��H=̗���ꨕo�D�.s����r^�o�c|�)S���fΩ�w�)�V�7�ĵv�{9�(�v����m��u�#�s �O��+�@�?'���`�6��^3�:�ܸzp��I]������Q�4�/On)mt�+P����ƨ�o{o�=Vg�������lĘ)�=
�@G��u!�w��I�H����i����<R��7��EX�ovϙ�{'߷q�E�l��BCq���� pJ_�w�$0"�g��{���\d�J!z�����X.�5,
Z(o�s�t�lw�.1���Ј*���}�q�vf�����R���Yx99y:|Uq�����Փ�tuڳh7԰PX���-a�J�7��}8�cX�ےU�V�	�L`.I�mYWg�i�����.CݳUy�ަ跎���1bx�]���"����3�5��{��5��H ��L��s]�;�.8�g����׆�pF�.AA�F����}FvN_�*H���3�N��q7>y�I2И�a�}ۚ+��W����nS�;|
�o�K�R��;x&-��7en�n�S��H<��^��˞���a��0f%"�&C}���y�LifJ�VuC�
WH��[-uUDF1�Ԇ�Y�	z�ѷ���-1�ڧ>��>SII��P<�z!ׁ�;�L)D�����BzY6l�s�h�yDZ!��t��������ԗ)��^������1wp�,f5r>�h���N��M���uz����(�+xp���n1 -Gyo�Xh�:�0�Q>���'$?�M�U�0�߸��A<U�A�?i�O���^�as�-�o�O��i����-T�G�ƘVntD�3�<t�Fu���f���=	�w�V��^����Y9�}z�<�t�O��dzפ�P���tEKIC�U�!h��V�o���0}�h<��W��s�B�ńzf�1�_Z��� ��y�8  إT~Q���bp�J�+��Zp����]S�خ�.�����XHOc�U��~h��q#<R���0��&n�Z3i2qbü~qPw��H��F<Ü5Ďj�!DƿcO�w6�̊Zض�F�#@.+Sd�n�`"�_���1ff�<!f��8��0���͝��Є:O.R	n���{'��9�8� ����/<JjAϵ��#�e��8�S.BBߡ��k㯛�fFw�l{ʤ���;���Y3�E,'��B��?.Í��e$bx�1���NF�.7`�1�
/c�`���GP	�_��.�!�*��M��k?�֑��:�:6'�X\�h源���AQ����`Ф\�b� �5���7<���Jh��3�Ԣ5��(qL��a�)HD�M��:pBܒ:o��w��'Ƥ|��i��l����~&k��� �[ޣSt�����/�y�p��R*�E�{����eIt���{W�<^��������`;{`�o�i�_��g�d[�:��#���_*����.Z@���`��Ҙ�!�
^��n��ؽA�L���)f�����@|�ɟ��.~Q]|���H��>�)s,��L���~�Y+�a�.�r�0���������RZ^�T���&�q黳���J�;�q4o^L�m����h�6$���o+v�ʈtmS��|��c���������PjM�&�L���b�ߧ%��+���%�u��V���a�?�i�mXz[�ٗ�Zt�#ҕ���3W@�t!�ix�]�F-C;�k7V��	��9�Q�k��̮k���"��u���8����4�K��ln�����)1=`����� �BR� oL �C����V���Ѯ��q
��3�\��u)��(��נ�>,s�Թ�N��Dی��{%����ALM�DDb2˄
�
9�&�}O
��θ����T?�c������������m{L�P;���EoϕBy�C� ���`�p���裨T!h��Z�\��W&G�'��/����ώ�))���"i���
C@�WoP�2�m1�-ר ޱ��x0���[R�zYqT�j�k���?��Բe1��R�c}!�N�~,�����r�9��=�9���ո?�дJ1G��V���Z���kY�����g3;�¨E\�(�P��T'La�ͥ����hF3c�����N��D�U�R��(̫1�Kc�E�N@�tP�I�c�\�C�xR�e���(m���$���[�k���i؟);m򩋗�j�SN�>�SPVH��l]\�ި��I�!����������O����Џ�OWsχBj� ���vL������]�g�ۣ�<�R){����Q�ZY'?�dR�E&:*Ul���˃>9�j�`�OU��<��m�ڠ���Q�o$Ɲ ���I�e��2�ё�똎n����Ob�5�����9�rA�IK��H�����E��ܬ�ù����Q����癦��W�«��4S�;���������*�톮Љ��)�-
oBӳ���1�T_b{���g0O�Fϱ�-���K�����w�s<�q2��������G���[�E�9�M2�nڃ����n��Q *������s��h�3��ĶK2,�e>2EltS[�h�Nq����L��C�M���muX����(8D��&�!
%}����z�I��b:b�X=����á=��U���v�.�R���-�o�b;OD\�ޙ�E���N#Cǆ5��"��w��q�Gv�	�׬��'?�M�w�>��H�E�r�Z�����y%����d��Wk��@�j2s}��:r����۹[j�(��3��P4����q�?5`�R��5�������Ʀ4�]Gcx��j~&�� fl6o�<f�����x�9U�&���6��u��ȧ��(�OOώ&?�1[��9�NP[�E?�V	U]��uf���&���NO��'����饞���q�XgĽZ2�?d�G0�K���!d��������K˦l[�"a�����W/��{]�}����	Ǩ���P'"D4���@�$f�n<*R#	%Ǥp��N@f�+�y�k��3�oz�&HɥK䖙�gy�i�о�h�%/\U���P1c+<MeUJ�ϭ;�_BVG��w�Dtvdn���!���[���6���#��Y��u|컒B�����*�{S����jٍ���<�T�3pR�O�sր(u|��$J��<�'a����$�Bz�,k�̔<˺�5�K�^a�0�Y���DZ^�m$�.��;�f_{83��H���J�~�����x�<Rt69����?)P�%��tb��z4B)3�0����م�Y�`wy{B$�-�-���J�V��2�`٤�&�����<Ӧ�}�/�H��.ڬ�ƅ��~�q�`2z��irC��^���}�imP��
P�p��B�jN�s�F�l��yy��f�8� �~�}�P�Ó��K��,}�6v�w8�ъ��� � i�iyL�#����a�g���X�^g@�tF�};X��5Vvxͽ��]���N�Z�WQSK���-z�U�Br6=�&��Dm�_-��=uS��&�qo���K8�U�c
,ĭi��.��r�G�?���$��Ֆ���f�AS��Y�U;[�}/t��*o��:I��8�Vp5����Z�Uml& �`{�?�ow3 [�q~4��d�$N�l�6�x8	�Wc�B�e��k�����eDGb{�/�M=�%m\$ԉ�4N�.}U-����Vz��7ѵ��$�[/]���!B�hyM�t|��!�[b�n�1�9A	C���Y�0⃒%::��>ND\_��yA�O�9qa,��7�F��6AG�|
 z�n��JC�9�%���u�
.�g��՟�,	���|�[�?
�9.NÅ;.;�� b �b�=��h��Ӹ����iK��(��1sE�d��	��l*U'�h����=(��D���D��vBS�%x�
�K?���~�Eyo][�.}�G�M]!���soSw�l4g�͋�\x��lB��(�]ƛ��������Y�^�L�����k��*Ħ*P����M^�Al6}IN�0���-�B���R+|�7b�ۃ��WdߛY��i��c�>a�v/�.�������PhD];l<�<���������D��)�o���M(��,� uE����_�ߣD��_<������l	�MJ�H1��52Y���>�+/���!������47R+�L�� ��\�8}��\�#K�y�H6�#� �.�7r!g�E��/a�oٌ=�9^�_���!���C^�%S&j⒊S���"���)������c�}r1Fe���XxY)AcG{u-�V�e���M��yGƀ�\-44�Z������5~�QK��ob�T�8�٢{˔C4����)�Js���qG��6`06�3!��DmD����fe�<8И�G@u�a�Ϫ�`�ݽ:��ǜ�[��]̸����*e0=�-d����$�"�P.��i� S�(a�Q\:Y��Z�<#�_G�o�Ď�T.���������e���p��~��'=�ڄ���O1�y�q��3ݬTb#fdn ���z��u�=�.�j������i��%�z�v-a_�9�*��iĀ-� o/�S�3��>�,�W�vx3e�`�b 酕9_�l�%`U��@0ɽ��;���7�&�L�3���CD�1Ŋ���k�B�F�_y<K�6��
cVއB��c�;\�!������>��h��{&�]%���@�J�����y=^u��U��}��'�P�S��ב��ժ@+@��D�mO��n���|Ӛ:9�X�;R���:_�Ŏ��'x�����qrW<}��I,4��T��L���//ZO���+��|m�('܏��!��T�g�Z��d��~��.}p_*� 5H�UǺ�ٌ�]9P�0H�Idh�|��?�2�J�C��n�]���s�D�5 d��{?Q�5_��}p��T�7�T�'�>"\�Y���qid,���M.7��s��� �Ā>	�Į8��hn�&�J����s���PK�r�GG�x�y�t���(x|�?���ޞ@�.���50���&�l.�iP����z���-"5��������Q:�����hi󲯗Le{!UU�s���l�B� �2��)9���P���i���W����������Q���Uk��V'L���+�ɗ���/�sF[y|��Vuc6�O��s�C��/�q��C�tlx�����	:��:��&M��Ň*3���y��9��K�d3�oǜ@����� +N��X����ߣH�����&����=e;>G^k]���̥��h�*�Ԝl[�j����8\�Fљ�\]����
����n$ŋ�I֫(�s�DTk�y�eHS����c����2q�O������L�{�7�~mә���b�B��Nm�1
�FN��t��0�I�������X���=!{噸Y7A�g���'�D���f��I?�:�k�ghTԝ}nC��2�4��e�t��U�������Iw�$ϋ�ٳ3?Hf���Q-�v�����qِ������y��%��Ag];	*�%x���pJa+��B0��$���:��,DD�