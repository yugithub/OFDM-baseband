��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛx&�NP�/��/��M�Џ���ˇ�5�]y:}�*Y,Ř���F��N6`�|4�����r����a/�T�Ո���l�A~��A�\Zp3��xwI�"�ڴ�͖Zke.Wr�}�u�g������j��1����шb��sQp+��n 늰E9)3�eQYU��P7"jl�(N�S�VUn�i�G��Qc����_�©���i���Z��91�h
)x�����t-lBo��g�R_���ҙ��\}����Tꁀ���e�v<�Y�}r(-,�@'?Y�#,}r���ƃN��M4�^tF�*i��ԭT��O������o(|q4��:Gx`[��PÌA�ٻQa��a�<'��ف�]�S�P�:�5o3v��80���K�����ٯ����H1�8J�h��lͿz����?:��f��I�m
��x�LP΁�d^��WN`hỪ,D��}��Qr5�T2<�L��0���Q�M_-\6>i�sBD_�r�d�NI��
���f�볇M+��j3���4I�h��e�x]����Q���Q�X8G�z��yUu�$ٍ��!.�Udm����;7œ�O��Gh�Ѩ>��S��#2��ug<ؘ@IԬcZ��	�v�]���J��o|8���~���4#>	R<˳^�ư������\l�-�B �	�?��2���$��-�A�17}bĐ%4
.K\�evqL\ Ϝ�����B10�͗�G!d��~��0�S� �����m�@�f�A��YLxnn��M*�62Z�Kn�钆-�[�8�F੏��C�;JyA>�h*J�wBoY�w>��g)�Vn���8]}3>�nu���AX:!��ďw�9��Kl���޼�ﳂ��q=�\�R[�)\��o?;�2G	p51l�]܎����p~B�'�h�%t��M��G^o�o��oe���TkѾl��)lH(��!d0�Y��_9��n��Ц�ǧ�9�a�2�������0ĒT�H���@�h*R�$��&X���y�Km��j���Ӵ��]�lw��J)�]b�E�d(>�K��cƥ��q�<=�v�.����ȍ��\c��7b���M��z�&�6ׅ@2���d �T}��l�!E}��O\oz��+�>�K@8nH���"��Ho���*y��| a�Wӵ!~zK{��i
�g*��BW��~�k'ssp�|�2ɛ�ޣZX�ݔY���|���o��5� �����jGl	Y�9��s�� �c�/����$��8_K&���Ji麫i��2=�]�l���[#i�W�Q�U�ϲ�O��<���m���8���k��)�z��	)�C^z��Z�P?m0xz�V�7���>=r���s&X��bTQC�#)2O�^���/�b/S�����!&�}P�w�������ϗkr�2�L�Mkc���H�Y��J�k�ݾ����8�Q�<����@���Ep�D�w.7e�v�|'.��؝�	�ɗ�o��I��w����L�oo��"��4V�6SI"<[�n4�Re#��h׃ߊ�Ū�W)h6�G�4�\?$4�����%<4#��w=�{;�zPI����^-ʳ|M��&��~��
K�"��S5���`�R��Xg=�`p畛G�R�gM�o om�ɽ�F��Y�*���/sc )D��y�����rwh���bjPI�6���<M�4�#"̉z& ��9��*������/YGW��&�ƚ���]*��ѠA�	����^R/+�q�w�-/����t����4e뭩~�tRk
�b�� ���!E�+�;	�fkzm�ݛ�Lx@��Q���(�H����6�E�M����G@��+��U�~p6ecG��h��P.�y�c�q@��X4�