��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�؆q/�֜�x���K6�"
Z����.��E���i�>a%�y��I��6��z}�n5�@���{�Q~B�J}���%"d�e7�����������s�&|I����P���
�<��g hR����tm
��6�Sa(�W.EC���|� /��د��E�[��;��'�X���d)19w��G��K���xO�$��Ԩ^����-h�`��m�g8zh�f������>lَ�l.-��LRaHb�{?o�/��f�Z����e�b�]vEj�����h�lC�O�[�2!cGf�)˗��-m�����J����L'vVk�u�Eԓ^9�G��Kn�z���o��|�;Ӟg�;��=�W���($�i]�6�6%H�sA�����3�Y 9K�T\�)r~5<��-@��=|s���7$�������"QÌ�W�D����L�Y��
���� `�Bn�i"O��M;i�xf0p����TT��{.��-�h�
�X���ٛ)WYc�ꞽְ���ݷr����7�+k���qpA
�&�P���]@X�l���jMش�{�������;5�8^h�%N6ǫ���\6i�2Ś�r&I������?.-T����iƾ^�F�":���s� oY� Q�\W��8�%����� �σ����-}|
�#���V ���)D@�n��l�֙�T�8@���O���D�[���� +�*�]��K�@˒
}��,�X��X���D�������;�O�F�{�*Ĥ,�����U1L��A��*6|����Pu�L����Fz�������J	�\g��U�aWVIJ6Ӣ����mEOs�߁�ھ��C�#|fh�,�ME�\�k��jS4sEOw����ّ���`'��Q��{�q�"�?��p�5���xc�����R��W5���?ǈ,Ï��#��(��xk��S��oJ�7�I�����JJ��m5�R����*d�ϙ^Y�Θ�9��
��߱;��;���r5i"����'U���J�R��֙�Yn��+�'7]��q��f����)��c����P����l1��S��F��;���C����nzM>���Nh �;�.���C7��Ă��b@.Z�|(R��Љ|������HXi�<`F��|v�ӁUٙ����31���Lmar���?��R[0�~�_9Y�n�!���0������Ƨ�jn���6E��M��5tx��q�'qH��ZB���|G.���a�&�)/�Q�	�R[���(��3ɨ�--r"3j~I�Bh:40%��=��lܪF�j��4*��}�5��[���{s�g��D�����k˥~�5Z��߱�;Z�([�x�鷥�ӴV�F��~�f�[�Ca�jmzSf]�έ�_>G�e�+��fy�V,d��c����n����)����l�%�cO6�a2��+��B!�s��-����j�ư�ِ:��)�[#1x(�;��m��V�^�\] @�Q����ox�Ia!ݷr]�Y���L��Ȯ�e%(�B��5�>��b��?��NiOvd��K(�d�͚m�Ʀ�?��d�#�ȾȻ���ػڬ�<D��N�j���Y؇s~�|�5����F9	�G�)#�9���W��$@��)}��`�ʗ-�'g+H,S<�EL�$���*���ӳ�:s�*p�ߏ�F��1u��U�.W_�Z��,ĚV7����O�����
�JU���%.zt��*^D��)杖aI��w�d��D�ܳC2s
� ��=��ț�#Y\n�k�Ֆ��->;?��Kf����d��r�E�y�N���%�^hJ�v���7�do�A�����/��C�A�Yqk�E��`�ض��[�K��^��HX���aG�"#��ԮKm��X�2�S��[�$g饠zE�o��Zv���U���xg�OM[?��Id�P�	@��18��2��`=�>/M��
��D�G�� f�:G�X�*�Ԏ<�o�&Q�,G��ËZ]�Z� v���}�7�cJ�BX ��n ��0��мE'3y�o�Z�e\`�yv:,5�Lx[�z�&w	?c��`]���'�F4p�\�&��������X�BU<��8"� "s��c�YKџ7��܅����(��܀PZ��.t��Ŀ���d�<)�l�׫�W
`.���!N!�;�����&E~F{}�oր�ߤ΂4L_��D�UI�J�&5?�v�
��`�5�x�֚�/l�)Mχ�%���'x�Ƶ0���>[ኀp��H��BI�q;2m�njU�Sgn+ë����� �*ͷ��H��;�M����hq�w?'X]���K�4�{�ٯ��6?7�>�T�5=�+��-?Z��$�%�R�`̕����cJ����aU%2����MF�K�(��x���5B��x�� ������	���vjP���>+�|�Omҽv����r�L]}�N�hA_n��_�<m�A���"��IM2D��n�1hwta�
���ܶ�O,iL]:��ܚ�L7 �h��q����7�m5� H�MV��.�����j�� �� ����Ɖ`��q*w���ֳ_7����N���Ǻ����f�E�j����e_��2\��%ֳ˞�FύC��~w�$f�ֆ�a?�Y�6P�{Q� �6l���$�莹گB�'7Lu��T��N�l���۾�9sQ��t��.�A�eeI�.og6~x���b2  q ;�>�q����^���&�v>�_!ވ��y�Z��oԯ�����$�M=,�@W�œ�k���(P��!66�1Z��v��F��|ZNi�/�T�B2��#�Ʒ���2�"��_�����n�i����QX��w<k���Tɭ�Y����W
�n� �b+1��x'���aK��F�Y��{�ɗP5��<ȣ$��w�njwR��=�Qr�o]F�5KX;�	�Ve4H�N�Q��c���ґ��[�p�BU���(P*"zZ���}
>V(�ݚ�NX�H|���}j�Q��ٿ�3�*��Xc6T�G|�+�.���.��$ ����8��=6JB��0�ҫջE���#���Gs�ل��vi7eMZ�k��_NWc51�zc�� c:�h#�+�������K���,I~9�;jȞ�7s�h�qDwr����U�K��pG'F�~@Yf�W#��V9�?A�����&��5���%�	я��l�D����� ����$.�|��/䥕[u�ve���1�bк8�����nl��-T�X߳�Ӑ��xr	rXV���J-$�Hh�����V;}���H�w(�Cv����s�#�8�X����)��^�Ը�bo`���+8��Q�"J�	�}�_c�ԑQ �����?��0x@�ݏHÒ"/���� u]�P*P��Kĳ�5��<"j�v� �p�ԋ��>��0�v�����?�Kd�K��ڠ[<_ف��jW�,DG��_�]�<���/v-�L!h�v�ص�` ���  /G�W���C����[N�JC�A�i�����:k���D��,�+e���| vӲ���&���>�� ~)��_A�ap�l��D���?���5�u�Ao�1dO�6pdP�+���F'ӝ�l���e����O;#g�Nc���z��I���2��w�'<s��X� ��G�i6!ƙ �L5��&T���~Ua�,7>����ov�ٮ/��W��k�� U���
�jl��k��c�9��٪�J�{��)��:�E 'j-)����fC���ٜQ��zD����@}Q��|�2����1z٨��b�X��+���|��"��#��,r���!��~�����:T 8�lC�9Ҿ��KA���6i/vkV�&�)#�	J׫H1�*x�~ixO_�;���&I_[z���ϑ�������+�P�w;nZ^SJ�Je* xH��/*���Zz� *}���g�;}�$\:�k
%�i+l�KcO$��o��8��k�h7�����ƚ���L7���n���"���`�^S�L٤�+(qd���(|�Q-�p���v[�^�ZTB,��B��栩���7v
�!qQ�p{�Q�Uo��}�����5�����\��H�K��M5���?�A��ctzAh8����1ѡ�Alu��M��,N�bɱH�Uݾ9�ɳ&��x�H!Z�m���G܍a��s�V�ܫw\�R[B��mY�%�@��_A^$K��6<���S�롈�	[0��І~��rMr�z��G
�o�{�`�%L�>;�/�p� ���{��˔�P�CH+��ެ�4���y��
8εϩCaM� ��>���@E&����
����q�̈Lֵ��2LX��k��^IJ먣�B���N�cM��?^]њ}�tN���VB�C�bhn�&U��J�*��cO�@^b�R�\{����� z�0���o$�b@Ӗ�%��j��uH�V֒�M�p��ht��j�5��G}��&΋۾�ܩ�6F���Ux��L	�00�:��(7�*�b����3��u#*�P�Y�qF���&=�YH�BVH���I"-Y\'j��b?#g� d���h�8C*;���w���H�:�=88�̚�/ ݇@	;�H��Oxk�i[��9�f�$��ف`\�4��Vk�c=�hD�������).d��/�	n�����e�(�Yw�#������ې�u�~#�K2('�=��r����J5��	�nI��R���7]fRj8�:�-Ж�O�Al$1n]���W"�|�y+Y����G�#�`gx"�@t\&EZ8�ׄ����K1E��V!�It����׸�Ht4�F �($�0��4ܡ�嫫[iw2ĠAj.$� P�ix�
���\0����x8��y�mP<��.z���)�6�����tjs2ڻ�\"�V��?2�
K��;��lv�-�kq�b�׮p�t�u�D��U�P��ܭ���B���w)q�@���	e~+M�0M��[`A�T���{2{6Nו@�>�S�a��h&}*O����mJ<�D�����Ԥԅ�'���d�1b�!`Q�;5�^;�kf�֋l���46���S��k���&ધ���ז��x~�i��=7�X�`-̓��πvi��ƝO)h���!3�Rߜah���=S!���(�2z�([k��t<��g*�e�hu ��>7[�f����󇥋��~Z���|.�fO�!��""�a\:DQ�<����fΒKr�RZ37�x��Q����oVL]�9K�j�}��3�GBn�|/����s$�H+�¢��$�D�Iڽ��� "H��z��V.V�\t�vH%�.�6Y��X��m�ǣY9k$
�C�?��������ԑ)|�-�4o
r����u�W��V�i���7b�
X����"N�� �fC��<�gF�$xz��[���q،����.j6����������"��z��>���×RI��4��E)rͻ�S<zX%�v��:�"��^\��������D0(<a���i��W) )����9����׮i�<T⟟<��Q6YBK�Kx����s}>���c� �X�C"ˊ�+ծN+����)���A�,��&�"B��kuK
��:*�'``�wdo�QݠS��{G �ߊߒ	N�|BB0�Yop)ō��|yM<Q�I���j����XR����YA�x��{��[B�|��:r��Po�������e6?G�D"�z���*�
e��d�u�M3��G���UU?�9�Rg�j��M�E*p#��3�9~�,�6�Sv�����G�Ouk����ߜaP��ƪ���� ���Js̄��cfx��ɚ\&hmٗ�̉���_��w"}�h�VK��� K@�c6ؕ��z��y�Ji���"�?@�_����b���Ɠ�`X�&�_}�Up<�[��_��*Owغ_� ?ݹз�\P�S>=��o�7#OJ&��$�(���(%�W�(�9	��B��k�!�����T��1D}��~`�eAd�3���k1zp������Hݴ��ZM@f����,���I�y���<n���'`�P@�?�"�b!�3s<���=iGZ8��1�P.[�x�Q���=������^�)�P���p�9n�7U ���^��Λ=R{d����7#�-j�V �?k*UI���/9Q�s�(VN'Gã��U��+�� ۺ��#��E!���Q�$����v����Eđ�ZK�����W�u�� �����o�K��g�y����>X�A�AP궘y4`�֘}�X�o�y�U��wK���¶9Dkb'��.k�E����E���h�Bql���k,eJhhv�ݲ�QW�����3,�-I	eϨ�i���>L��>�*�q�;�(��~'ˍ��ң�;����a�B�f��jq샤ʏ�oy6���4��i�4U|�d�>��ìwI"��(%7��t�P6��0�rgB�CTLh���n��*i9'��	�w�
�����V$J�(W|�W	��P��E���Ƭ��蟤�^�'��{�$��o���7�O�Ҫ�Og7�:�=�6��L�~�1'U9!�Κ5��m���5c�\�Li�*@����t#�@Nm�^BDF�a7��Ec��ݟ3���%֓$��-8QgP�)����1;�r�����dW���7��� �����z���s2E�&ٷ]x�zQ�=����6�dc��8�����Ivg�wK��/ʆH���`��+�P�A5}�)�A��z+!���e��ߕKX�1k/�"o����S�^��k Z5c��bQC-q�[ b�5�r׿��Ԣ�&9���A�&E�gB���g�G1���Q^.x�C����-����W�x����"�BW��e�� �����"��ds$����|ҽE4���y�_��c�Q�pǼl<{�6�T	��:I3`u$�p��?^s��ݟ�}�� �����%h���!,t�� ��|C}���8�����i��gh×wDvё�봋�o�w%�ԩ�0�j'�J�"�<�������CE�?��(���I�Ä�O8[au����f�<�g�n [��I�q�z�YluqM��GH�i���-�# �"�
á{S�"�W���LjǨh}�(�/��"��L�q�{��l���m��nޗI#ˡ��ɛd5ݦiz�>�|����vs�Nӥv-"�w�9]N���cP7<f�Ѽ��H{���<�	��1Ͷ�F���Q&Qe.A�'��g�o��皫Y?◨؋)N;�8 ��^y�����Pl������s���9xul�
k�w����(o��}M���ַ�#eK��i���5�v�>�^����[�ӡX,h'r�l�[��&'���B���'�I���g,����>3*2���[��~�P.r�˘���XeY���F�𹂝#<X���o���ۤe�n�A�v��/��A�沇�g��C�?�G1S�Y x��M��-�1�,.�e�,��e��S�U
(9�/�t,Oa��1K%�E*�:6p�m	�©�`�Ux���{�D㐁�]"�ި?)jrev�~�������A��BǇ�o3�����^����v)�1<�!��#��U�o�c�ħ� �����\R\�3]:�BS�ݰ�B)��O-�n�s��oC����m�GLn|�᪽H��Zh\R����O\oo�`p˲&φ}�a�8��Û�2 �
��\���dp��-S��	�
v�-�r�yy��3��8y�|�1K��2?�ԫ��a^t�4�Ձ%J*�_��Џ֛)T� ν �rq)�gU���A�升Br��|)��Wi���RJ�<.��T�*�M�.àG�3x�nG��q2y���,,�+]�"��P��NݺPO�i@�5��0���G��D"�"�60:�e;S ��� 1��xm���������xΓ����[�D9$�|�R;B3�e�5)�}9�&��K���v-�*X��)*�#��!�_��@&��ߌb̉�3�o�z��A_���Ìw�Y�@�F��/( ���,�2S"���{���b�y��{�s��#F������/�y7R!���43���f4D�=�1�*[5=�͠�`j8�g3����% �n5;Y���.�Š�/�4~�1������{�����Y���e&�HL��3�2�XN #�T�T�a�j�q�|gP��k���8@����A\��g}R
�"ͿN����Kg7��XD�*H����EIh��t��3gFӇ:{|Ȯ�ICa�C!�f��.
�u Qpd٪�j68+�H���0� �m'Q���U�o�H�>�����6;u�7��ق��Z;�?��
}�	 �SoX�N-dl�r��\��c!���4ǭ���6]ۋ�C^8)��^f׭[b����K/��ͩ��͔xh�k
�M�r������1�:�w�Ȑ�*�qQ�I����{��A���__�jY�������]'���Q�]�$�Z?����k���� Ϛ� �x���=��ϑ�޶�qԀ�����bN�ԣ�_��Q�3]��b?Ӯ6Kn�"!Uw�#��x����-S�g#B����ٱk�$��\^��c/��E�e�5�H�����#��ﻗHx�u��e� ��_}��D3=EjC�@ˤ�k_q6�Aa>
-?�o:6U�%k��N�O@���0��2J�{����9��Ҷ��|��p�g�֦�`�!�f���X/�λ�H:�!#AMh��Q]K�[��e��I�ejW�>;�|�|f�.2Խ�ނ����ՏV����tV[�C����R�t�YMB��I�\L�c9]�
zJ���]�Y8��%�/l��aODT���̨��y�~��	�J|GO���m�7���BP��{M`��J.8.���
U�[�[ͨOg����2�&T�-u��DvyJ�+7w�/Y$/�b�i3@�:�j���ꖸ�<&�C�������fkZ6�7�����n�CF�"}X z�帤��Q[����i�@`~CW�֠���T@z @^y,"a0'���|������m�K٩�}K�^ƹ�y�+��=�!�ȗ�dUqlD��[�
)�eԆ��זI�;W�����,�i�$�}b���q�W����@ť��������M�*{��U���=�|�C�dh�1YП"�����!a�K�Z�5-4�*�v:b��Gb�C�Ӑ�U{cDڈͱݪ�����Sc>wL�.O���ʧg�{�|��?��I6�[��-���Q �]��:��/�8g#X�7/�)�F�R��f`2ӯ~z����;�<�ȆlJ�Ȑr��t�7�J�T!��'�q^=����1cg�M3\������
@>�N���X�&��}6���(�7���^Qε�"t��2���xw���A�oB��@݌���k$_9�*}K��U�W>h���	w�'Tb�YP�F�y� �B2�6�G�J���[N�_@o��o�~�{��}�r�(���TG���/�<���mp�(�n����ݚ�9�/�ym]�����9�Z\��
o�{�ȁ�]h�M�e��o$6�U����Ǭ���2��) 0�'���9���v�����F�@Ү������}%n���J�<| 5d�}� �$�kr��f��9/��C��ΰK�'�`D���U�#��4�4�(���4��C���,_�ı�
%;��Wý�A���aC��	�ۆ��Ӊ�/q1$r��2/�)'�dȤF8F�{�-�� 3�A}�X6�θ�ε��63�.��d�-�si+Y���~��M���ǌ�DSq޳��`�ww���u�	����дy�a���v��g$��"L:謴p�h���X�HL�;�݇�-C^����Ո��R���,��[��9�]�G49h�O�<3���ȷ�Y�p*ƍ�FT�
4t��>�������?�ָk��̹"�	m�f7D�Ć�E�!�F: �һ�!��}2�㶒T����;6k(H�[f�w4P�su���]S ���.��X,ҤbD�ή>�eG-E�/���,+3�N�<^���	��	�´�28D�D,�����Z�԰PJb6�j�>�Zq�-i?�n��J������S�(��i����|n�`Ǒ�b� Bz
�
jV����b貥(�m���9��έG�����[oAL?����E[��T�]c��>����� %z:?u�X��$�	����O��;��n���^Q�ĸ"�>���XcQ������Uc�� $�㝿h�d`�=L�%-j�)�ނP�.�����6���y�������ah���:{�Sֽ.�;H���6�!��*�n�R�s��Qsv�Gbh�\�p'nӍh��MYbf�R�A-P���ݯC�z@4IƷ�	�>j�A�{�'��[�?�X �ӆA�N
.�~ת����~�+X>��)��ҳ(��d���A/%���Ҡ"�G������Xg,h�;>	�6�k� yjvT��!.���e{,E� %"������;LȦ���ʀ��ƪ&#�Bˀ1�G����ug��(f}Q��u|< ���2.�FWI����v&�RW�R�=oG�3��1�\�v�|LpC7Bz.�����>[�&�sV����X�u5&���+h#n��>���{��?0�,�JCBɇkl��*lr��u�C�w2��M+������O����
K#Æ}@�fz�L���wU3�<1$W�|��h
VZځJ����U_��<���#���Z�F\'�;�KI5�'��jY�u�w5~��cG��#Mc4�."D��a��Q:�Mg2)y�b=[�5�-����z�q�_��h����|v癗\ϲ��Ĩ�~5Xk���K~u�_yqǄ�?�O\q`�Ƨ.�����m����wmȬ+y:T��K{T�S൜�"��9Xp
�E�/���D*��G�/]ӭO4	c]��GH�sT���̚>��6t�VB\>��B'8B��E��N�)�\��a����CL>]`�M����I0CШ�|W�6�i��X�p �!0�)ڤ��wNJ}U��2���n�N����`zc+�š�"��
�ƚ.j���d��r�PW��m�y%�v-�b
,HY�"�W�%��\bM}��,�XrYxF�u���cDO�/u���������v2�֓R������<�0p�-a5p2��Q蛦*�5��{�C�m��H�2u!p��Ҡ#�gwb+-ĳԃ�92i���p���` i"ʔ���e�խ9�{��»Ƴ-`�\u�F�j�o\���r<c��g�LF\TURq�	Ci�9��N����S����������:Q������~-�I-��$�s �������HQq\�^ x֯�G�F>����J����N�5$�����})��(��BQǏ�F�j�29|:PO&l>��,��U��s�+�BT���1�:�Ě��p��?{����B�y4Q�C�W1�._��33؉`��"�� ���$���!wZX��Y��3���x�JhҊ�4Bt�G����N���^Ƅ�_���%a�ხ�(�&�g%Rs�vG�γ��?�-ϵ��m�M����w�o�h���T����,A����@��l�.�������`��68Sč@d}��4��](k��U嶈%�m�܂��x�����X}��
jy��� 2�;�ցЏ,�w,
�w�V�|L�Q��Z�W�V�kF
�(CI_�7�W������HT��Ĺ���B|�)�0���4	$��������ӲMqtS���#����k�IY�JUC�O�$#�4R�T>���d�5]M�.�E��6��u�@�罨 М��FZ��SB�Wƍ�ow褪���k��R\�Ѣl2eƙp����^��p�����a�s�
;έ4�[�|ꉕ�%⇽B��{Aފ9`�EF�eN��6Eb(;yذ��*��<�Z&��LS����xL������] gEr��j��̶G4�`A���3]ۅ�Z�/����T��P�o|��@��U�t��N��B��
n�:�������}���B��m�*�։��7��&�TVԋ܉�,�3lY��g�F�/}���z�|�隫4���&=Jn/�� ��4��7Q(�ܗ��ް���C���ͧC���xf����������䵨Y#�7C�li�g��*u�e�Hv$���*��`���r����|-��{8L�&��bja��1SpO���CR;����<�i&q#?��e:j��4�R�k	+e{7B��ܨ
�j�!$;��t�34���s*�U�ౡwjl2����G�,!x%�r�/V[ Y/�Wd�n��:��ھ1zN��q_g����2�ⲓ���z�&�EJJ:������t�/n�םN7�l�ۿ��Jwy���$�Q�*�A���N���Q��-�|��W*�;�wI,ﺨ��be'cu�?�IYA�-wj��N��� � ���Ԟ���3�pA�6��M+j'�Uo���V��^$]�gC�Ե�g9�vӻ�~�q��."��	GD^���v�[��cM+�!��	��pV���>��@�b�<M��Gb�+2�Rx�#��'����0�EB�2��?�,��4bf9��\@��� ג�)d�;ɨ�ޥ���w�I��^(���Й�u�|Ì1Gg%��	^55M�����5K���-ۑ������0�T�:ڈ��o�_�#t����%l�GoL��E5��ޕ���9T4^  ����2��]��i�?`�+���V}����/��yb@Q�xMD�z�M�	���<!JT��
&ܱ���@*��a4��`Gk�p��Ѧ�Bn��b[S.<���EE߶M%��(KddC���I�+��~�� ��2
J�&��Plk�Lw ��}3�De�tD�Wg�|5�*#���q(e���XV�{��Ǻ;�N*J$'�ތ��*ὗ3)���4�QڡT%�k������T@4lUf|S��7Ш��j/�>�F���e+}PZC��|��N����Ć���wꝑL��8����Q��QAn%P��>E)�pϨ�~7��g���aQ.i�c!�k�kt��2���\�H���-{_��Etx��A.��r�/v�|t��Q��� 񍗝��`�$#..���zvu�Ȣ�d+S�/O�"���	VC��#�(;���	)Ǡ5�'�h���	��n㒞aۧ�r%c{\��M��~ڐ�]���d*&?MHJ�����v&�OM�u�b
	�uL���hE��^ya%�>'��C��2�,eV�Ty���%���<�aUG�����j�NX9 %���Yu���o�~��:n��qj������9�]l
$LA����PA�>mU�;�Ш#�&}�κ��0Wå��'M']�9�ۭ��ƓE�*�g����LH|��,l75�s|�Adp&NK�{�Y[�m��!g��mg���P�[Y�{f�NF�Ɯ�t��Y{��,��x����y��5*��wEh|�z��`�5�z�'���2��Ӛ��{7-���S�����Hv�y�����+
�w�+i���zG���H�e�{�mN�'Xj��e�JI����{6 �O;��]ƪ� ��n5���e+�jv��-P��O�e�x<�Xa:_ d3�=k�G�8��O�\��_��S�ǂ�� 0h��	,\��Tm4:��t�mV�}H��{0ܩGm�o��V��>��8���`��/�V���o��΁�_�3i]�-���q�'U8�/�َq-%}��δ�6?�5�}�ѡ��� ��������լC=ˡK�Mi��Zn�BV�.��5>H���ll�fN�jV� �eOJK�7����յ8S�JJ1[��Ljp�,���~���:𞂨�v��ŉ�z�fD��Q����@����DNR�ȯ�҅���d�G����������}�F�,r�-��&����P�=7�ԙ�����]p\�ps�X��꿓D� ���\d��< �͘{�դ �X ���WK������h�`�/"s�!�xtTDx�m�
>ws���8Q#.���!����ڨ�	����4
^�cE+(��p� u{�!�Γ�B���(�L��JR���w��,�*�-�q�̞��?�C�lݗ�Լ��`7��ql��`��0�4v�p��$����U슛��ڹs��8��X��lg֮d�z,�����9@}�?�7,�⯓R,��ʐ��ӼO��bF.xpu��,��U
�B1��̮b�Kr�p{\M_�%j���$<^�{�D>�5,
A�1F�W<�3~,�o�"�Hs<����;��O�V�I�,���6�ۣ�=���9�:�k�\�@�&b-0�o�kh&⽞�*k��11xs���>W�/�8�A�;%Ǟ0�>��߉�a:y�j�	�i�X/O��b�y�-]�%��l{;�=p�&?9�l$��bB�d��Y�Ltu�$�B	�������u��|O����?��֑��Y!��X�N� �1$R���]o�����wp�γ�Hg9��\̳q�~�B��M�Q�����x����+`�:t��s;�! ��.�֌�����#��;o�$��Z�6f;e-#�Qn;���Gt�Y� x�u��M�0?��Un>Ӥ�@��>냞��BVJ� �Z��@���7�8qD��Z�zv��//LT]�k�����R��ջъ�@*�{�yU����AY����R��V���z�B��x��;�)p�8ێ����դ؏�U�@���k����NHw?nI�.�����x
7�,����h4Y����C�(��K�����kZ��(n,�}����D��}ף��r�L7�]�䨧ETR$V�+Y�$
��c=y��e�1וr��V��z��a�S@(:�r]p�*�v{n��Lz�,c��{\��=����Xm�ŖX3)�m���,��*/��O��qh	-�t���ʲ��LOd�
��b���_�ٱ�c�I�8v�������C�9���Q�|lX$��Rf�$"7�]���w	�R��q@O
��7+㤎����ֽ�*;s`˓�S�>�kc���F[ܵ��T_�������4A&�@�K��`�6� }����.Z��T\�l�]���Uc�&Q3>�.����3n����I��m��� t)���o�@��2H� �Û}� �o&���F�WH���n�����!�~��E�Q�v�6G̮XW�xE�Qԑ��_����&���Y�RO��>�����w�s���)i��@2���Z��Gd
�gT`Z�y�O_��H4�-M�	� *��2��oG�I-�+^I�+�x��r���i���{**�*b��c�V���Ѽ �Q=���.��I58L���9��-�\�o۱o,.���Tc;S�ҵ�6�TS �$�� Lӽ�P�����o�Y»���ik�
��y��KA�r%ҹ�0��->/�v���k����9Vf�/T��xU����5�I�Z�Ǧ�/�n[���To�%�K�:���D��));��a���3�<��7�	{q���Ng�]�ޯr)�Ӷ	�ȇ\�B����lS&jɤW���N�3�r^��Q���a�E��A��Z,_��L�����Y]���3�>�!jX�[D�0���b��9D��m2)�T�8H����sS�u�J����,������:��	���K6Uz
)����Ч��*��v��\PX�f��HJy��C#	�	�򘾅P홾~Xk�vgP����g>���ʳ�hV��C/�.ư�b�-�|�»�j>=����,���J��x[h��@�d�Pѐ?XY���H���Us�w(E�a�n9��	��.βY��H���1��2�a��-�A���;�	giIo��{|���i���
bV��!�6=�O����(Y��?��A�_3�mϫ�iǎ�<���A<W��4{(����xXA�:��NE,��s�]@���J�9p�hh�l�ߔ�r��_�@�f��A�Ӷ&2hd�$���Q���^���°_�᝜��3���׍�}(�������VR)�AS��v���9�=[N�6�^Iղ>t8'�?vl�7�BPC�m�'�S���d�t>w�ϒ�C>m~��~��Dʩ���; dC�������v$���X��Y����󿜲L_8�Ht]�w��\��=Hy��/L]K�^�C��س�3	v�5��W��³Wa���mOh�h>��	�Q�Y�c=�J�2���]�T �Tc��k���v��YՒ��D�WDU���3��i
�3f�-����ᝑc����A�=:���F�n�
������������8 ��^]�Ƭ�7#p3E���l0�^-H�`�
4W��4�����v��+{5Z��^�y���z�)����#$fF�&z˴�Z�jPBs�J�afE��ee�F��b��G;N��o�N\2��>���&g�\^���7;��#rG�h�� %�9�̣Ko��Պ��J��Q|V��7��l -6ZNե���o�įt��$-��y��F&q��U�,���+[Z�1o��(������S��Pz���5�<N��]	��&�q�9�⯌�l6����#|A|#�'��^���÷��?c=��"������|nE���h$���㾦^���'e�_�?lR�%F��E�0�P�N�c�_���. v�N5���]��5�☡{I�,G�.x�����0˩���RY�57��U+�m�]��{��\s@3����|-��F�v��1�1�O�v�d��h"��A	�&]����t:Y�y���ޓ�(�Ź����֗��6�xX3��F-A?k�1̾���<K��� N3ר5j|w��SM"�Uf�m��,���C�t�%Ƽ,1�^���qA�>��9�9!�jo��v6�mn����˵Ғ[[p���-�Gr�_Đ�-t��Y�>f��v�»7����E�"�ʖ����qF�<�<���m������ɜ�E
k��Dd��X�;��<+n�l�Ό�(φ�V��3e"C��G���&�����Vd��ނ���=��4�6Ϫ(�CH���;)�E�/���&
����L�Y`�)!���H`nX���(�ۻ�f����x���� ��W����FťJ��Sv����Z��,n�RI�60)?�dO�EDE,{�Sw�m���7�~�����9�K�e�#v$#h9Tq��W�����x޾��>蛑���3W�j�-��_5�$`��v��9��zA&t�'jg�j6�����@k��	��M���Q$[5�
��P�]: �Ӿbܝ=�{s��$_(��؉���x�Z����7B�>ۧW}��b�*�����b|-��ہy��j#d�R'��4%f��J�1+;d4�֢_�mm&4��q�� ���f�v'�c�M߽��-��:A�%3�0��֠AG~�ؤ��������R-�����H#Z�M�1�^Z�*Ex��U��V�ϝ��U�P���?� ����0>�:�My�[J4Ŝ�<�"�<�Įgx��'"y�_-&��Q�G�n���\Q[��5S�x�Q��67�^� x����BD.d5�h���5�����g�
�ПeU��ʬD���^�{�ß8#�����{y�U$l�`�"#�߸�)'P-:��B�nph6�L�yy���y|���%Q%��U�:�?�D�z�(��R��A��:��$��u��4xԎ/)$�ӿ'<� wYb��z�� �@�?�0�\�����ig5v�X�X�%PG��i����$��^{w[N=����ƣ�)i����i:Dw��T�Y6���I���èf�fF�e���h��\����#�#���ԝa-�;�ɳt����I��0��Jyl[!��/�)I#S�m;[H��n<��YFtⷆ�Ȋ�#���i3�}Y�1&�����f�����2���:09˲~		t�!s�ͳ�AM5�:x�U�ή�g��<s�%��dQ����y�F�WB�5�y@�z�#�xsFO}��O3m��&�����b�F��ө:�� y@�T��L�y�w�sU��'�ޛ���pE��?�g��U4*݉��3=���i�n�>�\ک�.��B��^�UW�~��	g���N�Gg���L�OfZa4�/R���F�<�7D��:o��߰R�*��l�bXq?��{X��9(����	��zƎN\�K���a��G�����'�9fT�N`ҡ97{2����w-a����|S'ۂ�~70!��YL���W��n�Ϳ��v=�h���}Ʒܗ9KWIEEϏ}�燒�i0�t�
/�gSX�
.O��B�Mٌ����.�M �T˽v�:�����Y:����-��F�x�I{��r|·R���=��Q t�t����̎p�jL�4��!K���.��$��>/&V�t��AN"Dz���$�U��qg�n�Cw�]�Ag�B���Hh��x��&Q�]�2R���C<�W�RR�CA!W�N/��)�"6U����Q�=�3�� ��P�
�72��ǥ*���by/Z��o��JD���g||�PM>��a䖛;D�1�����k,��C1��Ä��v�"#1y/rω���E�?�x��Ѩ�L=�����K��8npbs�o�L�p�`ȕ���?6gjjVo�=q{��Z2�Q�$��P��-VU%�v�4^����p�K���U����3R�S�r��P��N�؟#D���UmY����ͬ7���XA��miI"Y&�'jgA�eWYi�g��1(sk扥
\�iC�E�y�����^x�ON�X�WlӺ���BV�3rk�o�5����=(�_!�	>s���"��&y��/s7]sw���6߂�9�fuPk�AA��C�v��)]��uAĆ�b=���L(�qFnh��w��?��.���E)Jm�r�
=*n������æ"���v���M��&M�^��Q���9ۭ!��tOݖv���!�'��wȓ�V|� ��
�So�1:�D+���_~$�ѹ�zJP�GV�FfL�&"�q����+�+1���o�W��JI3��8\o*��}�Tb�(��H���x���Kg ���M0��h��uƦS���8��V��spn�(��s�d�0���v�Rrz���]����׊4�#-m5�(�"i��_�q^�����h�F<ڠ��e�\r�SE��
��k:قQS�j9��gp^
.ٚ��F��5A���.s��;�\�ݏ�S]DB�ă�x�-�U��HT����_���&Z%��C�ў���w�ro[[Z<5f���\ZW�#%�L���+���h�Hm�e	���� �Ң�V�3Z�^�&@69-%��Yʹc�֦��B3�Hm5���xճ�@˪�Z��w_!C4�=�]�/�% �"����Td�f��H1�l���E�5��d�R��u��4q�-�t���+�ݦ �Ѱ��b�{?�}O�R8�����ԫҏT�c����[=v���dW��'I��l�ƞ�{�-p�~�<l*Єc�E�}C�o��ah���Lt���s�]��ӹ�����E����ҳ��X6g�iS��;\�H ��ǳgstl�����D��]B;&����P��G�Q�5��!���z}��h!�:-:��K_�(��+�׎��9�3���Q�YQ��P'�#^��E���c���LY����e����$�b�@�}�l����[u��w�-V�:����4n. 9�����WDIA5F�L�ox\Q�|<�k�k��vKyI�� �,�9�/�Z?�Zs=���ӄog�G���'c�Z�,�	D����(�?�W����CŞ�ѡͲ5�g���io�"���z�r��<a���'���̈́Y�4˩dU��*�u(�PE r`K( ���Ǧv�`�ݦ�g�m���)ߎ�Y!	(�s���]�˪�#�_ƒ9�^,pz+~$HG���_�x���\s���$����1�@��Q���yS|�{b�ݘ��7z��M`�������h�^��,�T���%����9(�[Ye�� 3�6�m�v&
/����$�����XR���ヂ�I�h�������}��=&��ƣa(�X�	Յ���z]��;��.��l~}�T�9@8��Y�k�a2`��2���uz\g��.vM���;2@��aQ�	�IHiHp��Q�(v�	���_��3]�K0%�x��:E�T�R�m��Luo���b�e��d�~��P��a��� �wB�� ձu��皸�̘�v#�7�h��_�G��wk��D���Z"[�r���eH���*Y�A��`��\O�Ow�q�	�p4���2Q�hD��E��>�WӴn-k�DF��Hn�hSPWj-7�@Y�_7�g�O�H��ϠQn��D-�L~����S��g�Uh��6i��g�� �Q�� ``;s���rE�,~�K���?s6�}gl��"Y�3b�Ng�����#g�R�.]�+o|�����,�2�(��?2��Ս?O��ʚl����(�K�P[�90��Z����'3&sޛ�|3Ԩ9"�3o�~����+�!��P�`y'�Y\3<����wθݻ	�D�;`�to��z?��Gp��!5aI��|�_���A/{��'�<��l��]y8���XA�h�6�7�K�b3pՐ�IOSb�\�蕆M\`��b�ԧU=���%ݦ���ñlv�G���Cb�����c��N~\����A<t�������]
��ى��z����_ҭõ8���K,��~�c(�.�ñ#Qԙ�y��<�J\���Q}��IFV�vI�&o�a��%M��R��s=��{&�V��ە7�z�(���2lY��b%G%.��a�Y=U�Q>n>M�-�y�~�K��������V��%�|d��eH9>p^�9�2�W��Ws�Vw��y��,���s�S��!�����gi2��|��W�e��䟖!��y�������J~r�\&���Z���t��-f}#� ����_�s�P|��X r�U� %^5�k��]��I�P�0:�����B���C	����
�_Խ$@n�-Օx\��aq�����/W|Ԋ\���	lp'el�7�K�_���02b�rrf��l�
�A<�̐�W4������7�����r}���7&��C�k,�����"���+��S�xg}c&M��;Yn�?���2���NY�_��t��% ��?�����Ӝ�nq$�4�=v�F^�o��R�~G�<O]��5�N|"�GT��<�άI>�� E�%�����ـ����ݒ겄�H�z`�S+�����O��@�zo�0���0��y���_@�+n��Ę!V9�i�_/���j���= ^�m�������Zt�`v�G'�(A�X(,�s�N%���]�кbc�/�R<z[��P���~^G����_2B�p쀦�|��~���wyYJDs�S/�f����	�E|��&2�GU(v�ֶ�������`��H�QPV	����9 ��T����%��g)���J��C�H�n��p`��Ů蟣��܇�(T��0�̠�VB:������܋�H�l{���RZ�N�`ђ�	��WC	t���
��ʁ8��m�_��g)�;c��f)T��
���q3�ע�i^��,n� �-EC�4s�f//�;�Zi����� e���!���#_������V}=lT3>\h�����UB��D�[�z��2I��z� �/S��e%������jl�r�U��1�^��D\=)��9�܀�#���_�-��n��xb5W[)Rr�|���߮J����#
<h�H��P�ۃ�͜]I�����ƛ�7�x&���B;�vK�����*�ɭ��/�8�7f!#��5���\_�_��J��j�9j�}�fW�~�I^q�(��1�s�k�>�h�ˮ��ȬU�e��`�q���wֽ��P�n`�\�F�i���5J5ᙂ��{�$�z�f_,��O�p@#{��gJlS��t�AsCxo�l�Y]���c-�0�|ёd�9�]:m��oCfa���+KҬ�^3Y��Y�=��W�(xF��,�7�Ͳ�$Ŭm8F����#HlWK��AMy�����G^�������@���?�؈�W�O�X����5#�>���~p�@�N��nĚ�%aԥ9��L��a�
�Nb�����YH�G��-@�������U�`�$�����PB5d���o,k�
g� ��W�����U���3����ѥ0�9y�,_P�~'c�� ���2��'�d��pE ��g�z2����&�*r	@�C�ۚ ��1���f�s����,t�F7?���i����vfq�I���o�b��j����V�3�o�fөN���	�z�%��W�jUvvN�Z�Sp��ZG����Xy�m���r�X������T��S�A^�Ʋ��
���]HJ-&N�H����e��ɥV�a�K_�'R���k[ ��������՜�~��Q3�2g@>Y�ΰ�	�&� �倕V[P�Ԯ�,�{)O&���?f>\���4'6�N�(�����񼔺)�x�i��!����ys6��N���TԜ>L�A̵K&(�W	59��W$`c�1����E��O�����l$E����3�k�P�R��1`K�O�o�%��F�"Y�W��f+�����CmΙ(��^Ɓ^/���÷4�K:�т��g���#�*3IN��+�Ê ���9~*�HV��[�Dh�qf2E��}�!����y�/x6^ȹ�Ҍ`����;�W�A��Ӡ"� �8��^@��v:�s��R���]����?]̄�:yjr�'/@bJ���:�37�,��	� I�[+��k��>s0�8l�R7�s�;\=l��C�������$�9�}��1Op������)1~+A��]J�tR6F�˺�!H�� D��j�g���&���7�~qGa��"�$����3ˮ����Trj#�VG��jw Ĺ�����4�WV����Jav�e�P���_=Ul���y[Y�tuu�� �����f��V�d�=/D\���������PN���!����C' Yu��S�Ύ�Qv�2��eڣ���s\��G���h;6�O�<�'V=3em��0�����*����`h_�{�E�.jq���IY�cTUJ��-٪Z�bɛ0�r�+<��i��������N p=�uIU-�5��!�$��eR#��J�����~o �61���}��gg�M�kz���2Ҏ?����>"�#�L�h(�Y �g��p�7ڔ:�[��0֕�p,�/�M�i��Ɗ-OT�����ʁ������ڷkrO]PK1�ܕ+P���������TP{*�Z�JtP>7,^?w��b�9z�H}�c�;���Ӻz�R��7JI�2ϥ��&ъ��0B��`7�5~b�p*Y�2�`������N2;�9/Zǒ�^�9Y��m9 ^��#C9�1����j�	��1�_��:K��F�]���T���erR�����>����KO?BD.��^I%	jU S|�xKѰ)�m���,�jz�����%G�f�]$W�V{�����3C�����]8z�s#]CZ|MLIal�7i�.��L�]x��p����Ή��F5������O{ɿ�ě�,�_�b]�K+�[�����8��|��AIyӋ��o�����I��͛\�1`����|j0"��iwWh+��Lm]��C�:�Poc�^Z����7H����h�A��,�V5kcQ�f��?w5����:(Lo~1Ӛdx���o��F�9��8>�]U��UB �����0=$�ww�{2�)��XL�K�0��p�3���#�)R���%5��\���>Ŏ�èWu��Ui&r~ea0�=�K�OM�O/�5t��'��O��m��Rj���]���yҶfN�Y3sw�4����Ԋ�=g�~�K�te��b~����U�\Q\��ZX@�C#���>�M}��^�>�2���C+�w��{bŖoSȨLi�alE�+�8Q�j�I6˻k��㿙T�e[�j�up��x�N�{
t|;�BP��+�Q5c�1}r�o-���a�rҶX{�64ra� mg���l->K�9�Ȩy?�VD�b�z vS�A��ЇR���E�i���}_�d��!�?V��&j���q��P�.xڈ��EE�p�	�x*��+-bSE�J�����u�d�*C��F�� ��:���,����D5���H��>��O�ͳh�c��T���������Py��v�$K9Pa�|%�q���pVb��4���-'Xm���BF=�*��m�[�����s(ԗ�֒�o�K�/\O�iS�2j�{�>j��uu#<P�[���!�9�u̂�َU,�Jx!� �MR������:�)�uの����Zk�`
�n��F_Э�P��D�(����
Z�x�a���G������l�����E� yJ��m#ɔ�C[Tv�*;���I�T\��}X���5����o-����h��W��AY�	�"���b~��dP	.���p��Y.���452t0	h;�H���N��(�|!M����ӕ�y���\���>�ZP,s��{iU#mI4�L�H�+�@�),�IS#�o� C�Z�Hc��(�-2�W� <u�"�܅G5[ѻx�:@'�h�xja�ʜU�/8C�\��u���A=��91`��{�aʪ�3���Pu�Ɋ��v���]�iϭ��oTh)s�0_��i$b����$@v�o�盹̋��Wy�XG����n����"T-��=�ÆE�5`�J a���O��[�DSt}�tvľ�B����AI���q�^��~f�m��
ҥ��;�׹m�<�أ��}�X�rY��3�.�W���)�Q ���-jP5�`��|��Vd�h��L=�� �J#V��i>�3�V��XT�ᅹóx�a6y�9~���_ɝ�Ɋa]�>S&F�=���^ұִ���]��܁û=k��<���($Sۉ5�-�����P�I�v��v����Q��Y11�CM���CnlI��=w�Ym���)�~�eP�
[r�AE��׸�\Za��1��.C�~Es)
��;!�̑ո�z��}���٘}VfB$����()["������]�.�s@J&Q#�@	ZK��,�������R,�-t��}6b.�A�f�;tL̛�]�{�Vzx����b�Sx�_b
F�"#&��ǼW���f~��TO�FM}wg��b���+a̹T	���܍�vpX��h�~b6!
�� ����W'�[�����3�q֯�K={�]�d�E����(����
�s�4B*gNG�VTE�	^����&��`��氯̠��,4��h�_:-��"�n����Yd�5�l\d�|k=����+���C�O���&/�T�&�~�*��)w����n��$Z��!'��S�.����GNG�*h�Z�o�D7���V,��v8D�)X#V�=B���A���\sNu�2��WO���H��0��A[ei��-�N��q�̫6����Z*�:�� �@Amc�M��q1�p����}=�����W�i����B��k�u����������\��:��S��3b�&A��!6w�i�_O4���'��*���#P!�.����QC��X�J ��02�Ň�`���o��_'G�b��a�q���0_K\3�KZ+�6�"���=�T�c6��������j�����;#ĺu���G�Gc������VRx�������Ik8Y�(7�]�ΆG��?�Z������ts�}bP��&����?�_|��+�LQ��]:w`Z7�>V�6nQ`��*1�-$)^�@AJM@M;���*�(�h(�d��1��U�#��1�0X�w��EKchn�׌F*�K��D��#��w1RŪ�=��D����B�t����_!��-/C�S�'֚a�S��[6�K��5��zY�'\>���n2�C��w��[��-'�!a&���p؀������h1���&�>h�H0l.��&#�����> 8�;l���ME*�7	hhm�������[A�/�1LpH�&{��4�R��./9�M�{�9�F��hY�܃���	I�lE>���	�ھ:��V�aQ�`��V��%��v�F�3��P�pdw��5�]��H{XV����"��d;%bݞ!���M=܉K�'TQ�a��*t6�ՓTH�PwMmo����	0J�x�T��I���������jX�E� ���#���:'�?���r�w1ey.93��@������e��.����uz]J!�d��u�(�U"�̉��L�u���p���ň�sY����]��!�����̗S
�O�v`���i�3�����		it�٘m6�ϧ$U8`��"������/Y���
��$O�,��#dT_B�F\�w��*m��ھ�-aN����w�k0|$W��˚eZ�A�<�Q�3�Ѓ�3���}����9��͈虅�dN�葮�1��鍕����c*{�����k�P�S(=x-�d��O��FCE3do�<���J5e� ���3��w�Gs���N/��^+M��}��Y��n��_4+�S����F�" V����J�b͓%���)��i�£�"H��wUq�/�ʤ�L���}ə�Ѝ����,Hg�z�S���f�_z��LZ���ۯD��"�{��ȫz?��\����u���T���12S"PP���w�^	�;7��b���~P�m�ܩF�$3�(�	v2�Io���g��=	u�0Ym��%d���@s�b��
����jl��Siz��$��p�!>��ϏVn+feӠ���X�l��}?^_�۱kA����z��' ��P!�/����>��k�A0	�bU�F�0���0��-0ģ�C��!(^g�T����˭Ǫh$sК����d)��I}X�/��4"$��M�=}����z�)�B��rs�e���L��AQErĔ=��KW��y���_�nL�A��k�T�����).�/%��ݘ���\^V�i���exq��{��`Ir<�bڑ~������%�������k;ɏI�bMT���㑻�����߹��Z˨��:�'B�o��!�*G��C�������M��Z��"%|Q����)����dc x��+�*��ɘ-#Z?z�b�y�K�l�����Q"Y��Q��u��3d1<�D3\W�B}��q;P� \����ų9KH�G#��X�ׯB���\�P�@��UPCH@cM�ο�]��u�RJ��]��r;�IX��4l�܃�.��������X�=v�Ao'g�r����O��e\�ɑX#B��_���3aw�����'�U�]w�q<:w�.kqLT9��މ+������ŧ����jO��n�#�Dc�?�%7r�?[�R����$?(���5Lde:�I�����&ڿ��̻т���@ {)߉�7�W�<��&�Ǻ�̼�He@Dk����b��������A�������A���AB*�eV}j9��+��S���&���	�s����	�]r[�- � �9�`Y����̘�����̑?���Q��]���I|�y���ɵ�	XJR�A*O����V�$�No�X ^�$	9�XNhx?#�~��R��{7�V��F�"��nGM�'
:�&
!���x�ȋ��i�^�S�Z�9���n�ؒ���ڢ\!�B�'=�%)4:�,������?Q�m�W��[�G�A� c�Di��L�����~n����._�xv;1��b6ftm�(�w:��,e����V+a(;����&�Ay9.%yl����. nv��Y����f�96R���i����[�  nču��`��X4���dc��kܫ��X5넢��l5jn-�~�,`3m�t��ł���7~����n�)��b�{��*$��y������5��9t<-�d@'��X,��Us�|Z��̔�Śx�.������01_����KϜ>[��χ8v�^A�P��򐖖3�@�6]�uɕ�	����[�}�w���IfpwD_L�8�m�7�6��l�U%�G�ʽ\�!\���߶z4�kG=��Pm�s��=���M�*#�����QY��|��v�L!�hW
�n�0����)�0�R!�7p-�^]3� ��z��]>:�Cd�M�,�byF��.wb�������N0��-��	�)��Jz~���Sn�� M }��u����ufA�k��S\[�\��7R��I:(#B��ɛ�# �-�U@C����--��ZhJ�G��k�%�.YS��B�m��H	e;#�I��ݥ?t�S�d��봴�5���L��-��g��Z��J$%�R�/=�k7�H��٠��}�н�ODӈ퓜�C��0^����ث��di�g6W��y��R>�<��1��r�V�/�l�C���uq�~��G�$T�9M�:�:�fz�ޓ�� �Co���ꊕ�b2��)��3� W
�J �����V܃�u�^`"�L�8�8��0���%���7�9V.>�]����쟼�j��פ#{Ue��Y�V	=L��s����=�^�4�1A_�H�89�� �g�TדjCe{y��q ? �٠�@y#Q�6�I�3���Y��X'�$Y�|�\�}�$��A8h��}��G�/�=�bK?�Z�	?(�'���ơp��z�<X��U6���?�w;otC̎� ��*��k�`7	� �+:(L0a/;x,�(&���UӀƧ��p�u�.^¨n���ASv�e��߼h��y�d��y���J���F����+;��[{�Zju�~�������zx���8�g�s�;Vˏ�C�/D���ϟ�x^^��lv�������m��;�z[R�����r�!�>�wI�(<�q ���Kg���F��S�j+7���&j��h��S�D>���o�X�+��;�b#�\�2�/�|�=�mH�7nF�gD?�b^��U��׌���u����7ش�6e/p��&�3�ן��*Gq��
�%ۃ��*y���~E[��8�+ ��UG&Q3-��"v��Y7zrZg	I{�vǁ�g��F�AxE�ha��v�b�$1G�����ъ}F��s��6��KT���
@(�P��%��'�06��!���s���4	�?��Sp����d�j:vO�VQ�����ވ���*Mz��I`�Ϻ���lN�#��F6���UcRq=領x��gL�&�����t���+� ���ǩ��,�p��"i�����y����
�qF��4G�2��;y�Ё�?{���eޣ����:Ք�ZZ!��[nw��j�|�$ym�9�	Q�ǃ;����٧�5㺾[����hJ��b��W��6G�@��~rl�S)��h�!��eS��8���ϯ�M+������I�����T����A�\�����tL��Z�}tO4/�乐1l�u��	���oS��9 ���u#
�J�R�&ʎyY�K��[c�74p-Y�U e�r:�a�K�J����F�v&Xm��/�ـ��]>U�zFu>ƹ�
�713�����x$���:Ll`����9/ܦ���;՟��`������I2�5��n ɖ��ya�	��/gxg|g 	���u:�{�%Y�8\J&�y�a���e���ݢ�.(��y���:�m�h�:���+J�M�4V�|@!���l).T��O�K�~%(�5HKs�@[�n���N}(�9C�0�˿����C뚫7�����٭��e��^_�|�
�]ʠ�ۆ�����;����p.�֦H�׹!k)�aN.5>�� �������EjJ7�SIn�Վ����_����P���@�z�d�?^k�O���m�y������6�<7	5�e���dh�k�ԉ�/�j�FJ���^4rHR�Ѿ���ڬ0����L�>�b�GEbʿV~�R�O��r0p7T�5�����g�YB��ȫu�� �6�➇�N�İ��UT�V瘻����"Q�}0[e?#�I��v���)%ѫ��i����\.	���B;���*;���<���!ۘ��nk���s���1�o��'�7~+:Ė[֭��2���[��0�Fd5��`����&V 9��D���*T�p������MɎ�=��$X�F��e������ߩ"5�����,�Ϲ�	���k?�]dш����b��Y(� ��������Zͱ"��@����;����`�|̝}]�g�%qY�����zzŭ:�S��)"�*����2F<�0���^�`�T~����R!������l��W��IZ�́\��
Վ�ra� �ɠY0R��\������l!���L)���aI	Fb��y��u�W����/��p�Zms��ſ���S�f�e�9���n��Qx�z\g��<��7�ǀԹy�������͜�_����d�^�Հ� q䠤���KCC�Q�&����p�2#i.�3�s�R�n�բ���c�~���"4;�*	�d��ݒ�6B6񐦥���#�3���4 �"�k���g�Ȯ�։��0��nǋ�0���h�Ӿ{����]J_��K~m'��H��zI���p%ɪ�=���7nN��`��c�Lk�������2�b�iċ����f��P�z��6�ns��.,���mV%��s�G9��'�L!�R���@�S�{/U��7?n��s�X�ț3�m��{�	)�{tG�`<I迡c�r+��G��z8�{�ʊЁ#9k��k���=L�3�&�K=o\�U���3[����.8P]���(��r!Zb�vI4Tl�ē�W�?�\��
�3~�V��K���+�e<��!:T��MA�U,v�j��D����|`H������IvMu#�h���ꈦ��}�1�JI'|�	G�?<�r��=��e�Z+y��B�`�2�K_�p���kYP���4Lm  qE�����	��sg�����b\т���X���[Yv���5�C.p��#���n���3�Q9�&�|o�����\��s��O���;�X�#dv47�G�~\��q,v��<`C��s�lkpqY��1i?��l~���b�)[Dz�j��u�� ��C��wt-�i�C�:�o�.G����X����f�D�L�W_�;j�l�#��������Ȯ��4�z���أbf�Q�V���
��q��/�l���D�w��>dngL�+h}BQ��a$��Iܓ��x�y�` v�LmZ��/�k[O� ���[&т�f9���FN$SS�#�Q�+�O��uI����w���6�w�l$9������O.����bv1�;<�a���v��6����{�H�MRp�m3���
�70�z�DES�!���^�`� �ٲ�g܀ͧ>�2(b�C%��uSKz��g�����O\CP������K����{��Kn��:z�����K�g�0J��W�]C(ֱ&�/A��d�OS�~�씂�e����:=�4�r�Jgdl��de�l�f���|��̇�A��Z�S�A2�7[:�w���!�ơ]yLh/���j���b-�i�cg@͚C})����CW��0,h�!���%��^�uxX<��@��L{0��.�>�U����Gť�;��Iaj;A����9����eʄ���~�`�����Q,o���%��I78�N(P�)�A�G=ʪ���V^>,D��!�F����)M�qQ#%�տռS�C�9���D�7B���wsA1��n�T�?���}��uNS �L�y��,J�0un�1�֟�XY�Ҕ�uP��]�/))[I	�+�g�B�Ǚ<$��f���-X��&0�N�q�J#�q!��P�����_&��ƧH�y��O��S��jǽ�hԀ�3lf8i��w�������t&n��h�B�����k�2�{&Ɇ��|�m�б�|�Ӄ���Z&b>�����'r��fX��%5�^�r(.���|rk�Qeƙ�3>_�+�%��mF�"��.��s�1@sv� �_4#9�Z�	�}�G��r�I�:�`��D�V������^:���^2_1�+��ôF�2�G��D
��G-p;�����ui��@�3R���ҽ:�kwX��WZ��* ���;PjY`��,��j9(N�}Y��R���h�C�R��#��A ��S/���49B��Yc���U갞�v���qo����t�J�ߵLY�j
<��������"��d�v|5Q6���!�dZA��H���٣U����"7������FGh�>d-��j
��u��H#;��U��uDG���Ilǖ��p�J��.�6
f��;���{F�����*���no}69=o��i�~V�t������.�w�ì�~ŋ��OyM�����>��k��/*{�}?�2'�D�B]jQ�b`?I���yB�n%��ثb�QF�5��3��Uj��V@�S�F|�s��F�>>z