��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6O���b�;�_u���戠��Ŕ,�8O�-�7�"�������Ya���V�FZA6��%8&\�������A�)/-|GG�1>7Ň��bA�yB??�;?u�gd� ���vJ.qL=�۫WI��~s�E-1��2J���X��sT�<4���g�P-�W�� ���T#N��[���8���
����=/ �B�d� �.e����-�|�i�Mp�]s�we�L'��P$��t�u-���v������e�)�:�f���n��ϵiΤoY�"Uka9��������������V�%��FtƳ��a�5�����
看��~:'�j>�>�v�]|�n6��s�M�L�!��&�5=�Mx��29H���z��k��ASY|""4���~C����}�h:��D�W����fk֩�/���X6�n
����4���?�-��
Pg�l�i��wZ�����  J��5Y2|1�P$)țf��d�Hj*���zT�:��ҟ��n&�oF�� ivR����D�����Z�������a"z����x��$���N�nT�A�}�g���:''�)���x46%�񢯳���X(O�EX:�����gE��.g�`���ـ0QR-���N[���s��#;	��R���ٌ��>��������1�Qg�p��pp�;G]��w����}�
��v	/�By�h���_<���ٓ�i)\�ѕ����d���sc�e�%�2�c3b`��Y�����eu�BcN�����h+���솓G���384&�G�A���%ю��:f2K˼4֑,�8|���D�wW;��p�)&���B{�Ϣ .��'���K���+�tfS�Ut���PU9�`�����@�'�����&�i���w�ک����E5��>{镃ɀ��:n��f

��?����hnn��l���i'��z�bk�
j+�+�`R%���q��Ũ�]GK�r��Qk6�`� ��n������	xI���S&���������Nd�c���u9��0�w�� �1>�Zk���%�Н{tL��<��U��z�X��Wd�H��^�>���G:�]��)��G��a�@�U�]$��*ta�(�$�+�LxN�./,X��:�E��O�����T��Yi��U��Ps�c�T��2K�O�vf��U�N)����L�9Ll��k�O1�?o3b������s��Ҭ�9?��.`���-J ��v��yi�~��E��(�|=<����Wb����C�o-�6	nu��7c�ㆋ:>04GOv�|���d^vՎ�3O��,+�4�7�9:W��/^P�aIޏ��=S�	�* �B�LH/β(a������:p�f
�կO�u�F�7���E���qL�,fp�����S"/�[Ɨ�SU��g�ƓG=�66�@(4
�s<���F�Z��9�_��]'o��u..	NWos�!W�e�t�Ε�I�l��a���h�_B������E"�X.�(�ݐ>�z�[</얱���1
S�k�G�����GFFM�W��S$�����u��;ح��\�G����SzN�z���_�ģ�C�Y��xE;p��<q^���A?�<��W���k���cV�V5x�3L��ݽ��:���ǣ��wx1g�W�ç�x��^��e}��"T�AZS���R�ë�J9p.��|MҀ��4�y<����Z��ktp���dx/��Lh�S�o�S�V|ٳ'$`/fp�md���ϒ*_C���l�\ `X��a�Ӂ��h/������KȜ
eR�hY ~6"�i1&E5�PR�ډf?�m�53RGfa�",����k���ǋSi�-h�/����5�C	�Z?�Cm9Ӟ?���t��Q,	���۶*�31���L��YYl2���Y���d<�}�����I��Ab`�0�ZzO�p�g���H��xE���_��QG0��w@)L@����T�n��H/C��"���f�!���{j@�t�j婢����fgx�ʑ�(�_ܚ����%͝7���Q���!�1��uz�L��A�^!)�Q��Z@��D���e���PK�iL�ފ�Г���sw&}�2�C��Rm�����ҐA�xޤ W3��=��%l���O�H�W��[r��Q��v�/�-��7�D��h�ۚD�QLD�����z�&%�b>�(|n�⭐ʳY�7膍�N�@�D
���9��)�۵��Yؔ�§��s(�o�x��Le�-��L���
Kݩ�)�|ʅ���8��o�v�� ��Q6$����t��.�y@���n�!�V�닶^�+5Y�d���g-���/�{<�l�j��$c�6o?�k���/�JOh�D�Z_B/�Kl��'Vj4L驡pM3��ɜm(���S^ǌ�C��3`�	!�K���4
�mk�L��nh�k������,N��J���M`�jd^��x��K\�㽥�z�;�q&�L�hg��
%L�*=Lܲ���~�/���>-e�e�!�/�����e ���<���/�6I�W3;����"��r{���F<��(j��~�37Y�/R�y#s�K�4�W�&2č�k[�� ������ʭ������
��mUIO�	��N��f).M�f��Gì��!�4�`G��or~�Q�t�i��)䩴�,�q�0��/�2%�X���_A�
m��/���F�|�ղO������y��i�}�0�o���TV *R��ao��ӣ���y0@4�A��KbF�,�AD Njh���}U�,�@P����^!:�ND]䍘���p�9'�7:�Rk�������B�Bn:p����NR�ndÊ�I��!��|~u��{m8{O�p��m�%_��@�$9��ћߎ�ޞ^�e���҇�R�#u5���LWxr���'N�O_Rq�U�s.�)���#�d��	I�k9���:������+C �so~�Q�%�@�b�EO�\P|A���/��:A@��\���7��8TW^��y��S������#R��d�9�'d"+^�����G�+�P�7NE�2͈WC�am��5$�h�������q�Z�M�|�3
P�}8��oH�j�5Ib�뻸t|l�Ɋ�fT���70��_����|����o�-���sB\*�v�1Z?A�\�|T�3U�ݵS���q9%Ф�~�c���EO��N��[�!P_�{�Nm�������ΏgB��>���b�$d�����CČ���oH�J����iw1���\�q� ����s�9.*���!���n��Xe#Z�[�B; �t�Ipp�=Y��m��c���dK�9	��2�R���Aϗ���(j(ѫs��F4�5/�i�<W�@�I���sA�f�^Z!��&ǚ4���=��������c���2b�2 YĖ��hBd�O��T{��@t����H57�����Yt��ֈ��5K���?�_�a9Y�{A���.�E � �p�ù��������{CL��#���1�Z]joA��i����.���kz�3�K�����D�3���l��⁏�;����%0u��B8w!���y2S@#�x����L*�Q}�f��0�����l���?�y��A�3�����AG$������r��U�r�k�E�� [�(&K�}��2�olgs�ʽ�^FX`#���F��@/�y������?5���F�юWf�ƶ��<��Wv8m�C�~J5��W
��#���G��f��c�'>,�0v���li|�<�X9�O�5������=�_1�C�́la�ق�w�70؝���|`��T��9O)j�Ku
+��=�� >����16��ܷ`u� ^�.�F�I�H�Ms�|�'r��QE(`� Q�!! ���T��:�Ot�;Q!S�
�[ף���F�o�{S:�A�Tfv�*��<z�hN1�B�q,����C�2�&�Gcu	�>YgY�k_h
����ҹ��{�#��aI%ial�4'�k��L�{���qFA	�R\+x�ݙ�l[�]9�+ߴ3uk�>�Iy���
Q)�i̹�L��$5��x]H�ӂO��;v5�|y`�o�u5�rhdM�fVNк�|�vi�q��?&�6��]C������"5YE��Ђ���[� gUo�x�;da��"�l���A�H�5�K�9��6U̠��!������P��U�"�)���gY^�F�%��#VD�7����~	We�'7��Q��1o8{�[�����T��~��x�m8o/ʮfo� �R�0Q\��h���ܥ�ύ��������[�!zsFq�v@�3P4^���E&x��`��qa��qEH"�E5�&�b\^�_U�f2i^����C+�� t���֎_$��1{� �rp����pv�<G�_Z�[p�u���@�?'˾jBv�i�ܾt��Q�.���_�����Yx0�c�u�����,��<?J�^�O�#�q+�	~	��ÿ��T�ǈ�.?�q��)|�����+f�m����;�Ɗ�79��i��]�#[�UײeF�L�]��fx��Y4��0��.;�[�l�t������z^͖���(�Y��Ӧ���w>#,bH(��g;��k2~4�F��HPc�SV� B�yT�z��Z�қ8�3Y��j( ��n^����m�o�(s�p��闭���q��נ��q>4���z�L�����H�����MC�}I�Ss�I��Vhh����*X/�C�k#�Q�Y�dX�ǣc&�� �uOל	��_�)ʥS6����Q�k�U��c`�t��+'Y���� �'��Ϩ�$!\XV�ϗ��
���"���Y���Cl�LNf'0�a'��fI\.��SZB�& ʒ*k�#C�cS1�r��u\z��;��Bs
 �g�ReȚ��噳LA�t�̙�7�s��+�����K+F�0����S��Y�}�x5�dɈ�e��ġ7N�֨��)C��8�~TV~�&����W'�'@�+jUG?&>��7��.\����oQ��Tz)�
��H�:§�4/ŋ��:k�p����/�ح����׳A���R�lŔ�X����{ۇx�-��Ku�1�IEy�G�ȝ�j���釸h��)=[E��+
�TV�
��z�7Q�3��i��O�5�E�Xv1`�c>��Fv"��N�G����@�11 tu�?a��w">["3������{�jD��o�Q�0��ӣ�W��|�����ݲ@�W���z."��d'�D�(����-k|�j�� l��T��N�����o2�̓7�N���U�.�K&��_�=���T���kE�#λ#��Px[}��s���Bd`����hv��Ԯ@C�@���c�6��DJ\:h%�A�����ۂ�n^�n��L]Ɵ����ؽ`���I�����-k�t^z��~Ad|>)����)����
x��*N�����0�Ƞ��?"\��`,�@�a{��%;I�½K`A����ߟ��xUS������m� �#_Z}hi�S}�^��$��Ǐ0�#�T�"r%���i�(�D.ҽ2�4 U2�d���^��̞�`��?�.��|i�����~¬~� LЭ$Z�\+0F� �Y�D1�sj���@�`"~i.��5�3�G#�Ǿ����g�gJ5k�I���Uy������4μϴ���&����.Wh�����
>�4��cU!�����D)�XM�����S6��2�]	�Y�}�sy�N��0J7����XɬD	�*n�s���xX�.�o0b��y8���"V�L~KP�^��B���\�u�Ab$��e�m�L6d-�RJQ�x�x� E�r.�`u۰�Q�~?�_�r���-���������^J�#��0�qA��{Yk?cy������U�^C�y�b��X �dI���=A���K�E�x~�\/�8<���:���A�{�y��RR�h�ޏ4���w��<��h ���i;X�L�3�����.����G�Job1�y���ΰ������nX�4�����>���O�<���5�+����Y�#�B��3'�Ot[Q�I�]eXގFF~�Rl�����zi�ݣ=�-t@����M�`�/�w��\�^B�\�����-h�����Ӝ�W,���q��KUBC�[��6ӧw=�^����`-Ĩ�Ys�d0�!��G��x��:��!<�C�9̻����[��L�������cS�s����swU�L���'R0��}1F�.q�g	��.�Ѝu�JG��-A%���)��I�N!��6��f)���X�U>�d�6��$���	}� /��l��� 7�4cCpЫ�5����#�+�"��Z��������1����^�N<c���O�m���N���=N[90{="�oQˋC華C)�C�������7zY�:k���~2c�"mc� ��pǑ�<Q?B�	Mb���1� E7��z3]Fv~�u¥Sth����GW���<%���\0�2KÕL���(�e�7�9 ?v�
Nϛ!e��W��d�䴠4T���o.i������0�?'v&b%}�L�Ke�Y�G�Y�g 6�� �a�z�I��*���{E�>w]N�w�r��y.1�-+�(��9�e������Y�B8�?^�Z�;[KV�rՈ7�g�ڋ:��n@�`���O�}=����H;�0K�ƶ�f�C��T[M�,{�,I�7c.q�S���f�������6��+���	��`�#�Q^�	3M܇����/l��}}����n������7E�!��x�j$����l_9��zޤ�����cWviQ�K�^��fͰHYf4C"��?���B:}��((� 5�qy����2�����T杄�F6W�$}?��W��lђ>\ѡ\=�������2��:R��n��A�;%[Z��}�D���y��r�8n{<I3�G��*�
�����k�4�%���-АW^��IG��u�3r�^9��T�6(�3��^�Z���$������[ȋ��HsZ	�u]������m���� �i6��'�~�dd��ǈ��^�`6.��b����:k����󠀾�n8��Mŧ79g�v@�Aķ:Q@*ދ��՛�O̓t��gCoW�r�Y��=;��l��p/J1�T��xF��|�[.g���G�a?:+��)7ʢ��nPB�j�0�Qq{Y�GS:BY�!#���q۞QfIﴔ�� t�2����I�#G��#]7�bL�s �wD�:�k0�q��|:X��}>���<uW�B�pB�~��T�rm�t�w��֑�K)nPΥ^>ࠃ��C���	{)��UO���\�'9��`0���R�����_˟U�P>$w�ӂ@P� C#;4����]@tշa��3�l�<��K��?A7��Ol��"�یc���;�̝�W�_�p�&X%LC_�)�e(�!Ce���D�v��V��EەX�M�ϋ3�n�m�G�im�a�}V�IAK�\T��?�y$���4�p~��5t��b���?w���K�W����̮�nX�)Vv���Q�f�_���0�'�a-�v�'���Z%�_�]�[C��W2�ע�굊���|�
~z��[46enS,_��)0j�(w��0u/��o�f�ExƂ˘�"���i��ΏU�dمW�E��h�b>A��c��[�=��G>	N�bS��Z�rFI
�7�׿@IQ�4@���i��\�Ɲ�7��"�r�=����0������v���l�VzuZ^#X�rS�<�.oP	(�p�{~��Dw0%ŧ"�R��*�� ���M�;A�eG�"�X*/��_�KcU{]ij
C-� �v�H�\��7�↓J�p"��,����	����lQ">�,��<�^�͞7}=Bhy�<-���BR"���
׏<�A��>M���ŪmUgXu�G+���rL� "� �>��T<v����H�+v@�Q4M-?���|uu�ϛ�
�OVcUF��.�����lb���8�RK���]*Ll� ��Jp�R���	mH<�j��ue�&�7���j]����6�U�U8��J�����d��h�P7�!�9^���f�� �D������ʆi�v�5�^t�������N3��s��ra��'��g8ٖ,I�b�Hg�3'��U$l�]���E#{�M�j,�l|��R��p�m���L� �����$5���K��~S	�\�A�2�ֺ����4�l��W���ǌ7�g�W�=ݔ W˛:�	N�H�����4���N3o���Z�|r������<&��#&�u�Z� ~�N��n.G&DZ��;*D�:r��hZ?��N�y"�����R����x�)�9���<4[*i��$;�7��8
q
"�y�F!���Q[�A�݁��E��"֒�~�[���{�z5M�Zz<;{�XqWR����ߩ�F�����מy�	8^�
��_��`�y&��s<ix�Mi�����l��Y��BN�����b�
�D�s�;�i$?BR9J̥$qZ�kU�~I�z�=��]N�F9��s�������	�E��f+<��(�8]v�M�
����kUbΰ���}+����Iʎ�ƶ�.�zO�P_�1��fQ)sP'�]�_���d_9�,崃Ԟ�:΍j{�C���p��v�RHU}Lt�H�e���y��h�,��N"�x�J>]�_N�l�4Ԯ����J�����J{B��8>m,��D
��GDu`�(��+�q�c��'X���%b1ǼS�/1g�R��I^ �7�������<��+N��MyL��Ȫ��}嶸v�j��v �i�������%]B�n�@I #�ae��'f�UOb�Eە�Ԧ�Zb��JM�=-H��/��W��Um�E�b)�搅ޫ���D'��0�e۶O�Y��?;0���>�����LP���B+F�寫��F��ZZ@�A������9�÷O9?l��,�]�FO>�e�H�<�g�GX��l��� ���R69�U�K���B�����b:W�zuG,	��H�iKV����Ɋ*/�ƹ»,r:Vƈ�6̰[�� $s5{�(g"=�ױ��
�o���S@I]p�<���p'��$�²D�8v@j��v��c�#�Ϻ�?Ǭ^����c��1n~��P6�&�lӱ��)l~ϵ���˸�O'�$g���d��%H㜞��O�.|o�wZnE�H�k�E�p2�{�"��y��D#XN�6�tx߳��N]�AM ��:��:Q̲`���t�{��S�ۖ*��}{w4�S����+Q���������K�~�����NȳND0G�z`��7���G�/l�a.��Y)�)C{�i��� 3��mf��;Z���A!����t���{y:��a��o����r����g���
)����sʶF������E_�̩���e�<YAP]%�R�dx#�-
nsb�����������Trt���W������b�Y=r�{E��~ZN��ru�Vl��%6�8�3ϰ�bx�]E8�n��u?pwk�F~�oK�*�V:�ɹG�m�K�(�O�q(z\�ђ��<��e����eA3I56Xu@Ifw,�/�� o`��U���WC�3魕;KlŹ���ި�Z��pB������?򫓮iq��~��~<�+t$(7Ȁ�;�=q��R�b��9u&�
>�EaAMF��2��1���>�ϣ{&}ك\���8Wb�BM@��fo�%Z�� �d)��g��xd�#��"w�a��6���ג��,Q���7̠�JA=_1D��J��i ������-̛���h!���5�J/�UM�`D���}	�-)���"%��S4X�B!�u�(�������F13���W\����O�K�0�!;�=c�9��M��特*��M����7z ���;�0�l>��q+�
�L"��u�	A ��SЍ���a�j|ۣ�M'zF��i�i�b��J�d� �ҮY�zԍO�9 k��-��}��b(T�M���l�G|J*V3Yz_&�HŔ��� �܀�+;3le�#�N������k[�xn͛0�Օ�*�0~o���7|A/���0i��.ƉI|�4z
���,��w�9�,��7���x.�{7z�9�4{�e�"'T��#�B��s&�qlv<KASƹa
{��t�$�;Z����������]���08&b_71�y��S,yO��r��Jc��r�em�?)."�xwXK2FMo�i�!������Bl����KA�[@���I�$�ō-��+Rj�b�?20C���>�f�o7w����0�)�fک�i��Q<x/H$�<��{%�c�p		�SY�k��<����C�_�K3�+������θ�L0j�
�5��8���Ӌ �*O̪O$&���]~�����b�ʆ"%y��n�o�1�6x�쉈����ew�k	���$9��Y@�WR;�\_�-��ɠ��w�4���8�:ӹg%���-W�%ּ��?����h�.TV����Q���z6�� gzZ�����dJpE`|O���:-��h�1W,��P�I� ��Nb�v���d����I6�F������+�9�I�C�;St&�"U�m2^�7�¬���_=�zm�Q�g�|��FQ���Q�k@}>��%�SO�w=Z�N
���Ο��6��g��B�a���[~~����\��l`���5�<���L�@�m�J������/s�v���������#��S!īS� ��AOc�|W@�Ǹ>�GŪ��腳H%������Hd��d���潭5	�C����?I,	<[��<hj�Oܥ�S�g�mF�k�[�0i)�|?�Ev�*>�^`��0�l{�����p������l�H֋g���0�1�f5'��\+�ϞzTX1 /���J�����=��>�k� � W]��7�*�qGȂzw�	����`z'5�W5�y]�!�i��ej����y��uH�Ԯ[����m��_Ӌr�C�W=BU�ҷ�cN���[r��b;�ҡ�m��r̢."mE��H�O����v�q�BC��������?�����HQ��k-Vh[��T�o�HA���ܜ-Da���;ç�q�l�a�<�m� ���6"�X+j��v'94��k`f������Ȩ���|٬���K�k
��}��2s ̎7�=���}o5ck	����CO�6����V�	��R��ۣ��#Xag��--�����}��B���6e��B�,���j|Y%�xH�i@iY��d������4u��&+
��C�Ӊ��}�5x����;/a2>��`"6���Z��'����B|�2�9�q�Ⱦ*����U#�Ƒ�!����:.-���
�(�-��or8�HԔ��Je�R�-��5{�M�\6�b'� S�&�I�;��4�.+Qilq
_�����t��'�����8s�gUVu�7�9,e��*uIh�vشlݤ��q��/�6�%��ODuqAbH=�4��a+]u�k'�U��d�D�%hP4��sz_�ea�'��3��\�u�1X�bS�F�ږ�!�����������|�,΃×�/"��L� 䡳zxm�gvQЋ��`�!���#��"��JE0��j�&M�<�ì������.MK@�q6Y�#��|�T`4?K�h5	.���i��D�d���+b��d��`�(BV�m�i�G��@��4��.���]* � Ř�)��n��_�Ir�����X��x�Κ+�U7�A+K�J�&���kĳ����H=2�v�C=��Xs��J��v���t��ɝ���5�7����c��E�7+Dٿ�5]�}�Y�Ě�ȿ�@������c-�-�Xĳ5G�K��ČZ����#���ѷ�y��z�e3��̝sL+m6MI�W�G�5����S�B�"9��Q�~y� ߶���s<����.��-ע��F���|��+�M�m\(}��,,ɜI�*�b�"�v�Q#��ρC����?��Z!�5�K]¾�RS	��0;
����{���ݢg�5�K5�ਖ਼j�_�@�����O���)Ro��ۦ���������N��x)�����!d�L�j��M��'���E��r"
��oLM���a�\x�cy�-*�s߼�� �4L������ۍ����J���_����0p����q�y����}&Y���[�"�i�"�2-u�V��-?��Źk���R��R3�6
�O�:a�� �b��8���_җ���N$��2[�d�o�u�l$�q1%��V����n��M;�Z�Pc�������g�-y�I� ��Ք�Q��ɃM�R�J���I���7x@�mP	e�Y.X3�[��9Ol����8��A��{+�*���y�T�O}���}]����k�u�pNc�k�v�Mbo�0�� �9S�[@ Tg("��
b��]*
���s����{�a�~�	_8Z�TZ��ٹbɁ�jTA�t����4�wl^�4nb��Qu��,w��v�(��\n�l$�Ir�G��V���u��r����|��_�����Qե��a�H��Z��$��%��'[y_���	oe�s��f�A��H�q���J��*�u�(�%�����|�vP1��������|n��"��[;��e���T��/��VP~K8r�$R=�d��y�Ư�c05�I�������/�"��\wW=��)�R��V���z2��]k�V#��ޭJ·&Juݑ�,��Xm@P@'<���G6��E^`T�ڷ����aG���q���G8~�M-2��z��q�Ci� �+�đ�pJVVS�/�83Q�D� X�
�&�&�G*��X���#-��FC��Jy�g�3�Ps�b�oq�iiO-#}��At`��c�i� J���Rx@'�lF[:"��*C�ɰpk8OyȘ#Q�ڲ~?<�VoZb��m{�KN�-#|:�Ҝ�54�0<��Dꖚ&��Ku~�W��~�x4#k�t�u]����i�Cwb��_�G��O��Ӂ��oF"��q�H+�����~mO��,C�#��Xb�x�x&i������n���
c�ԗ�y�9A����6�BH�L�?�3QR�5���k*�]�v���W�q�����W����L���l�����������%�ŭ��3�����s�D�Ӷ�c���F�:r ��d������a���=ʖ^���I���� �	_�Ca�61�`ǆ�W�՞ƙg�����dRޡPm�2N���� ���::!q�u ��l��?a�>,}�n��W�^B:�VQE(��6�rJ�~������2�YA8`\��Z��?�_;^@We��>)���Y��b���P���k�x�y6|h^ˣ�>�Tf��V������~�H���pf�%�ʜC���29�y�AR�0"F��d7/�t(*�eՃb�����q����(��D'�u䄼��i�u��r����+��m�L7�o�BfU߹t Oh$�=6����;h[��*�!���D��6�|�_vE�0N��i�}'� >�_ ���ŋ���ˉY@�]o\��&�/o��Q���}@����-Z����L�Z�T�yɯ�k0�&%���7̨�|wcA�X(b"��o�<o�^\���rD��-�Q�0*5�@�N���}�LJ,�M�:{������y4tbM���]�o!���U)�2�E�d��!����;!�]���Z3��a��|�K�C�|�!�Y�={O�"�����0d8�lE\`4��!Y�	����Fྊ@b$�����b��.U�!�W��W�"�
��'$\������]1V�UI�,�D=(Z_xt�nc�j���˭� a���?Pu΂6��=ѧL(T�t{���\w*]|����Ba�ht��<S����2��������k�#;������n=�-9���ɞ� ]؝�P<e�N��;�6��T|�D�E$lv��`|�ص�'�KHI��JZ7�o�ZO£��W���Ҝ�)/���|����Rr�Ht���*:T���	5[�RtP���VM56���- X%qҕ�܁r�ʓ����Ν�JsG�߼P�m�+߹�v^#��+��z�����Y�,�y�/K��zB����}�n�*�&�%<���K:DH�ߥ5�K
��� �	?H_���g�u����x�����V�1C�s������Q�������`���D�mѯ�U�����.MO��Ekp�w�sx�(t5�a��,���pa�1�⋮r%ʝ<}�Y�u���؉�@��Ɖ���u��9���|�"�́3���u�jC�Or�ߙq��	����z�8*ן���05!/�q�zJ���ƭ\���Ydh!v#-q�;E�<:XZ���a���9�~_O+���.Ozg=�cBk�����>���bI����Tx;B���ՙ������"�p�,��|n����'ش�h���z��-�ݢ�x�
e�i0�7��џ���0ݶ�yj�T���oJ�>�~����HF�5�]�X����::2Xj��3��*H��߅�*��@�>�_��"�B�
a�Tq	�]|0�]9�o�&I�\qX&A�8��I�	Q�	�$?C]�ܫlؗ��/�b��j<A�ސ���-�} �c`m�����@p�ϳgQ��C��O{��(����ĽR{�͛	�b "�Bk��V#�1�̸�+�C}�L�yQ���}@�Ї2x�L������ag�A�����n��|s���D>�{��r体��7��z`?�&�3��ntv8N��m�����so�3ur3:�f�X�zI&)d#}�s|'g����YY���W��DN�Z�V��o}!���m�de� ��(l�3� ���d|n�m�2�����2N>5kYFa����Ӫq$#J�=؈�?t���Z/�9'G�`F��?el ���@ض�r[Iك3�}�g4J��O��S*���T`�=��bd\Hb���$�%[ ǙI�bt�p&�Y�n�������g�r=9�R9hlR�wm����*�ٯD���-o>��S7���p��ڢ�כ/���@�����Tdu�H�V�����+p��dD��X�U��'+�!	�����h� ��,��qF��\�� �Y:Z��9�JBLٶ�r-���0{t����[-�~?��oڢ��a<��e2��N���0Kj^2��M�f'�X��Qt;�[�^�WE�f�X+�� �۷˹��MV��~��t�O��K�Y=}}UA�'If�`�:_�bIהw���Tm/fkϙ˴��q�7�,lG��@�Bk�ը"D�e3���q���I��q(�̕j�6�CQ��lEZ����2b�ZY:V�9��u)�2���H���Q˦ǥāl͚�f4��F�T�	�/9QgK-g� �|ԬP���=��6�^y��xL�d�d�T_o�/cܮ6��j��u7V�c
Rsx �1f�/x�[v3ٕ���Kذ�����$Kyh�t���E��Hcm����"��r ����t$#K<��}�k:��7�ה�l1pӠ������wqkV�����UV�z��� ��9ɟ��6Cジ�
=��� �i,�3
L�=�/S�f��x� C�����#��kM�NT�%S8�?��Y�42e�HJ� �\oc�E���_� ����bO�\)�"�Ew|#z�R����X`��x�!�51�3
_��.���6��Խ�����*��d��AY{��y26�h�� +Ɣ�v�tL\��\]9�HiZ3��+��xZ/��i��Р�|���r.�p$�/�,ӸVդ��& � ����ڞ�qN��*����܃�w�?���ez6��v�#�� ��غxm���t�2�u��7���j���r�d�F����{���*�n{Z9��=@y�l��/%�������܆��Ƽ��{;\A�գ}ڋ����#(_���|`���ڰ��5�l!��WI��PC�j�/Rr�#�<[��m����\��F���˻�T���?�r(��WfHv<�ߍ��1���EK�u��pJ*��PP���h9��2��On�y�{��q���XN<.5�u�aה4e�u�×���-�Sμ:�y���g�26��|���{oљR��xΔT[a����u����[J�=�"���e(~�^C����J���"'VNm���S�,��� 	��5���&��������7&h"
��$�)E�2���Į�xR�v}bx'1�S�!���#�ukG���Q�eUJ_UM\�Q*��z�,b]��0�����?#!�(�Y��y�{$�ݯ�-t�˟W;�����nۨ�B����ٔ)k�ݱ����w>V�=M����)�����ʨ�f/�ծZ;9�k(�A�NxHm���xA��Cl�wB.�է�{ו����l�u�ij��$X�A�NU��i��a�-Aj�#!�yA-�Ϭ=�w����5'b�}u3G�����Gӓ(E1;
Z#D�b$I 8ppW_ �`�M�.���Y*��q���B�c������`�X��æ��Cgʻ]�9a9��X�
+u]��-�~Z���w��;���P��5��/:�����4 �'C�V:t��T9*�K�78��N�Ë���F�b|W�N��f�����u}@z�uҖ��@}�#��e��Mc;-�/G�=,f�˗B�2M���JU���x64U�W����~�m/��3{�9��i���АGv��)��4�M�+٠��X�a��	=�"�V��ei�!M�x�ϟ�e���Ak��5xU�,��.�����2�O-�|H������ư�[�:xԏ��"}��d������qT� h\ǅ9PG({�>�E��UR�<I��(t&Iw_��m}����'i����($?�O�4�N�1�5$�J�"����!��F��j��߁Qw��ډ��C'#L�f?��0�A��b4?����錩���S�g8��t@����ǫ�N�s�r�����mlo�@��lĀ@1J�r��z���V����J�������)�!u;�fc	���o+�3�  ��d�O��+��9��Wr��`���ڟ���}�Kf�eg�;x5���� )@�x�p"�P�[V}�O@�e�D�qw:Z�'�,d�WS<���sw`�Dkv6����� �M���v�S0�i�~e�bA�%�Д�i�7�Ǟ�5Bt��E0�Űv��[ĭ�")]O�����Yh��^�J\;���j&P��0�$h����R\�d��/m�U�$M,p����nx��ki��mTDœ��+�aSD�M�v�X;�3��?�Ƃ�%$F��u/���v��{���U ��	/+�59H����n0�G���.2�9$��[�'["����_�J�c�VO��l�����,מ�F�T�%}v�Uk�b%���x�׳(+�֣ʻ��FO���ěT��S���<3�|G�����8�1&���=xل:��8I�Z�w�i�<Rpʺf#d�Н�i}>X�y�V1&�L�_1�h���p���|��=����g��"�r�<�ؕ/J�)���(/��$J���w|]$b��K�m���:�|�t2��#��ձg/�p|X�X��Nx��l����6���20���H_>j��<�>v�D��a��L��L��W~�I��6|g��c�\T��^pU����D�~��7�Q7��rz����8y���@�S*��>g�:�T뤜��w��'�o+��l<!,��P.F1��^�
���I!0_����a��Na!�Ҥ��H�o�{Ij�W?w��N��O��
F��pH�  �!Z���b��T�:N�
ŀ?�A"��C�Mz݃E����m�w�Wz�.l�^�_�0�J�H�ׄ�<&7\d}��0@%y-��_A wg�ܘv�^��$b\�j�Ͷ#��� �j?�z �ƺ��m{z�����o�+�ї��
�w��id� ��0�Ԝ�Je<�Fmێ^4(���f�*n�`�z�?�@�ǆ���ߨ����p	�N;��YZ��{�YO�����Z,���"D�t��q}�_l���ݦ��|��N J<�V]��Sm��V0"m$'�<�)m���^K�
�Aթ�tv��wHU�����R���w GM���$���?%n
��� JP��S��)>���h9[ۨ�*�}��*ba�N��9�4%�;�jH���>\J���h��%���l�����u���)���!Q�>��1������^���R�E�r�����ڧ�ax<�y^��|�J�KT2 7Ϝ5�{\��)�&�@{��6Zк3|}�i6]�M��R������"��e������}�`�lP!o��f;g�W�<��W���HPLkіDp�
�A2g����{f�ץg��n�GV��71_������Ǖ���/��c���{�+�'�)����g���Z�z��Sb��^�ù6��]��Ah���]�aax�\Ұ�
�#���7Ҥ��'���J�S�4�A5Rs9���/|8	�y ��#N���!`�N��Ee�D�>^�'x{؎1�t��t�*�NO��k��d���e��z׵�Imr��4�m[�qIQu䰓��z��A!�BpO�FI�8����r��}�?u���>`3o`D�&�P�u�E�%����,,&�	Gm�$<���cv��n��sA?��j=>I*H���6���3�̨U��6j�Pi�S�9!��}@���@�fz�P�?yz�[�H�3�:P��bmJ��X����VD�g�Xѩ�����-d�&��Dt��z��0H�lcR?ՔH��j,��Sج^�s?y���L��T^���=�����A~�$�Uw�Z0�߮�5���±�M^�kL��~�����^P��I9�P�f<7����,�y�&�[��Q�S.���:�����
�O��h�/3�ìw]�<�.@]�1�@��*�_��L�5��gwQ8Ѳ�H�rP"�Ԫ�l�:=n�w��v�o+�sf��˷G��q�����K��+%���g(��O?�����.pA�'��Ru��?��d�F�h�/��p�K�!�����S�󎛟�w����/�s̻
�hu?�Ֆ!nN�3�Cvh��X�f�8睔x
V��a���;uCs����bL2K���R��B圉G|7��~�yN܆Zl��8i�� ��>��������CN�k@Y�)}c6��pz��ixӑ��N%��t�F�bf��fKM�]���9���P��cc,��h��^>�/)��w�R��zY �ѴB�r�O��"$�&��=���YRI/Gd��(�,vpv�W�;_���$JSK��c��LQ!�F0����qu�b�8g7C2�ۼ��Z��p�憑4�e���_9i!��pF�3[l��[�=L�Unu$��C�|/滱���\
_�#�h5��}��K��1�(��ni�M���%�l���VZ yy5�|��?��%�R��j�@�Çj��K�M[(ْ� #�KUq?A
�=�����?9u�Z���p1�;V�\O��?Tfz'/0`� Dᦶ`�4��װT�sȨ]�6�;�� �����`�խ0X��#[,C���g�jz[�B%0��l�|q�^J��f�ꋗ����Vg%I!o�F?���P[�J>�%���o�/\��<��.Ƨ����]-�� ���V�։���Yd�vݏ��rScgP���d��������6yN;N����'��[�1R���V�lE���:h'��`���1���1[Y���� ��P�EW���3r	uf��.��P�a�V:��q^����ݔU��������i���8.%��i 3��br���%n<�������L=�y �L|1���_W��[�{6�4�|��M
�Ɂ���8N=g�9��a�G�3?��բ�f-g?BJ)��5�Mx��C�{?�5:c'��XMBPN��FLd�[ոi$,���ܣ<���j�\&Y6c��?p�4pLT���E����skVd.k�H��:�v��G��Ӓw,!��u>�`E$���Ze�`����J[qi>o���^�����Qٵ�w���;��ٗ78�b�����
�Vq[�lX�/�gX�V�6��_�8
�oN�i��d�i׷���
Q�g,`��#H�u��mE��B֗��k:��,�)�H�M���1?�A�I;�z�"��Fn[V��}q����u�e�y�����q89mo�@�Y�b�{��m�党)'r�:%jb�q��o���25#p��`H4��Sq~���ߌ�(��M?��=L�:W����w8i���y��&� x�Xҝ+��F����;�b���%�jzM�C�$� ��?ao�%������a�l��̥t0=#:�As��̹�$e5�����u���1�\g�7C��#�[�R���_-#�%e��>G��HMǿ܏\×���ĝ+�i�e��j�c�X3��X<=餞�26w�v�����dH?oa	%��0���+("BO�DO�}G�ܿ�� �?Ők��;�t�Q��d Z^�f���R�/�f	�F��_�y�6�M�z�j��^K>]�_���/�����B*ǝmR��J��&��Ād�v��\�f�:��ֈC^�OSFB+���?�0j��k`�Ep?�&ßC	�<��U@[�x>�pQ!OѴ��L��֧"��B++&k�[�H�i�æ�XC�+\��n�]���G�S��I�ۜ�xν�,ŭ�3{^BV��&�RGjL=�~Unw�"�~iF�H�A,� �|�g�L0����4f�O����俙�J�޺��]A��fΜ}�b���=���s���8c���\̜@��B��<_��N�I�S�P�G�k̹ݍ��[P���T%G��=0L�wlf�2'�?��1�n���(��k����;�8�c8��N�oI��V�a5	85$M�������g�}<;��+|�$�$��&317���Ng�}���uy�*
��OzքTV���W�=C|�N~"�R�m讋��[<�m���hB����((N_X��I�Z�AC�a�I�cf�Y]���J���`|�zb�����7[7ns�`黡�i!WJQ�?�=9�v%yfvp����Eމ mҟ�I$�<b���r�j|}xlJ҈�r�G����/���3��]�gsP����!j�^ 1 ��jڻn��p����jt��\6`�}=�cǰ[;�s��S�ew/���͇����ч'X�E�B���U�H����Kpjꈘ�X�b��0�[]	��|��N�����Β䤷�R���ɴ3[�{8r]Aۼ��6w��&�	��H`�ⷴM%��Y��*� ������![��V9�D�u�/z�Ӑ	���PR$F����s
�(���v3,�c�|�P\�D�E��N`4{qP�rHMK��q��^;����=����7���`�9�ڴ/BV��ĦBf�^
L�Z�/��y�6�<=Ӽԭֆ�����e�|�<��fб)u��l��������3c�����;�]���8���3�h��}�v(K��y�%X�l(g�����(�iEg׋�+���s��}tJ5��&��}֎��+l��U6"�����6���w����=,�uF��A`���O�>(��7yt�:���>E�璡h����w/�X���\d���֪^Z�U�gh �o���E�g�m���bt��xv$�1�N��� T�)�Qf$��E�S~{���N�1ѪW�J�@ʫ���Zv��Ą�a��
�_:���ƻ�7�>4�G��Z�8��Ѱ��u��r3�f����5g*�����K�0��?��q�\yJ�.J�Ja޸�(����� T㙳�[�g����Ӽ�Us��eF^P�%�h���z��:L��$��Џ�f�ЌG��ad5/-��=��+���\�$\Ă�J_�����r4��lK�����
�-G�cj��Jt�D�:j`���XR�k�\��#}��ޅ�3�m�̶q�2YƂ1�G������\4���n�K�-T�a�	j��\�F��5x2�9�{�Z�Y;.}s��p8�PS���R�������M�V��=J���\�3 �am��ꯞ��~�af1!g<3za���r������	Z	�~�'�6��#���ƾ:���5�3k���?L�Bls{qC�͟f��zEƅ�jf{#�����M�x�%��ԇI��R�PQ��G��.����Zq�Ǖ�rm���f���"]ƛ�T�N�WJ��y����j�S*SA��Pջ���*���ꝩ�e⻓��0^�Ep�s���1����V½�cD-�;������{��,���/���Ũ#���u6�Lж6��*&e��{�\�gT���Ep8v��o���ȗ��eր�ݣ�a_0�v��[TK��3%�fvDr��e�Km�{��\���F:�
��<�n/���H�5���G{�MѴ�ym�գ=����bIP�{�O�+T=G���hLm�<�vAC4�JlD?`Tײ���4�a����������d�c��taf�5�pn���Pu�CD�v������W���>��5��)9�)[ Bk���2C\�� C�:�t@�5�)S!����K��)��V{�댒���
�/�&t��1�~8j#�ٴ�/RɳM�𕅷���Wz�_�x���v������^�&��Ba�nP�k^���V�E1($"���QbAi��%DЌ�w�sv��%�vv'�ƝQ�������(N*7��!!��濒����W$��Cj�^Zm��'���ݢ�gl��RI�]�v@3���h���?ݥm�Z���<�䤜\*�摜�����jO!������/|c&�� ��j<%f05�����m1DX ���.j�)q��#,����3˖l¦�)�P�m�I|Vc����s�3\�)wn���#9m�M�o�2��`�� UC��RH�yS~���F��@���0���������w�;��Oh����?�x/X��ʉa�몿��=�G)ڡA%-�b�e�?�3|�0�oy�NE��fX�노Yy����-'�MM�ޒ�%�4���޹O�U�V8�@��%Q�eK�"lD�s�"|���f��#���q�/��u����"��gI�R�M,%P�sev�Y��ξ�:o�g��%j��O,]���6#K����QHW���K�Ed�S7��Ћͮ�W[�g�|Y݀Y���pʰO[Ň�i�"%������fқ�[.~�bM`b�t�������g���Ci܃!�C���?+��^��/Y\g��k�A6c���$������)�E�la��0;��}��}��t��Tg���VG�Y�x&��\��k�Q<_�mk���g�p��!7���aG��q#
}�*�k�-4l��t����]����-R�ꭠ��sb��ېdB��%+�đ�n�xLcZ@j�������*f@�:�j����8���]C��>}�ɧ-�9�	��@q��l��?FV�v+�O�MT�СW��{��M�y���$s�&
��A>����!�#;G� v{�!5�|F����2�ٙ���OqZ�fa��j��g�*�����_,����u���g��,�/ӵ���$� ��E����3�ڥu�sIz�i~%��� V��:!�*��Rp���h`��m����YW��\Ӷ U�2�!����^=H�[�0!W%&.�X�{Jk
�>��0"�	=F�����Fa;��M/)+ի*іR�E���������+�!l�t�^��"��G�Ð �	y!�g��e,����%���+�-��8�S�7ˑ�f�u\�����+Y�`��]'�J%Y,>�uT�H�=��"�#�4\�;�L!�1�$j��+�Lfh���X��f�g�;5*�:�l�.{�[H���Y��5s��ttȉ����aZ˦����oӞ�G��.�B��O_?���E,/�br�����5�_O��Nx� ���i���`�����R�~�8���RBq�6w�ٙ9�l���6�7 ��/;���4�b��h��Q�Ko��2<�sn�U�r��h�6QA��z�XQ��MLz�B=OȽq���\xpyx%�ן3������.��`���o��K������4IƯi)왾����{���jK�#"�J�,9帙ZK4�,�z�7��C����-��"��تm�m�?xB�Xw'@`9�)��ҧJ|aδkBW��@t�E��[v�k%�� �����ߩVK`I���S,�Ӽ���eE���/�A�-lI�RP`g����%]�YRHj��D��ݯ�_%W����8GK�o��`�ׯZe�yD�cpa@��`TAS=,ѫD`ig������/d�kh��k�`D+nZ�5��>:h�i���^lnlܑrԄ&��.��S��|O5��{.���7��ĥҁ�N�x�#�Tr���y�C`�BF�"��k�Yx���G,���r�!�ʂ���+�L�\�w5��>W1f�����|�6�	b���\4X-��R��샂�[l� ��v�X
*�$z��J��k����jq��3A�c���[i�'y�X��!�6�d���&Q�,��0)� ��=��$�>w�=vkG�kkF|QM�����G���,���o��it���;J��9�n��]�?��;Cf��c�75���a��+�@���D3����R� VLp�u�Nn~�[�;�nBFK� b�o{����;X�/ ��e�`��(>S�r֔K����L����!|�&�^��� P͉D���5lH�,��un�q�I��9C��?��	3ɭ�tTc0��(�C�cٲi|H�%v�N�ϵ��'��حQ���{S]������^��c?���s1�66Ϯ�?��{<�(�K�A^�����~��D����3T���;o���j�5ҁy-�4����T��6�k�m����=;�-��#R�(��ɚ��Nt�� ,��o3�!�F�K�+-J�	S���<=��2���u���=�4�Q�Z"j��g/)��ͤlg*U�$���$Ѹ�}��2Ѩ9�b-Z��W�.w5ִ!�Ȼץ%>��Q��j&��V�/�QL���ɺ0{��͔����V0E�7N2i��0�bbc&��5��C1%��'P��B��v�Ϛe-���ѽf��sIϮl9T*na��G�sXÇ����㟑�'��/�Ǫ\�0OZO��Z�U�_��������x�s����,2��MM.l�n���5�y�3��Ϧs��e-�ĕ�����=�]sbʖ�ǯ�<"�ab쒻{�`	6�����G��J��,O�"A������
jQ����d����ۺ���V��O*�	����u"c�W	+����IOh����Z���#x�Fw��C�ΎSU��~>�9N�*������*a��,��z���\_�M�xm'�t�?Q�y<P)ԸA����o���y>�]"�0'���S ��sl*��`��ϿU �#��u�r.@xS{�*x����~g
n���o/&0CQ�T��qp�7�VMˎ(�ʀ]�����4eq"`��se����܊���jR7���	�r�i�]�5��v|�qg���"��p�Wi�gh���+���"��݋�����a��ITF�[�L���>|ΤV�j�{�_�@��r ��$̀yԆߩZ�;��P��>�~�y�� �Yi�i��re�g��9�b��|r=t"���:	�ŗ���aY�K����d�W��z��v��O�f��)��p��(���@K��
�:M������[�7�h�Z��~�B�*!k�8s7,'�t�N����0�I�����`X�I dds}�r�˹Ʌ������貘���Yw�^=��&G9E���{ r���k� ��6��m��'@<���*͈�w�>.j*�h�$�2�oi&o~�;y��uN���>��,���?�xp���hƟK!����y5e�-((�]�0
>���c�^��9aRƢ'Ձc��lV�f�?�]�{��@ԧ� ��ݠAw�!���!
QO���A뢿n���*fUF��;-�4R�M��h' lV�'�`8�G�״g<{eZ�q��w���8������h�O�f<�ۼ��N��j�D�5C��k��D��R��%m��]�z���vpX�����V��#�����M�`H��/O`�t�s��I� ���v��g|��(��Ruj=H��`�"���ظp��⾣f4�>W�Щ=W��#:$$^ҋ�̠�����Ѫ�"��9� ��R���>ƂZf�6����.���BH��N��@��� ���g6ل�JdjX��U�r���O�4�@��ڮ;)��l���Q�����Q�\
���y���c�Q��]ڥv��B���L�ǵ�HW��8�M�K�v����cAe~7����4$�1p"���`tV��t�o�9߀�#��$�@��D����3"�2.���Qy��������]���׹esN������.N�����:�w_`�d7ޛh�gֳ'ԗۇ�9�
�s��h�2�7���;���0�]��,��๦h�!�%���_B�y%�p�eka�o&rT0D�ѣJ�!���	�1�@��%�{���~TQ1����t�*n�W�����&�NA0���fi1�[�y��1�o��/�����$4ݗ���TjI�d����]�xW�e�jPޚx;�lx	�+\���6��詊�HAx�٘�BB�YO�k � ձ �� �d6N)���ki�z����g���x��{d�P�H�?Ag�ҝ�E�M��u�qO5t�;��]�;#�b�����{�,ǥc/r(��J��Q9~�r����=�6��~D�R�yٳRwYv-��z��Dg�L3T�\+�I��!���Q`�B�Iȥ�}n�;���jp�i�Pi*;��1�IZ_s�.�o�ZIՓ����G�K����jV��e�S�^|[S:��t���T�?Y ��ڽr;i"�(�1��������b�5`�{���b�p�I6�u���t15��~�A���V�������K���r����I�K,=�!��2/{L�j�F���=6��C�����i�m/~�������+���>k"A?���(B'~�f��/���[Ψ���\y����@٨��&�U�-��� M4���C &ʊ`!�=V��.d'�僤�)�z[p���׽e�/�6�x�3!��v�\q7�W�|��(�X�U��q�� g�b�Fe�^��ރ�0-��r�hV���2-#E��Y��-�%�F�Uv�Җ�ŝFEpRZ u?|�K!TV����ڻ��[<�{j��S�D���M�m�]�w��1�x��Oұ#< �q��	�RUM�:\�dN��t6�m�>����a���9��,���a�w�N#�dN�Pɪ#m.���O���S�*�f0QZ�?� �Lߕ�����9��%��Kk�6��H2r��J�6�Mhj�X�Ǻ�)�](�[:9_j%7_���,��8�z�p�}п�)����J%�{f�K�{6��W��c�l�`v�����z�y��M^��\��4�@m���K�r�9�5�u�t�~�δN���#��<q��*�X�G�_�nnE�)�P����c�f��*<x��J/��`�u*���>�8;3Z�h�X`�w1����}
T*%<[��ˎ{����Y~@:
NW�9�}�U�h��&��pwPM�JW�x���(��[ǐȃ�ʋ�MQ�����F�Q'I��ʳ�������O%�`Z{��կ�i�I���������Z5#9���4��J��YG�.0��
��{ ���$K	-�)8��,�.��?N�9ׂY%�{� b���q۾S��6�	܍�k^XƵ�6_ހ�]�>O���
�A9��v<����*;*�"�U��P--k�im���:_����ր�ڼ�L�u�ڶӀ%�Q�
]ޗ�{��0��8]��t`�om��H9��[��ԕ��O�%͢�U��}��]G��d��WIu��*r�!��2I�ԑ����Y�[��h��l�l̉
0c��yj<�g�Yo�(�>��LiHg�hxp���3)���������t�l�]D;��lf���s&�f�)P�o�s�P$ǇBE aѐ$=*6�![>��] ��Wz�d~���혝%&��|�~It<���-l�s	��<X���ˊ�N�DC�kJ�1�ܦݏj��޴U�&��τKѪ�|A�W�ߺ#$/���eHB:t����ڃia��x���Ԅ��(c�i�GD�n*����^��K`V�,������&߂���p!*������H7ӽd+�Ļ`���ު���@ �A�L����n�ʐ��gڙ���c�]��(sH�xo�9R�*�����(dI���Gᆴ�$垝���R�[�o	";^V�"��VM�6���Se��_�N�m8���.�����J��E��:f{ٺ_p�ݛ�q�m����t[=��.���î��(�7�������Eq����\�!��@S�p�Kk�l���
�7#u���Ɣ(@~k[;Q*tM;+ˢ�<úaf���&�%%�U���-�S+� P��v�&���o���$�ne�z��V����2�i��e��rڑ�I}���$ꇼ ��".-��&�Er�D��@ٌ�K�1�Ճ�P�����P�����9�<��^���j��?�� /�˒]�(��	�EVGƥ�W#�� ��i@�Qʘ憨v �ihs�/�D�̋�=�3�׵j�������7��}�����=.Q���:0Ν����l�p�0q�Y��9W��G��t��E��$R��k��^�{���$`���G�>�*GeU,�k��C���|��fC�ykc�!Fx6�����,�&��pLp��ё��~7����s̺	�h��,�m\�|qEN/X� �< s���B���j���r�{�5?o�U�a%���l.���������*י�0�_�O��&���.�#X�R`�2��Kߐ�,���Q�;	*�%G��[� 'ZJ)�y~T�¸ =�b��X��\I���ܵ"~Ѓ{)���'#b���'�3������~H� %����#Wഛˆ�����U��<��34�u�a�fvIl��=�qZ>���"nv�B;�so@Ys�
j�\e\��B��]6��u,#�a#L�Q�>wrbώ�U�yE�k=A[��+R�tX�<_��ѯ��rc��r���B{��D�ĝ$�acD��6����
ݺ�yE���/�_o%Z=yJ��>K�V��,����	�)�U�xu>��LlAD3%�QMUp��J���
3�m$���7�������d�SJHM��:С���HP���]=oJ�؉\�!�7d<�����
#\Y��AI�?53b�0aq�^�Ev�*	R�̝k�}<z�t��}�q�SU�����&a��	uJ�C��貗�ܿ�5�-�k{`��V~�m��r���T�?[�PW�A'Y�w�g��a.� �б�J��y��ԇ:����oD��S�nC���U�?t���s+3U��9G�7���RMiQ��1��� �/�G�/,v�&�P��L�t��ǅ/�@;��@�_�a�V(׹V���̯��7����]mZ�|g��\�r(��a���s{�z�P�����N��"z�_����m.�ލ�TV��<Q/f���$��'���E�}MzAmѽ+�E�g�0�Y�z�ag�=�BS���{ƛ�FFIJ�V)m�6	����aI��1F��4b�C�pΏ��cUL���������C�*(�n33�Kܢ���Y�/w��G��G�
H
EU��U?;�N��u'3LO1��.M�a-<��+*8-:�M�@աiZֽ�g�W�8m�l�aAT�^�E���#����01ԑev��[\����2 F2W��v���4�!���U�����k�&[��q��������:� 0��S��@lH{��AUv<L^e�~��g���K(Zyzz�U@�(Z7w�	p8,�ҢѪ�}�I�K��Ds�����ތ�p�J�;	����1-��#\f�ѩp��7E�� \x���Mfu�Nq�?���UM���l�}�n����c GFܬB��Y:8���s:���R�ffۮ�p#�q�s<)�#�4nM��Di�چ��%�LL2���DXgCD�E�<o�%PĿv�y?�˴�zZmh�xj��7�v�� ����d�d4�L	]i���jW�����9h���Й���~>�U��Q8���Je�ݤ���^�[0�φ˯�-Lk�	F�����4�-��v	�B� �-�V ��o�1?_�iR���l�M��	�FQB������kr�[V*���7=y�z���Ν���:r@�[S�dlhb�4f��U��.<m�!m�ge��2�V�S?H1�L��{���/��!��_���O�1���W��`����?��������W0<� �()֔tX��^���&�I�Ąe�*Vz��:�F�X��Q�N��ۘ7x@� �ݗ(�s|�N�{�EB���I����:�I�#�V�����&����T}@zz�X��]����zQW�&��v�Cg�1dvd���	�Uqxp�2~���M"9�|5hW,� _b�H�>P���_�뉞c����V�>ۂI�b�"`W��k����)e�m�Q������$��#zDް�Ӏ&����/v���RJi�U?'/���"Rڢdp`����X�%�%�	\�Z��`��WԠ��<�-�36ή�&c SI�;:�XKX�Z�'	�;C��C����'�Z[K���7M�`5^�Jka�ܛ��zJ�LO�qŢ�-�֑�3�O�3�3K0�9��j����J�����ӥ*[�A
�(�T'��#�� �ܐ�D��L�yM�y '|B�[���\�
 �jYl�3��6�7n�$J��[i���E|�C��N��᧗�-��P��6K�{��bD��>G�N;�V�%iDW�%+{s̃�_� 
	���ì��I�V>������g��vL��ڟ75$K�NX CW8�ϫW���/u���Kiw��{���T��;	|�y�	�K��"$��K��ش��V��8N���;��E�&$ m�.��s�gV�ac�C�O��<�{Ƭ�"�Ր�<����k5咀�%�q8o��%�"��B�4���U)���6�z�k��k��N)T�XE?`�m���7��S	6���=d�FD8j�t��K�P}j���ǅȳ�y����W=e��u��R��N3�.N�W/���F��yC�IF�F�(�!�ypWe�|�?(*sz�</�h"M�{2*�v�U#���� ��  �,��QR�1� 4g	�A���o��|+���,�h�̰e{y�ݍ� U#�΀+Vy/`E%?�5-�hRw���*���W�����gDK�̵�օ��7�QS�Cxh׋]X-�4���^Ao(f����{����F�uY�����Gkz�<lR���9Z��0�p�%���F�X'��.�\��ėe\���b�>�,�k����N��:���i�,��:���z�k7�Kf��x,m9ۥ�&�� e��irw_5ll*U�L$��P�tF��`[��}����W�����|;��*�3�hv[����@�,@��(����u���2s-7o�<�5���@+lHnw�!���GP��4�H��kOr<�I�>�a��&����h�[�D����=}�|�� �Y���#jE��~���RA=%K�?�X�)�>�Ȱ�!�s�+�ۖ�M9#��\�c*�'��?-�.R2I:m/q��'�c��K����*]b��H�,~�կ���?�5)��A�sQn27��8�NXP��q�@���2��,?:�v�8;�A��S*4�)�{N���PԿ|F��9�AZ����v"�.ʅ�}"��w��da2�[�\]pق�aP		��u��i�y�vϧ+&a
�Fh�N�m�d�JF����C��gƐ?���_�xP����������[�fњ��A|�0d$Q�D������Ţ��j��z���ﱲaY��
J[���/��cy��O�$ �Z��g���U�
�{n�R;^�C�r�>��yUC��W9.��L|�N�+JP�Oq���}���nG��1ð��H.�:~�T��L���x��t�q'�PO���H��6>u�N��80ʗ3ҿ}],�)�-�Z�(�(_�b���J�BN��qX]�Sf�W�����8A"<0b����y��g+�R���/=ߞ,�~
��z����PE&V�OH�$4�M#Kv2`1���9tu@�f
��^�������B��]J��H>"�uO<���խ����D��~&����5���O�~@����rA����v��Tn�y#q�SFU}x�3��@���3�)�zh�7�\s�3�@D�o��g��AL�;��h[7�O�����"��u$J�r�o��D��vM�A����w��fg���/$���nԨ*c)�}���q�Ӫ�y΢2:+C��O�}])fa��*;	ͱ'Q�g�~X6�D������[F ���9�AR��jэL��XN�&�|9�����N[hCpb�t��*_����-�!��U3�d�v�%�7,��"��t�������;�*Jej��Wm���"���MDe�)Gd�F�<(?����	-���7�#&�.HA�M���B�e! �m}�$ׁ��������?#T�;N���H��V����)R�;f+�f�j'�a�3�X尜��
|It��_�ü'[�bos9xt����	L�bG ��u�8!�3i�� �����c����E���a!=[��:\a/MeՑ�d��a4��R���q��*i��B�'�#�@����b�!rC��H�M�j��U�wŢ����'4[��#�XӒ'��No��,����	3۹S��EUBY@ ^)�,��)�u߭�#q�ZI�m��i>Z�����z<���R6����������U�z���|6��<tA��n��h���C��^�gAE�u����!��Ɍc�eAߑ����F6�\��:@�%%w��j���aps�����9����l�:@�����<��R��I�d�(^	�q�z�+FE%	��o�z�+��e\�?*�蓷�$�hmnv<��6[�m[�_��=T3���K��f��kz���"����_��(�ǚ>�pO!�tӫf.�<և�"�Gq��� �p�&���4�=�� 饏=yEK#��x���M�qG���a�?M0h ���) ��U��I�J�vo|v�'�"?̅�@j��G�PvT�nCtր�Q�6�R9�9fe�ˤ��$���*��-L�,��/�Rk�%��%I<���7�,�5�+���J�? �V!loC->��eG�^�����WSm/�cq��&�Dk�� f�u�'��7]Y@!٠f8:j��!��	��5�p��?��{,O߳;�o3�ȶz��wafB���> ��{8<�ڟ5,h	q���PD����1�I��p�W���#Ѵ'.����x�.�܋��v,HS��[P�XG�s.�}:,��v�v�g�DW���8��=�2�b��/,����=��F�C�N��CXb��R��1���u+�3#�QPXK�@�`��|���4�.ǫ���1"y�.
m�|�{)0C%��M˘%.��]�PA����1����rӫ�[��1~�P:���O���E�N�����"�w
q`��g�@a�w��*d�^뀴�/����X��Q�D"���+���؛Z~j��7��Ӝ�Ҩ`	��.m���{ｾ?E���Xg(��:�M�y\/>���db�Ga�V���[�Ť��&=�q1��*x�vuM�n�_.�rqA�b�IT;�gt���u�C�
�XF���˵z�>�y�Xz����|Z)�ٙ�f�v�X_ШE|N/����"݇�ʹ�o���$���ـ+<n����ZX��=��o#`�I��T�{ ^a�����%m\��(�{7����|��F-�wg*Pm��'��"�ԔRL����
lY��]���i�:��t��l��h{���p��.#D:�\��g<�T$Ow�9�p�`ׇ�� 7�s}���#��v�Σ����J8��q^�0]�'�$A��0R첱b����N&7��1⿽]�If6`�PD�,��i}n1W8��cr�2�"���zK�$C��s�&�>��<��G�FE�?�Q�i�'�����s��w��D�ZO����HATE�u꜔;S��j)�9���ȇ �C�I��Gɡ���	/zy p��c�JI�}4Ӊ��D�&��fљ����(�D�y�3����JY�mG~�KĞ�7�������l�7襣�TA��4��H��C�G�f��'Պ�����*r'T�DI����1K���G��K�w���K�}���J_0^l��㗣_�z�&|x9"�����	��U9C)<�Ue����%�T�5�u^W�f'�6Δ��@Uv�F�����Du���xg� ��y6�U����4g&O��u&�C���~���<r��/�Ǘ����őp�e;ԨId~f��n���7HiUe��¶���el&���m!f?�����X�`@=��л��X7��<�Xéҁ�2z�
���0F�������$zv^GǓ�%��qKR�0�v��79=��.,$	�&U>h�9��l��|��k�cQ�
��f��h+s(y�I����������C�����4�����F���]���z���y�N��0�ӂf��uٺVb�e
��6r������2c��Th!ք7����8V}(Z-9���'��NRp�U&�?S|�/ud���c����J���[�N;���ѨY���%����B�5���
ۉҜ�К-���^��q�7�$����"#�U�Q�ݺ��O�pN͚�W;7\-I�L�\��AY�<�&n��c8I TKR�Wu
�
�}��[xW��K����b[�nvV�{�jB��U�Q.����=%!�a`�vy��ě�x�n�F�����U��}V�	�|G:�t�.*�@�j�'������ F����=��Z���<��bn6B�F5e��$rj
Q�4T�4R8 =�(�B��%�O���H�3�㷏q<FGkj��QO�Wm[�Bq�8�-�Q!Y���\�=�o�F�kd}�f��R7k9
�y�J�QE�?�E���)E[�!���v��Q@oa��i�P�d3���*z)��X@~8`��A��j�����`�g˔Al�n�$D+O��F��� m��;�GHí6���΋F�>�D����O�B�#�������7�Z7�6|A��%,��gZ }C�OJ��HQ���Y��OJ%�&��'!���`Lc� �e�^���L��4*H�Q��a�K-�u�1�g�<;�x���$3b�^fK���*���#��=S�sr�\�8��w�L���gQ��W�׮�1�#���:�Uyzx��}�D8�IG|���\b��c�pH�u��_Ō��ud��?��5���:ߙ�li︳1�1i��l�r�o��\~���'9�"Z�N�x��^�i�w��i��Rd�2ĆJ ��I����&9����zT�z�P��%ܱ��]���y���e�r.����ܵ,�vϳ�cj�u���#z�'�<*�������aŅj��^5]�[v���^�����y�rI���{�V#s2��^���T�R���^��o)��2���TC[����e��i�i�l�w��',������fG��ʢҵB*$��9 �P�Zd)\e}U���W�'ݡ��k���e��L�G+�<���n�E-.y('�����*a`�ҟ���\@�C0.+�ߣ�檊h�%�xB��7�2�I�6�ٍ6&p��d�E�@g���V�z�	��س��4�D����M1]T>r�'�S��/aX'�B��&��D�ߗ`iY��aՙ���򷃝���a�1���r��_�ታ�i�O�$
{e�hs"V./��W�;�p}R�?���l�n ҕ�� �$�)��&�����U�'��Q����_�X>1(�<���v���Go��X���s�jIz�v�������и����tͱ�Qv�DV�J9l�h3��'�i6���%!O�G4�:�X��w���͛Y�`q���ɼ�&'q��R><��F�_u *c�)B��s-�X$��w ?���13�}y���́��,��.m��G��@y@|���ZO�'ȑ��#}:�����2�����`�`�V������%�j����D�'H09�R/<�e�ndF�T_ �y �]����� ��E��ԠJ.`l�1wˠ����A��`"�:\�8��T*cy�7�'{��eg�� "���Hn�r4h�{�2�
ؖ��D���y$á"�1�7�P���P�h��R�+Ny��z��Q��O �ƶ�W����B�/Y�Ы/o����P	��VtDNU=G�\� O�]�v ��x]�٣��t%�ﰤ���	�^�.���;}'a"W�4�%PK�b�2��RO(M �4����sti�D��$��9�A5�k��[�i+�k�`�4��]�j|e���uξY)	�Q�0�I�[�b�K�����յ ˌr�_G�HS�3�̭zZ7���.�z��'�x��'��`,3���8�/������v�L�GsW�vs�����q����Э򬎺A�8��w6?���$�mw=��{�b����*yʦ1�� yך���6�Sҙ��T�$�kui���ƽW\�m�_t7L�CR����*��=���R%~Ή�Saa���)�{���a���Ah.>�J����a�?Z�l�a���Q{�7��0h�ꃧ�WJ�SW9���u=Φ��t�e���|�s��}zp�s�|��ǎ{<Y��^ݭce�78��<Z8�����ƭ�1s��Tto�/$,����������>���
��y�w��8i<Z&��_�����y�����b�	�L����C�pm�ng��3�n�:yO�o���d��i�Us�aEoP�Jh�ތ����'�XiM��Q������1k�"���a�o�I���í64$7�h��3�
�o��]4��l������s���<���ӹ�@�����0l�J� VN2����thr�^bi�����j��*�d��l�m/�g%ӗ������pk�&�.o�(-��p�1�$����Ř�X*���NJl�?�
�:WY�1ȇ�e}���6�����P���:#�ӝ#����/�F�z� /��嚚�2گ�r¡�b�,$���'L��v���L�T_X28�3U�61ګ�Gm�R�:�@�qg�)��f�liE&:�K�Y|�R|<'�!'R�y[�-�";�J/�|�Ǥ> JL,���CN���y)Z���Z�R�=݂�!=ߡsd�}�U�!��t�w�m����˔C�&ͺ��s�>�^渦:�-k=�6�VvȈK>��ݨr�$�ﶆ�Q��YFa��ߡ �\uV�?�T_Ҟ�f�����r#ޜ��4���6��S��/�	/�r�P��n�ב�����M:;�.?��F�yz��]���wz�~�P��B�(��PdH��� j��P�迳p8�{P������#qi�z<�]>P�V�0��n����7
���Ic�ۖ���W���'��w�y_�[)w|3��_�p�U���������t�ˈG�L���=��e�>�e�e��J�������l���Tr���s|V7ޖ�V!�G��?���
�6DM��#�\�� ��_=���q�e���Q�_p
R����F@}3�7��Hp��g�Ԡ��CV���dt4q)9%3�u�	�������_68%کm���G&�����R����8_Y���_ ��z�p#�c�g&��Χ-X�j�ݲ�?
��Z���{`����{W��DX��P����!,���\��b��]e�$;(R�=\���d�X���d��3 �9�ˉ'}���%���'��lAydQ��8}�gO�,g���N%�(�^��6n���(`�M� ofm���SĜw��m��In�0�-]?�?`Ο �J {��fp���u��j�-_�����ή湧�S���v����ӎ�&`���F��E���aB�Γ�j+����2ݻ�0�SC0eB~�~�� ��i�6��C�t߸�K@�Zr��!s�X3�n��x$F�5��x���H�{���������Z��ǉ���&n��Қ�`"s9Օֆ�}���UYh���I=��<�`��Y�So/�x�ԗz@�rߖD�[�J#.B1������g��K�6�-�k�������	�낃T�c�>,��|��X�Íà�[��t�gy��@3҅l���֍�tL�4�o���j¾������PLz�����ať���Ɏ?�8���Yo.�3vl���f��E#$��;���MD�́F�S��xN^{�=@N|В���@�M��m��RP�FP�D��?� T�x��Sr��O���Ҹ���Š(�(1]�nR@�1�Lp��]�}���ZY��h�.�
ؙc�	��N8�}K��(�r�3,�+5FǽN�qVZY$
����{ ݬb�ږ��~d��[W�6/�_���F�t��{r��rS;�DN.�W"��V��}���|�$ʸ��m���)ѕ�h���ʱ)�PTYH�/��du<r�'�'I;�!���S-����j�����I��䨚��R�����Y�d<<��0К%�th�4 ;i6��>P��]o�	�5�o��ǂ��O3�H���	Y�w����B� V�%|Y��f�D��� U�>+�X)��RCk6��\ݸ3�<��ᓂ�\s�ז�xz��x!_-A�v+��)	�����j�1�K�EQ��nx�E�;M�G9���/�I+�Q�����������c\��e6���׺����w�|�[��W$���g�I!c�؝�ipi� CF���)��u�X�[�/�~�f�����|��o�ߛ8��h�kѻ|f�!���6����#��%��6��P�V�Yx�k0R�dڕg�P�P��,w%�q=���	�>(�(��,�_�H'ּk��T78Hh���/]|��̕`�y�L�қ;�-ʤ��@lX�o��<�T�!��Z��u	�vɔ�{�?w�������,aM�GV��_ك��"��L�Ro<����塕���'�ef��5�@���l�A�lv�:y�LbJ|5?��T��~�w�Jb���u���5)��ƕ;?	T�R����߄Bu��]65�𹋾2�P'�I�Ѣ��^.����i���;Ǌ^���h��uӅ�.�Ȣ���3.fg�@fVLB�Χ���G��W�KC�bTtK�qi1�2m��� �?��>�9�=N;��0��֯>V9 ���-@�a?��hz�տhnd�'����1��C��s�+�����29��N������G���o�t�!�X�6b�e����%\��z�C�����������&��2�T�
�����֭pT�8,�
�i8�dp��
��Q���}�p�v/����Ĉ��N���rZ����q�!�ک(v��,/�i��4T��i���3E%*��ק[����m7.��뼬yh�3��:a�þ$!�5���S��;|����e5���½@��^�JD�i��Q�6��X'3kh�����\���%3T97F���m�k[�<��1���$�&y�0y��IT�	J�1  W_�M�ⰧH5����k\�F��������v���Kv�}pQ���|���Y1(ksM�l������bby\�oi	�g�K[��=M;~'-����}��f�}�P���
�Ts�x���(�Sɉ~���7~}́����d��ܟzU���K��S����dҭ�$k���R�%�w��{,�90�t➽�E�|�˪g��v��p�N"ek� �&�dp0Sn5WRl,�O<�$օ��\\��sH�2幀�*I���Nۦ�r,F����נeK�ly5����7*~�!�����҈���+�P�f.:��\��e�a~D�� j//EE���4#[o���}`��]�|�)Ifa�Ha[��J���|��[�ae��oCU�K�Qf�'9^�M�T��(�,Y�GVGp��+:)֒���nd���p�y�|M]�T��Z�R���V2��]�D�d�g�s	ad����p%�k��=Eϗ���rIyt��U�~��_�\�R�,��`wD+^G�Z+Ͻ&����K��m�^Ó��ڒ�4�����贕C&�Y��?��(�-���[ߏ.n`|W�iP���������	̟\��4�5�"� k�����d�3LBQ�=/��1H�6sDY�����S�y�G��ae�ט���})<m`�c�TO6ʂ_
��c��t$6��ة�sW�Vpi���<]u�!i����b�f&�p˯�J8�.��������p�3�� 7�]H���0<-�<����ҽ�o�n����j�|l�2S�؞���)l3�'�X�z�,��4`g���@*�����!�9,�2 M �˳���� xɫ�}�HY<�����\�
2�q8d@�/�Pm8�"c��WY���s
����c�,�_h,�z��Y>��T��O棏[T�ڑ=�Gf|�V��~aکi�$���Mt���E�Iqռԉ����ߡ!�Y�j�yƪ�gc��cNo,.��-ڷ��cFc�_��I���Yܲ��R�[�WJ���r���KDfT�vN/�����[6\�K�c�s#���6�I�σ�N�F�`u=���3�E��ډC��Vx	���J�]�cq ��͙c7��<�C��1�6��?LM(��E�W�ӱ��}Vɢ��Ȧ{�����k�H���; ���\�G���ǳ0]b6"���\�9�x� s�#9t�	\��kь�܈x���4��,τ}��&�AH]Z+G3A�zR{WBQ��k	rdd�r�Y�CBvף�±���v'^iqu^dU�B������Fca9hF�ŵ6�;3QzW�E������Z��k����':�#�U���i�J�
��.e>��͓S�O,�+��� 3w&3���
�-w��8c\7yA��Uf�sa�_ryx�� ׳$����_�>+���n��|��2d��_�����j@Rt�Lx, [䂬$~�?8��B�'!�U�դ�12�s��&��/�s��[3�{���2�Ӟ,5�	���qe������ETC�&z���5Z{k�"�P�)�}^(��*7��!.��P���#�|��  �r`�w��c$��� (�Ae�/e����_�tբ�"����-�-sWH�u���Ǚ�c�&�	\�������W��@HB�|�@[ �Jo���2�`"�Q��D�_]����<Cdn��d��R1����X!z5����*�x���伴+<U��~�t��S4�|��?"�^T#��6 �+۝�����%4�5tjz�e�;���*鏲�]�w
aV�q᭭��i���×)�����[��_4c����-�b{��iُ|ߌ���9Z��.��ư���8g�"	�!���sg]���H��O#K�r��k��|d��������r����ɳ 5&R�n7�Fx����-Ren�
iIj����抪$A&�5�^���U��{e	����5Ni�����[���8�V�0j��k��W��}xt�ہK4�3&���PD��I��J���L�o3�T?�l����"�%Ȫ���k��ZPQ�4����?"0��Ź�Ьo��+V{N	��Sied�H�쉒e��[
��Y�)�&�<ڴ�DJuv��F�׹��/��Ռ����ֻO��cU����h�
`>�+����4�!ޒإ�2��vF��,�M/X�b
ǀy����Nť�MW���#-;	w[Tܜr�EP?p*��oY�ޥ3l���"�Y!���!44��O荂.�˖���Uּ?��i�fiEsZe;m�m6�A>��R�jY/�8�����}y����n�L\���R+<A��o_�d�OhɈ2_�C��\���QҸ�ߴ��O�{�b���{8{�{�.r]f0��d��Cc���G�
��<-Re�p0j/�F��p�6�z�)��۶�yH?0 �@#LsK�NG,]�t��{b�G�Z����d�����IP�;����s��u؈���A�"Y\���c�q�e^8��m6ȻrBD��Q����^yĴa�Y��F��$���h���%wz�֦����z�<ZF��X�����[�=��V,U�I++�&�[��T�qW[�,?�i.{Gt<��$�RM��@ѩ����]�y��bRD�D�y��n0 ι��=�3k�B�0�D/�ur2~ac_�|�w~V_�re
�ۗh[YąB����z������cj�t$�S����H-w9
��ߝ�Ԡib���S��_�t�X"�οO���z1��TdU S`c����碛�MS#%��r�K�b����<�=���gN�������DU6�N;�3:��H����B`*7x�>��
�a$��0����7�Z��1oQ�S�b*-9��	n��U�ɇ�c�A�%0�F����te�[��M���0mE�FD�yB�vh-9�賋�(�p�"⎪�ۿ���!UQ;���J�͌�$W�s��6������ Lۡ�֐4X�^��_܋&���f-����tj��{{x��´pQ7� L�(h�s�e��XJ4�'9||�R�kW` 4�C����'Qǌ!����V �^���XR�/%�+e=�r!��zユu���
,�5�a�*.�O	ؗ�߯k��ۮNJ�	�l6&�Qy��l�O�e��08�Sǩ�,�VZ�
��h����>!Z�����
IJy$-ob��d����|��26�D�6���7d��V
��1n����tӧK���X[��b��++�N����B��o<3���T&e�����GUIf̦H��ÞfHRPU�|�k�ڶA@��5���+CKN����Vj��\A��;��N�5.��m� R��X6�~��C�Tb���q���;�3K��Ӯ���B�z�DN��CDc;eB�2{{!�B��}V]i����ۛ���S��r	5[Ч�x�ئ^�� =�e�w��W���p<�w\:��.�ga!"�MN������i�D���͒��}Kn.���q���S��zz�͆hez�o������9u���(��)L�22U9��+�IFa�e'�-������U���[<z�߳�k�&�/����oc����V�ўI�W�[�I�Pҿ#S��wJT�� E�H���3 �q
�4ZS�ץ���w�#��7&Њ��0�ޱ͟׼��\,���3 ���9Qu��|�lӴ	��
iQC��c��]��b3��r��z��+����Av�ۓ��M���G�2"�rH���[n�\�#�;�ߞ��~�S�E�BE��o,��
�~K�'<�p�e�`�Lp=aU�Q>�9�4B�rYY��k�+����w���፧�Hc��3��T�\�i�	D�MiU�X�CA{+v#�9�T�i�K�R�4s��׮"|����Sˏ����R,��
-��Vgղ���ܯHa��̭�Q�ݚ�z������~�4,�(?����U
j��_��9<E���B1J&�0���GE/#�0(#h]��?��5��'s��-Ļ?���_,C�(�� ��?&��%H��`,@��Ի.�پ{�AQ�	�8_I��&z�'���"b�U3Z˧�F�.9�������1h���a��+n�E�N���d������2z�@8^#��)X�E(�} (G�Wy>G��A�K|##�6�����g� �#�v����[�b/�٥9:�͌�K�mѿz�1ẺHRf��������.� {�/���=��!��P��0ڏu!�kRT����VR�x>xg2�qj� ��ZШ�R�޵��B���n�J:=��C����r�K(�E:�.iO�_�*h��P�7����	)�#%�n��tj��;��d��*�:xͲ�/xxD�uѫ��[� 3K�����Ÿ���cl�Ԇ�����yi�{�]����%V�;Bn�:!i�yW��RO�E�K����?�{mw�±>v�� v�]�j-A��J�mψb��A�#�k�B� �2�vs��b���@��P�Щv�?�;����s
g��TF�K%A���~��3F�4�J]�h\�/L���p^�$��2�ʠ�tT�c�~�'��[0��a2�H��0�����qH�L�������ˇQ�}Y�!`�[0�>d�W��:c%Z>�fu`gT��!�Z�O���)C��z���Eз��M膓ü���b�I�q4�UZe`���]��{*s���8J�l�Ob�FCI�R��¹���dĐG ���f(�B
[S%�L�>Q�/���ǻ�����G�_�T]8�e�ݾ�H�쎱���vr��x���PB̟�IĦ��W�caM�6!O�P�ağ�c��Uf���7|&e5+'A&-��Of�ޣ�l��1٦B,�a�K������]�I��~��7�=�
�L�wS�Hw+�f�@6C��ܐj��>C��R�P�^N	Z�D[�[q)�0ʹ��$e�XF�
�ˊ���R��XN���6b0B�/]S݈o�_d���mI��}�|�����MX�3�K=a;���N��T�ڣ2�ⵖ˫�����t����m����)/�s�z��cd,���F�$���7fQ%�?�&A�p-��)�Gc<�^j��22>4��a��@��~��2�ů��[���6���vZ�1�m��z}�0E�k���ii��3�?�b�� 
��Y��ߣ~�`e0��Qwy�ْ������(�����B�Ӣ��-`=Ԕ�u�]��[�;Vf}�w��R0*��=p�����R�T�z=-ݬM)�R����
iƍ1m���bX����~pČ���<���e0M�;j��o���,�J/)D�G�4��+4ʋ�cm?�@L(�������,�y&B�9�[f�%��P1�ȇ{�x#�$�dE��,�J�U_K�/��Q��l�I�r�^�?�-ʈ!�5��>�&>;�r���.�|D�����5��-)#�t�� ��Xa@j�BG�ɲ��sS� ���#
��*�QIhϱ�����?m�0����K����$yWjj/|��t���YOq(k��o�\�! ��%}��(�`����03d�@%q0��%��.�=Q�48\y���ӕz�U�gp��10^�f��N�9���i݄[G}m�q:�}k�E�3����<I%�K<�N�j��O�.���R?$�H�)Y��O���//���0C+3�0c;}�"|iݏH�u�y�d)�Je쬰(���x�?f�S�+P "t)l7�])�*�S���K���E��Iu�����`���� &t[47�k�&��?����io�P'��uC��-��o�D�M�2��.�3�#�$<�ݐ@4��I�cR��N��?Y����4���2{S�P���q�d1��������W�<��0HҴi�|����A���rd�"K�n~;j�}EE��Ҟiԛ�^q���@~�5�P�q~[�3#��� �r�.6<�8W���s�&Ѹ�Gsl�i<��4!��A�{����_��5"V����T��	�������ƪ�a���/I��LVҁ�T����>=����*�,�/�9A@C�r�ˏ|�ѻ��3x���1-h�!n��]=�g9�p�O��)���HS�[�Z�c4��}�[k��z )�O������2�A�t�@H�KN�0""��[�'������������V4]C�C�݌>j@��#s)f���i��V����`�^����p����I����W܇!lnjsB~5r[��K��` a��Bc��3~���T.��é?�����S�3��-&�!I^L=�<��焂�.E8/(����[�e�w�й����aB����msy��]rʶ����ɦ�qI��MXFw�U��S�1�:�L���Z)�:GF����$j��V�(P�*].���{������QG9�J� �A�)Q�\}����Ԑ���3��VN>g	<$P�ɚ]㟐�@���'���n�zǾ/�x�' \NȨ9�U�F�s���?�h��բF�d���g-a`�n}��}��h��f�ᾝ2Q�mi�32��M��g�J�!@���|#�lvϻ��Cv��x�+dD�Fd��i�̓��Ǆ�h�۸���	���92�ܣ�*Q�9�y�t���o$�H+�H�6u��y�Z|K������ۚ�i�Fy�z&To�[�Q>Rd>o&e����Пu|��J2�z�����;�m39�xbv�<���v0��w������U���?�7�R����C���s�J���'�#��sڭ��c�M�'��Է��ŤV���A�;�g��I�<́��Q���NK�K�窙i�Kq�e CU�
�VX�������vU|�}VQBW� @Z���zw��r�pWp������X��d�����Ҥ��^E��I���;��J��&_rCƻ�Mcq���IR�x��G��ͤ&1t�r����W�qh06��wh��25��Bp�)zpkTcq�P]>H�N�3s��dz�a�&,�;������i���>�xh��p�[L���s^W�`EB���6C*91
-9����cY��
�V����q��#���=�i,��Do���M�GN���߾R˗�0����e���4����C4���1��]ՂYWv"�V~�YY)���ha�
�3;��&�n������Nsz��N4s�pw��Q1�a�bF<��&B�8B�0�l�c�)��6ߜ����%^Vv��K����8��C�=.��e�_So#י��o2#ahnY�̠T�9�MCz��J�3�۱�*I'k��dG� ÖW����_-�^>KR3Ƈ���d-L��d	h�f"����p�e��J���t{�]�=���ֲ�/�6���]5��i{��e_��rTe�K�F��C _�+�s�%Iy��*N��ygŚN��)}bک�*��=�^K�b2s�����x��>^Nf =}B�6sW9��:hÝ%0q�w�)�k%=t
e8A�}�@R����J���&��ţ���<|��}�G�Gsa�,��f{|+z���ƅs�``pk�����EVJ8R��>v�oƋ\\��=!��р"�^���]��������Y�ȳ��^fnU�z����E�,��`(5��>��g_A����ʃ�6�z�P$N�;�;}�B����f�O�NW�%�E/��xtmĢ��s_���z��h�ޔ��EV�AJ�� a��������s�3��|_���uP�6L�k���:W|�p��k(�2.�}��N��+W(K)Uq�ӋA�����#�pq�*�l~Q�*��i�C���27��0����=�'�<�~'ѳ<N����V��]�r/��w�<'"�[��	̦����i��@H�W*-���o®؍��^`/HQ��O~b��g*���}���n��sKDbBjR\t,~V�,��H(��q�HzW���ϓ����FK�>Y���h�����w��8�6՗�ӓqpf��.�w��N��M<S;E�J��D6�n�řr)��h͛Z#�؀��'��Hy�L-��9 ���#�u%�0'm&���W�A�� b�B�-�Cv�-
/6s�D�B|��x�X�u�7��:��l�5<��V�rӶ鮙uHE{���˿��)����ND������r`��c-�	�	��g�i��z>֛��z���wV�"-��J�(��%*�ٞ5��5�ܧ4�1fA�0�1�#{�2�����/�EY���N��� 2��Bh�1]�HVo�ƄHI`�]�8Ԑ�2׿!}h���F*
�m�'!ʣ+�������$�)-|�$2£��r����w�gђ�a0	��m1�.�s��ty��ؿdg�����j�8���4��˘RY��Z>^b���� ƴ^)���؇�pM�6�Z���"z$��&[Hd���B���p�x��Rznt�!�j� ��se����Y.h��l�q��oK�OsV�p;��A��G[�D��@�&�w�ﻁu}!!To*�X�`�|��ߚn��@��]c�✮��� t�b]��Z{�����s=��b l�W�_W�2�'/�ᨆ"�Բ�X�1��-eA�=~z��i��,�O�"_=(,�v����k]w�H<�Ξ4z�A����	ר�~�2���hx/	��LtW3�_�ؖ'm�'�dU��BjFB�D~���m�h�Ep�_�����I{j"�γ����',|��M�����s}��Ba�?���׾�da��U��ĴD
~P��D��a�C���
���>K�m�0�%��sr��U���i���?�h6�D��vT`o��(�{ސI��9J�ٽ�,�dy�[�Q�,�?�
��I=�U��`�N�� ��Q��H:��fh�XOg��Xl`�s�b�	��Zmţdo��u�zMv�-�<Q�:� ���V0��F
C'�B"�P��`�}|Sf��ڑO(U�W���C��Eb�>�~d��e!x��c��/��Lt�D���+��]��,�������5藉c���,�R�6��>����&I6bCOXգ�����'�����NXWդbU�QU	�CX�ю>TQ�.wp��b��k�c%6�G% jGbD�B��r:�t9Z,���u��..]�a�R����ArU�n������Ś]\[+{3�^�p�f�ǢͿڷ�	D�z�������OW�p2@8P�q���,�\���DbvA�d���7�G�R���wN�P�D��2����+9m�ʎ`�W.�y-�H8H9�����$�WG���\@j�r(>��.~��ct}�v����rOB�ZҶqt���w�=݋JU�w�8���}ө���WN��{J'�k���;���,2��E�݉��KRN!Td�-��o�!���]��Fh��B��
�lG���v��V�⹓p3\�c�G�f�_F�����B�Pe�Co�aX�P�zO�Ȝ�S�M>�]L1�Z��~��;_h��_Q������ w�h��	��U����&�`q^v��-/(.&�T-�p=9@o���W�7�R<����"[����j�<i?��e{�,�a��O��v����G�4S�ITB�1�M��gx�+���V�ڼ����� ��Sz�z�A����[��H��RyQ93�O�
���Q!�O�(�E������c���s�~����;��EA��l�~I;r�-�E�O`�x��RщB����*���Ij�r�=ˍ��i�J���L�e*
Ho�����{��x�R��7�j=Fz���)�{]�����<%��t͹��<j��N���stR$����*W���.3	�/E��%[0�
���;m?tdQ¾}aT�/�Tk3G�� ����i�Մ�3ˌx�k��V�Z��z°F�TX�J�2��L,�OJ����@MQ1�	�Ū#�E`���H��+�}�Em 
,X�����yq� �7���l��u����q�(�-�0��G�q������rߘl(�����Zx�~�1x�L��2:*c�Z�}��]}ב����+%���˱��A�[u���G��i�Jn�/Y�h���#��n�G�#�Y_a��=5�����D�f'Z?h�y�:�<�O�����3ǩr�_J�a��N��_�z���n���&���h�,�W�lP�h�T�����l�� �zdg7#��b���E����ZD� ':,{��_�#zb���*u�&�A�2�Jh>�e��}�OwEU��d���?���-^{0�I�j�Q:���7ӷ���9�%��H"7w�B�TR��kS���	�u*]F�<.��k�궕
	�%���D��R���`q��������za3���[�J{�<(���j�G�)�6�u�A-9�)G*�l��G�a�Z�Nb��E�c�E篑Tg����C���̞N܏O��9�A� �	t���K#b���\q��DԐ�!��m�kw�T��.+�o�X9=p,���������݉0��|؀S<>��������P_��!�$ܛ�:���v��a���^��3��mp�l��elX��rY�At@D�����3;�uy�����[�
꯳vԒ�EZ+[.y{o�[߳��QX_f�j��V>��T���ͰNÐ΍t�	�D$V����A�1H��������<�j=I�R�:5��8�ĘO��T���x�
+2�kh��I폀"Y!XH�لo��w��?S��g�O�����n���Qdl���T������Α���7��p���Ɔ��C=)V�(���5�T�ܪ\��K8)����a؏�2��S���Є����>���6ȁ�ZÏcs-ْ�� �T(nt~>������	qQ�v�<�/��:�1���Bb���a��Sw-Ծ��x� ,&���w7�}�n�sh�A4衚m=���}�x�v��r��x��=8�i���,�	��ezF;s�4c�,�]N|��_��sg�m��Y|U>�$�/tN�{���ՃH$|~w�ȮO�ÿ7s5��	*��:P{�6�R�s�5k�}���_c$w�79�%TaZ(kڎb�ò�_;fȅ�ޯ ���u"39߭*�u,�>�_׫6��1��'�;�S=#3�q�ڄV�5۔��܁�$u�q����)Zo�������) 4��x��j�w9Эz�v� �b��W@�gq��w,T\�r�]+��~��{�b�WM���U3�b�J�a} ��Y�5'ȊP֜f2��CMj=��l���R�@⟆��Ʒh�&rƺ��b�Ȕ豦��WK&�WÛ�`i�����m#��e�"(�w�L�^�L�1=;}C�q�t���>T��<a�� <~���jV��%cB�s��%��b��(Pv�Q��&[G��]{��^dG 
{���/';�/��{AW�F�[M�Z�Qcb�FV5���DeR�x���S#��D�V�bAy0�DJ&U[Y3�ܰ�!����p���
� +�Ą�HXQ9�����F���)�2^Q�{ei/4mcTV[���7^Q�������1ko�m��R]�W�t{uÓsy��<�K_7�K��;����8�/�(�iH�
�k���In� �_��g=d���q��]�t��'�`�]ɘ��������ߣ5�2�:\�Y�,_�h�C�,Jkl��<M����ڿ�����<!��;����j~E�k��UHu�5����'��6 �8���DPV��}�|�B ��g�ty���-��׽��V�����c�L[�n �>�U��3Zf��L��f|`*����3�Ǖcr��鈠r9�{���W�����]02/�t�q�������&$a^;�3s��iג=-�
��h
T��{ٹD�����Q%��Vh:- >�|Ë7�eF��0~�ѿ�D�Ɲu¦ͳ�����т�Ҳ�z�p�������)*��i��n޺��L�^Y�r/��#7�%��03�uy'3#s�'�NO;���VZ���u����њ�|��X��R)�m����/�7�rc��lU��c�|��\�f��k���\6�q�UJ�B��z+<�xl����{E�(����#V޲z��߾�\�X�]b�smi	7G�=�v&n�$Sʳ�Rfg�?h]���sU�����[���BI�4��8�~-(��f����E�Ӟ�V�A�\ܵ�޻�s�id�����jX�Xየ%f���N�>Y��lֺ��w�U�|7`��q;��oA����ɏ:��V4�h���Z��|�����V���S�H�Y��e�	�=�c&I0P��O_э@-�P��!~��h�����ڽxqM1�o��|K��Y�##��x9�S]"�!���r]#�޼�e���d|���V�f�s����Tp����L�c�j��ekՔ[(�%1�C�$̀�(b��q�o�ȹ'��;�z���U^��K�Ź�{��6G"�­��I�~�P��t����p��'N@L�����?��e*G|���YJ@�w���,��+�*�w&k#��p\��yhf�H1g�k�||����m`1�w�=�$���A}�����/Ne�"�U1�+�)h5k;&�4IK�?�^]���|����6|�t.��.hy�r�8#�*p����B��*KyhR�R��� �e�A>?d�R���&\]�XE��m�����F�<�E��d�
g�b�!"���B�@
�wV7����폶J��Jwxt�y}�ǂ�'�[��`��*�y_�pѶ[��ƿ�L�W�7+��ʅ�_؆ɼE�mKS��@������G\h�[�t
�I�����<�dVg4�b-ͣ�Ǵ��q�Wwk)r�US2"�3��PL�]M
���Y�"TL,�]����B�Iău9�7h��*�g��Y������:��]C��:��BɷSkꕠ���:��jOX��]��*YЂ'Q��>K����=4��'Q�D%�`Sc���cPBG�i� ��7�_�ק�-��fd�~ �0~G@�	�#
�4ގ
��Rf���2�!���Yh?mk���3ncu� ���妕�ϼ.sKO���Ro�4Z3���f�,����Zh��An曞	���F ����Ѫ��dж@�攟�o�P��
Ե��)8w�-��_���3�A5M����I�Z�I�S�3���et3sN78[���:���/�|����[y���c��qvR��2��!�tY&���� hGN��˶~�o4P�'�I4B�mff�U�~�q��\�9C��J1�<�`��*�k���vD(�~I����S+���3��E����J���"�3�Tr�P�5�o�|�����N躗j��b�^lK��{��1H4�:��̿Q�7���G���>Ŵ'��O�����_�}�`k�9�B�PZ�9:x;ל�¸>��Q�)x�d�k�jF&��B���ZȲ��i�
S3��l��hO7����<�Vr)D�G� zێ
0>O�&������To̲�K�^����jnpŅǔ�{-��p���>`�Z��M ���,�~�[�EBŃD� �
��4q���\s o�i��<�n5�e�����g��#��o���#���\̸D�oQ�[H�u�ب��,V��%|E�[�E@*�1��	���,,FT�נ�E&�Hې�c=+���A>QW���+
*�&x݋g�����<�7�U�EhR�9�U���%C�u������Vq�Jv��w.��g6�"�YC(\"ruhS v�X=�J3	_Jko �C"@�dh���U=��."�b�}u����/�m�"�']��[E�N��b��^>7���0���o�Ϻ���F�b�7�s6�# R}����~�r|`��j��]z��PD҇����oH��$�~���#>�e9d��P��
HI�2��&�L+��z��k������%���w���T^]�Z\����jՙW����]�KlVg�CoS���mD�P�����!��"vKڕ��X9�A�=�#�j�jPr9�B�!i5p�WeO�E�����r���gd݃Y3y��x����㙱8�T0��EgLs��yH��J�����<^oO;p_Z5��Ӽs���Җ�+݁.�N����	<���69���#�^�K����|ن����B}Ce�h"S�^�9���������N�!�6�x�5��!��E�e������P�֒S����`�i��P��@j؋�a7���Rm��i�����^�%�r�(�N���,�����|D�V�v�{dA���J���0�|�Eid\��>BF币�PJ-
�MZc8��b�S�[�eA�z�{7��p����{3�C7���3��K�U�y��@�Y��G�FFd�d\�_W~��V:J����icuWP�HA�4����{|`�t�[/����aD�2��do�o�7��Q�p�]��D�#0֭��s&�Q����X�[O#�F{Κ�B���9��nѰEվU�1!x���f�=ѩ,�f���r���C濄�B��� =�"��\x!�f8��,��P�C��(Uk�[p�R���J�P�7ê��6���1-X�\.�:w;�0�k���<K���q"�&K8��(U(|n�R�$�q��z�a ρߣWHR��!4s���EX%�`�&�
�z�>�� Xr9�#37j����`�O>���𷙣ī�6���.�:W��<�L`z}C��b?�C>��ܩ IQ�7[�7���1�Aأ^�-}�	��'I���i�/�uR3�8�+���\+��TIt?Ι v�"U���"^|17��g �bTO`�8&خ�kC}JV�M�A�]:�N���R���ʽ��\H� ��K�
*pgy�Ǎ3O�y��ls�+�H(��F�?n���A�y =ŧ�H	�n�Ѥ~%V�OQ���	�)��{f����>ȩ��M�p!)��i�ƴ�K���(���t�:�����*��nN�c��R��-�hM�+
'K�tq�`���ϻ��k
����Κd���I�bVt��[o����Y�A�Л�}^8�Ѧ�Y���\����1t�����;-��x^�=�|������D�4xĸ��k�QO?�$eg�C�[��yXj�����bE)��%R#��.����I�v�]<'��G�M�V	(?��,��F܋�\�.vOH��l��V	�fD�!N�^{�{��fX�L��*����y8;$�+)D�r�7X7���/���i`�1�70Ю�V
7q�I�.Ȋ�%-�I@d����Y� E�E I�����M������R�˕KIZ�)eн����xn�����{�(=oI��=ւ����t�Zˠ?.3�E�1im�0��c��=9yh�U�m�Qñ�zU,HPQ�)�A�hN�K�lD���5�� �}�z��߮?����� ���Su'��yg	J�y�&vj�~���0�i�;x� JaUͧ�������^��ͨ�!'��GwC��
����l��8��?���@�a�J-D�(�5u�/�u�h�{\v�D�nKY��TY%�d�I��=hݘr<���J�%RD�x���%	 ��`~RAt��<G@��%̂^��b;���:4���8�^��Q��v)�5tyd�u����?V���Ox��&�-�x�&Z7�S�U����s|G,�q��iI�~$�.D��~>��b�R��(Àrj��N�
��RX�(B�|Z���')���l�2JFџ2[�P2h�S{�,5�Տu ·��4�Л��%t8������Ԉ5gX��%�5.AQ��3�Q�o����RuC��%:ͪ�9�CS�������kFP6<}�4������@��H��#�x_�M���Y><lx)�B�.�� }��t�OM��#�ʈ�ѽe�4!{�"�2�Mr�hJ�p!n"�e�dt2����x�:D��l��S}F����a��Ƌ,GD�KX��Y�i0s�d��	g�OB�v�߸��P&L7>{�o�R���Ɔ��?;��Bej�v�6mdobJ�3�������)%Z��~�?lC���� P��4Y*��+{}���k��h"��2��]s+M��Ll'6�c�x"s���-c3Ǝ_�E�xԭo��M*�Ǜ~}+7{��D�s�J�������6gbu>�h��Q�q'��^7�6]b�QRԲ>:�U���/�a��˝�q��'Y�z#5W��D��$$��2�H�>'*zQ�[��ba�s3q�@ώer �*��>3��ة�2!;-���)]$mQ�V��:D�F>�b�끎EҀ�br	�J���(�Y�H$s��t�*G`[|��K��̈́���3�{?�H<���Aux��+=Iԃ��r@a�-�QqLkt
���	��B=��"b+���Aɋ^��YØFe$���ylǃ�8��(�����\���������X��I�܎��)��P���lD����4�%8�4'�hŷu^�ܯ �q�_�q�В+��M�Z�W�K�1��XS˾
�$=I�b��b�x��X#n���6����O���W'����Q{Bk���0�Ҭ�H4'�����]4n�Ť�E� ���pS��v!�+Z�H��J���U�hJ9��#�|�^n}�3nq�5'�Vl��p��+�̢�\�?Ã��R��r���=�ݷ��	�ý�ְۤ尗x���$�:V!�v�-vJh�1&�.i�^���Y��@=.�31�˱��S���V�*S����F~�`��y;�����t}<>U�$��N��bC�73ۀBzY��F�qn%`/ΗR�e�<��%wXJ��P�H�m�G�A��ɓHk����c_Ժ3��84���:�j���B�w��f������=�t�S۹N^��v��]ɟ3�.W�v�XP�&[bV�w^�q\
~��{�ߞ�_���]�t4
�[1�������%�Hʲڅ�p\θz���q�[	��Q�6���*s*���~���n����>�+-die�5"�����\V���\$����b�|��d]=����-p8�����{���c�U0}�	�@L�<xr��]��,����T�I���D��B���?��~���Irv�9���7����6��hS����-b̃.��(�&sgeB
�<HQ���#"?5��hni��߅KSV3�LU�u`�S^�l��X틍Kֶ�ML�����r	��D�4Ncgo�c��$}�HH����Z^��O���/�is�����FGD[0"k���ۇu�a2��{J��7�Tt$�6$'�ܥȩ�,EKd��~+v(���"��M�6T���;}��Tձ���N5zv6���{T#�y���D�S�y��3������|�>8�{2Y�+��	iQ���ЅX�$���?FR���)P����׌���%y��D���G5�e�lw��K�����}�O��>=�ƀ3�~���ٖzB� /�d���b��s��.��)�2e�\j�)l����4���^�z��օ�A����֓��d���k��0c���G�+)l�8�@�u�a���C���[��gΡ�pD�>}���9�N�5��9XnQ��N+M����0z���38�!;id�JJ��}��IfX�.|��O�g���^��� :!�ͮ,K#?��Ҟ���ð_dk��A�
�{�,0�B�E�
��8���|�cs^g���I���y��i�u8�������w��/]d�zRK�oX���Cq��-�#���D	.e�&�q�|br�~	���β�0`#���;p�!�<A��@��dn`�vVK�h�*2�΍�JK�##��i 	�m�p�R�	[d���8��*{X) �p$8���x���C�qE~hit'}Cf����,�i��#ceI��"i*�����z+�40*F&�Ă��a�j�]Ч���5���$q� H�֌�U~4q��͏M;=�hfb������`�̞'R���9l���X����~���h}�������H6m!?G�=7�ou���}�/T��+tiqh{w^i�U-0�k���ʏ�)�*���X�)w`u�R�U;6�R`b��3F�0�����:ћĮ������o�ޕ�*(M�[�;��ێ��CN��>D�=�q��%}��������P�y����_�t�-����t-�v+���d�H���ܰ�}�<�!�)}ukx��ێJ���R�4�="%�v�����X�<�)���ߝe��e?��� ;�=�cE��ߖ��T��2�� ��m���8���6�������,׹�.����ni���d�eMor+�S&�w��H6�z$���E������-����̛�=Ց��H0tX4p^��*r�-'�'�$��S��
��'෥5)�uÝ1���sO���
&�f3tCE@���U!�5:
������;�۬z4-�G8���v:k���W���-�n�����6irʒ�U�m�W=O,�<����F�>�G���6����"|Ε�4k��Kx�8k��#�������6{M�M�*�� ����c2@	$�Ԡ;�Adi�!%��$�R�\w�Q��瞫.4e�N�0�z�M��,�����1���"��9d��8�R�S��J�G���'�mQ����dJ�(���Ɣ�e�˫ ]���!��(�/^���Hu�ݤ���AǘVN*I�NjJ�f�}����8�i�b�d���w�[~A��IF��	֪��F\'���������;�*΋]�+x���e2� H ؠkNMg�6��5�����}��-p�#q&���K�f`++�� >qP�ǁz��s�Ӥ<�o�W���@��c�1��y�DWT��'��כP��9��PF�K�N���2�]�w��r�� ۙwj�E���+��	e�;����u��	�Z���.�%����R�,�����c�O󨨸a�)��*nî���{��&G�C
$/1W������������Ѧ�j� r���%���?�
�C�V�v	86El�r�&e09��Q�^2���ނ!Y��/��^E�#��D4�����+���,�)3G���QQBt�m��@4��f�Wl�w�p��H6=z�^�؃��x��y�+��Q��D*U���]<�m��D���#��?�}�A�W+�'��Sy��}�d|8�3���x�<���Y��R::)Zq|�sU�?�`]��⚖c@gR�Vѐ���I�ڀ����Sx̵�!Ў�����x?�:� ����G����kY���x�#�R8 ^�Z1��]6���٣�΃["J[7�"�1E��؉rV�W!C�(1��(<ү�ޛ1���%?|=��P0ǑN��-G�>�/F�V/ka:M3�pE�P<1�Cn a3��%K|��T9��B�d�����FB�0,'O�=���<fn3��$��={����.�L˛4�%n+��'j�O���SL[�3#������qI>�G���C0<3�Dv�+�����lF���`G�bvHQ��=O�j��N|��X�E���6���<h+��!�b����$!�q�+��;?v�<�*���S�g}��Kq�_�ĉ�~(���[��E-�h�W��X�D��AO�r�<�g���������:��7�v��H�S+������JH�� 3ӭ{��G����SQ�z��P?ˤ1o-���sXĜ�>���h�$vOD��Y�Tb�R��DuA�GG)��w��nv�+7t��<����s7C5�w�����ݼ�v���I�7�'�rK��S�1�j��SVŋ���ڛ����e���I���,-�m��)��ʹq��{�T��3H8J��Md�a"k��R�f�'z���#���[W/�Wj�0���q��򎏲�	�s�)J�j$���
j�L��{y��Q�Y�P@*��>V����E~q��B[�9��7�*j�f{����l8��Z�4�?���*�h�e�Y�`���l~1jr�NED�.���Tm�~Ɲ��U5��m��F�)�twH'�ڈW�ge?a}�	N��L_�9
���Uvp��#��	��*�<5?(9���%�>��o�-|v��-��,d|���{���Gƻ��ȩ��ԟ�� �q{4�U�S`��@�s)��c�ʰ�
@�ܶ���Hc%$�I0k�h=�A���KS��85@8�#8�p`4�TtMjB*!`�wvu��k��a*4�K��`_�����M�ƉG��<v�96L�]����q$��+ ���^0����vvF����좾�vMq�_6C[�:O�+K�+�I�zl�l����!Aсb%�L��&O�P�]�*Z{���8� ��߱��<���o��b��&I�A�AJ܆D�ø��3��ϸF�q>)9-/�BQ��]�ˬ�h����wW��<n� ?����"����D�K�1�D����V ��O�]�����\��<~(Wˠu�!a[���ơP�t[e�i��*U�(��*�r}�N\+у�0��+��#S�WB�0m����[��!	f�S��F1�r�*��u��y�l��ɩ��r�2��_�ؓ��X��鞤_��3����������Ԁ�Nv\�Irg}ǘ��	�pRK9wɆ8���� ��l�[t�7���OH>��-�X5�Z� KW�]?6qFqA�� ϴ�[��aT�L΋�ds�W���x����W*d��q��H�6��q�	3��^��|ǥM���]ݑ��E�F҉��ZP���_2m$�m�*�!5+5��ܙr;��x�����X�SόV�|��ק.��e�Vfŷ�i	t��9�Vˮ�M�_���r҂�=Z��!_����xKQ���rݪBR��Jƅ3�eh5�L0�;c�������e�r�	*J�]�֭(��^�_	��$�*��;��=�Uv=��綶G��X��s5#��=T¥��z]�f(�8{��>S��=ͥ�q�.��]K�e��6����g$���J��͔Cװy]�`��p}�gp���:�Aiv ]���� �f6��Dve����ܶ���J�I�٢&N��bQx,�
}��P�ɡl��D',V0��zm�5%����(E�}��l��Q
	%���9�s!L��lQK�Y.M#��̮��gv��]�L�R�iw[����5/��8Oi�ݨ���IB3>*
0m3kI��T��3�
D��w�h0�T:�l��栧$:hI��l�Ҵ��KC��S�G�D�NX�I��
$N}�fzڈ�7f���dΤp�pB�����[(�������+���
�)� ��_�P7:�� �V�vӀ[���4Xi��BR,��La���
Qf�����Af`6����	��б"a�Yqe��ӉvB�[ހ��j]ד�)��D)�޳P�NKl�;�7�y~�<	usI�	�̳߫�u;C� M��g�X�)��̴��y�{�d:�H��
`6�'�j���Y����1
uc�`[��qm�v�p����<��6.�R�MFr��6��
��a)��)/5R~+�	�9�|������΍�zL�x�Z-~�)sZZ��U�n����x�t�4���Y�L���Z:oV_G��s��� K�z
91c�M��P�N�Q�:����~��n��NvțS��V�a���×qH!�>~����eK��3�2��G�Gy����QN�/qE��o�bl���6�z��IwzE\��`�'+�����^���j?����"#$e,�\Ra-��YC�V�/2�Q(��{�;�1-Yj�Y�ºʫ��R��D��W	�n�a�T+�)U/97���qz�L������B����/�HJ
3^���MfR�C�T�Zh�?*���ǩI�9-�c�Ͷ�A�nn�BA���c���H~[�壖�����;0�3z.D�1����kЙj�k�FQ���t|m^��ܡ��OG�n6��72X6��R��A|��"S��}�r�`��]�Ų���c�ݲ�l���l2;��.y����+ S�T=ߵ�D��0�[�	9k���a���͂��SY��I�8�{�m0ʟ �ڼ��j>U�SE��}j�.R=8����]��]��>��x�J�Fq�x��<���	փ��Iw��������>�5'~���Rj����.w �qp�"�b|�pp�r��7�_k��0�\]=w4+=��<�����ʧ���AW��z�ݥ�{T	�}�_��#b��37P8�3�L�-����7�93VH��%���&^I����6*_Z����E}����\�
�"@5
f���@Wey�$�B�_�,v̶\�?��o��ڭ�p��%�O9%K/�ƙ�.��I�B���=��������b�9*B���-�u'�F���Zm�0�\5G'}	[ ���]��"�f�0zY���������X�͞Mn孶��ֵC�:�����
�ȫ����"=��Y�}?�/�6��j������.9w�ۨ.�����?�;�
y���~����ȳ�:W�I���m���Xr�����s���'����P���{�=�C�ҕ��4��ʃe�@@�
�̙�0l���I��3�_��Ou>&�k^�2bS+��`��o=�ҪZ�{_�_�QU6�i����Ri���m�qEWMK�٦�j˾VLv��Yc�?o�#�64��t�A���%G2�$�;@v ���1�o�����(X|g^���2u��+�#%2�@%-Di��U��kf�� 3�ܺ��H!$!2I��ڗF��g�x+L�Z�޳�|y���k��pʴ�Jywd�����2g�zΫ�a,xI���L�l��\���o@r��7��#��і�\��"�e��s,��x-%��]�dk����`Ru���de�Qל��7��'����6O�y]����%�xFK?��˥[l��e3���	چ�i��a�iM%�\�g��QK����>ɫEW|{y���Sq�>WZfS��t8�`>M��#_��{R!jʨq#iz�`�ĊpT�zE�Q��07�\��y!QH8�ߕ��_��DR�6{��f$�"�/c|�v��� &��i2�=Y:���I7|�pXǓ�M��F<Św�S���>�Z�s��7G����f̰�i���bl�������P��b�f�Yמ��:ӫ.����Q�%����͔K�VrݧA��U��!��K-ľއ�/�n��'A�O��o����=�������?<�2�5Z4��3��(:L�Ȏ�F$�	����c�q�1���D~��dQ6A*�,����&��r5C=:[���'��	fh��u��b�!�[��An]\]�w�B*E��<���ֲ[jH�5�N��۰|��p��n���>Z+�'> �U�b�]��-}�غ������8oX�@96�	`�9Am '�˹v耖�G)�k���X`�L9^a5&^��h^��T�o�b �p�7V�Ў5�p��{�)D��`�j��Zg9Q`���_>M�H5��]�C�;��&�nM������/:�w6�������%���F*]\%��������G�"��~� �B��D����2��V�c�q-	��E����<wU����KI4�t���؁����y�K<�f���8aB��� ����c0�wB��V'����1l���ݨ����������j��R�s��y+�R<9g��ni���;��5�Ĝ3��{R���!1��ya������Ԉ줔�u�D�0-����!2 �r�EB�pЭꍒ�Y��y�BnU��'k�@�r�u�D��̬J.��R?u��j L`;c1إ���*H#��� �|>�uceU��_}�%��&���P<@^��`�i�
�k��o�s7t�4�yZH��>��P�w�L=%/z�<��¯�8%+/O>P3I��)&r�[so�T��ao����<-\v�8t"��%���ƛ՘1�o~��d��?�\x���F
�t2�h�ڃy	䧄���M�|x�$���M��@��Y�5E��ۖ�T��gj��� ���ҏ����a̴+��ւى�- �
����B>,]5;O���f������Hc-p�O�/u������׫�fWҊ��λ� �!=����bE{��K@m����z�#,�-��c~H�� ��<e�Rgc�����_:�o�]�����xU��{�([�욞`3G�);0����}kh�,��9������[-V5���`/P68�dמ�W
��rbj�&�8�Ej蘛xf
.����~/|4��4���s�C�Id�*�+k���21D��$�����hpȴ=4Ō�e�p���V@%��'Ć:j`�w�R���懦�o1��KZ1��I�(���_�_��_��^��O��ֶ�[�`n�>99���|d �Y��Y	5p���h��Ҳ֧�� _O�R�yA狞\S��kK�vX��/+������N��u�x2�7dy2��9���+lHVSO|��TI=���p&�ۿ<��(�Bl��?ϒ{լ#�lȈ���w
��ʔ�G��}�N�:X��`\\n��E���n9�D4��P&�����:���X1���p���/I|����w��R<�'�Z� <S ��Ɨ��ԅ&�\q�f�Ȉ&C�ya`��󾻩�A��i=�/,��|]���U��&±�<�>�Ҹq\��₎�i�- !s��]���e'�����0n`�W�����RuB��� �v�|��,Q�y�7�1�e�ѕ;N��J�l�bJΖr��ʂ��>lV[w����U�G���r�{�),gg��q�����^�Y�P��v��)2b�;/�b��O����Ƣ��4��7����*��3�%�kѦ�uj�Re)�����Q����U���q�h�`ݟA��r�e-�h���2�Pk~�AY��C\����
t�K�v��uJ�z�i��@e ���_g�.y��/�eL�y𲛜er��^ƠBMr%��*�)r�?f���l}���L��7�f��O��2��=Gp����e��U�x��N����L��ىւߴ�U���$iuest�fƃ|!}�.,ͽ|�@5���A�+!�2��#m�?#�%	��$������ݰ��4��O:�����2{��*s����Z���qm�����&[�_+�W
���"|QN��T�13��p^�<��_�2>�ܬ�yJ�[��i4��h����[�qs���Mg�S��W���ʹO�-�n@O��4��W�S��!+H����k�V?J���W�A��}To8Փ\���v�}5`7ȸ��_�'�x�ɢwFu�R��|@�J-/,��/�TV�-l5�#@��+�7������F���ڳ�$��NHw�1����8�ۨ���6��U{�0�#tY��Q�<�]�!۾.M�G/-Hy��p�Mk�n\� b4`�~$�Zplw�`Ѩ�e�ZuY�U�=�����걤 `jb
ݚ	^*�$�Ñt��K!�yC��@"<wO� ���H.��� .�cs�i��2x���-�W��?�݈M^!(�ڬ,�),f7�Cw�r�[l�D����s��	��������nI��>*ao�ty�CӹR�^�f����;ݠ���gbit�0����7)9���+�D�:��e�@R���i���p�>���"8�ȃˈr��a;Fc�>��-��X����ׁ?���{�z�6G��C�1 ��:k8��斗�xvSq"��B����6ըi4�k{�;����kT?8t�ܪ�V�\iM��ȿ�%�����d�2mD�Ͳ	e�<#W�IP{I� B~D)/i������,���
�A�/�I+c([<ْ�C|�'��	�id��ͺ'o��{�e�e�>���i:	��<�?��:#�|(��-�L���}��n��wz�J�E�^0�э��9O���[��~��1ޱ̡����=���Uzh��~'��D�iI�a��CH�lO�����O��l	e�S�SZ=q_���/�y'g��8'�O��O��Sͨoe��^��_���O}܌L��˾ShMI
n�r��)���3'(+rRk�!Z@���7��d�3&�8�7��;��~���?��{tC������=W���q�#�5
�?v�:�8�}��P����P��K��u�S6�czKA������#�ט�<���c���m��A5ڦ��k�
[����z����vW��	��I@��r�ZI�4�S�z����U-q���B�1��˰������6?���`�p{ s>���R�=����#���7�@k>ë�j�oN(m����(�3)I���d	�\Tݣ�q��VK���/<�e$�-���jS�0C�*o�����5�"?3�9 ��+v��Xʸ�%V�����F� �c�Q�DA���t\�\��F��j�G�f��c-��`
p�d�����"��2��F�$�8ܲlM�97=�,�1RQ�g.D��AUD��k�����GDfe�5=;�?_�Eٹ����l�OOl�TDu�꠰�ϧXUo�q�Nile�Pl�=�O�?��Q���'c�ȿV/j�����旸/�#d>��·�,�%����$�����4z��!��n�t��5��)�=��N �8�rh��~��	���-��D��L�_��ZeO����+��2� %ܡ����,���wCb�s)�^sP�_R�u�� q���˼�N��r��L4�ShT�7}�j�5�r��5;t;�@���Y�w����X�+C�j�2t�%x��=�D�(�+8��� w�m��[Y�A� �KA%b��sȅrC8�C���ܝ.�ظN̽���C�[|e�*a�4.�y���oDZ�:����YZӠ3�HX5��!Ŗ�p��q��/��eź@�s���Fj~W:���Ok�ܣM��O�L���QUt/�~��Fc��JM����4t.�#*��L?�mn'0OaM���!8�ٓ�?���r���45
`��~��eI�"�;���e��x
${dA
M`ܾ�c<�6k�`s:�;W�yo/�v9�*�j� 9�L*���EOW�$�u�ejK�i���S�%h�"�vC�< ߲�<����V��� ���v������F�[�zb6g���&�&�ŝ�V6]�0�DwM��lz�C���3�K�q�.d���
㴐�?zt/������<����E��yfGt>T�#��ċGUj§5��b�U�8}�!*�s��?�!��U.�q4�=`��ig쨅@\�8���g&��x�m�Z�֤�l���y��@��'��ָ������6~.B6rT$��2R�P�S�jه��H�=��9!���WoCq��Nҿ|��?D�}��r�@.i�F��F��? �:[�w���.� �������lq�s�B���'�S2�Y�\�������B`$�3y�W/wNw�
k_^`����?'A�̐ ����'�-ꍆf|R� ��R�������4꙾�u.Ʊ�+ 
�3ǦPph�r:gwVJ���')82���s�D	y~dD�a��i�
��{U�js�mX��TX�������j:й�UWX�4 �/��p:V$�6��KC�{� P}�	�8�$�4�xƗ��(L�X���c�6���e�?ǣ��P�f�.g��nD�(R�/H�c	cRE;�
3�.��Q�����`C{
��e+]rYI\�Ѫo <Lx�M�!7Ŷ&]wA>�^�l��tH�L�g����/_�jL�Y-3o9$�uV���X��Q�xb�O�eF���nf��]�c����lF��}5C�Ds��uX�V��a��42$�T��G���i�`�x	��ɹVvE߼Z�}�?*�B��o`�*]��S&2� �z����3}k�^��IJZ�qo�B9��Hx�����
TA�jVă|e�n�	Z ���B**�ʮ�?!��H֊d���M���
�o�Eu�<���OM����Q�(>s�cx#��u� �'�N'�3������l����0]�\^X=MU5���r��Z)�B�4l�3��ʅ��j���m�L#�3���Z��I�#��R��G\��_��3��"%<'I�r?}�~��%��䎒�K
/e�qCИB���/^�~�cJe)E�O��|j�k=��Y���C_r�[a��!�Kg��C��`~���˰��H��ً4<T%�y�B���f��8��+���i[ؚ������Vy"6�5L��i��N�/�z�hV�87�NJ������c���^Q�U�!�\c����*��\	��&������@ї�i��������2��Ɛ�mt�2�\�Q��a��rٵ|�,����?�H)�]M.�GSQ?ә��҈f�;��/����۰;qH���8�=��1bI��t���i�&��c�w[�r}?�o� ��!S�i�:������\�����)�NJ�i�II����{���+�'�-�q�軴9*��t�	�~އGS�S[���c�F�0>}�J`�@R��lsf;�fZY����������η�G��iG���Z+8<rG�S�@F"����>1&�O��fe��Ou���K| (X����6�b�L*l��&_��l��
�61�/�8u}<m�'Ձ���~Kja2������R�ׂ!H���k5��O�L�u1LD��Ӕ���6$dF{H�xI��^��V�J�c=�JM^ Y��v�����.]�N\@?vf�rZ�SwǏ
p�67���/B�kS�0���["���/D������S�RA�Bu�!�ׁ�L�>�9�w֨�e�FCTgx9{TU�&-:��/04�i�R��R1/&��V.�����~��5��GN�G���3��޵�Dg�cyD'���D3�0��9-��E����K'Z������cl�M��qv�V�hp`���hr̙�61"��z���;�BZ�� �2O�[!���:��s��-};O\��g��w�PZ	�%%=E�`��3��̷�K1:���Q Tc=B�i���ޣ�N� ɡ���z�F[B���z�s�9n@}}Ϲ�Q?�B�:)lfBt=�^�6e�U��_��i7^�S
��/�T��}RƵl��l��D�$7L$s-�6LD�&�ܩ��cO>����^n�ʠ��.,ͩt��$�KT���.��ℱ�:��Q�
�xV,@nE&S͐x�A2=R�x�؍�Z#���w���Ȁf���i�{9���0�#j~���JG���\T��9��yi�L�`�C[4�#r�/����X�T����E"Q��m�����U��͘�0n�E�5��b�*Q�n,�u�#����"Z���W�{T�Z����7�P�F@�C:>X<�3�K�^���L��b.�t\�$���Z�	�{Hx��$P�]C/I�¸��~�D���=���"C��iF�K��>�f�K�os[V�:hh�f٨�����*�
#��~���1oߏd�L����"�Q���Sʍ���:������睵��2 �ڞ�:�Uv��}\�K҂'<�S���
�$*:qD99�U`��֥Y�\h2f�y�Îw*�	�+�R�S�����\�!�N�0
�{�x��{7�!'A�@<ۙ� ���}�c��j/߿�M7�?p���7��6L�Byd(�c_�;�-V]И����@�(�aÐ�5��`�q��/B;2����*Q��DY�rI���KQ�g�4��/gC�Z�\�c>��[��Bh�ւ����H��|4�"3?&J��ɩ�m�b*��_�qeNsY�u1'BM�����\���u@k<�߄��O{�eN���(�?V=�w:�K�x�C�(�p�Ao�eTM���h�H�"�_*�F�ꠧ�S6����+��� ��`�|:?�h>����._�RN5�I���3��2g�	'�d����1���p�j�z���o�"�)Y��I���H�%�ؽ&���
/��1��� �v��?��n]P�3�����ƌu���
�=��U���01�����uʆ�D�eog�ٝ�r!���}*���'�	�O�'��$�/�o��U56&
k�1[��c�<n��l��������2��6��(�!-8Ъ��s �g�w�Y�U&{�a�ɼ���,�7���kޡt���~lm�$Y{o��~v��1�xش��h]g4��{�Y�~0r��K 1�t}<���z����"
q|
q��2��\!�W�
�3��_=�_|���f�ԁ|?�0���	���@i#��뫡��'�GV���̼9ai$9KA���b����9
]�pM�cJ��*'�N(�(�F$�t��f��B���,Ͱ߲uU�.^�ޤKFLc<�Mm���bWoƫ��y��#�Y�S∺���kj^�7Й7*���ON�_�LS?fU@܉�/�����yH����.�$2��< V���D��~�"ǌO���):Q5�3�*�轆.&T��,��;5K��=N.��hճz¨
d�MR����:�����#O����c_�/��	Z��O��Z�X�5Lo�t/��l꧵�E&��Q������[z_[*N�k,����V#߭�ކ��!�Nh������.��aW����"S��?� ����бs	-Y4thH���c��]9��	�N�DE#�{�ob�(��Ʉ��-�!�Ї\���fe�>�,���gvV�w�I�l�M�ܢ��Ӎ:XC��1���9�b��d�y	�a`݅r���%�z&���<�:F�����PV��]	�pq`�����Gt��ҥ0���ڍ�N��2�p��y�-���4Η��8�ԆR15��E��s�	VWڈ��ƛ����%3HХj#�أ��N(�=�^���G���`�k}� �7#��r�����a�If%�k��C���-Hkg�4�v�$@����m��IRU���-ҙ�r�a��M7��*5�F>G�"c���h�7/��rQ��K�1`���ք_BOb��c�Z.�=�u]�ݙ��7c�@6ȩ�_�1#�a�"��$���fv��GA
-.5|�q౾-#ǳt�e��_.!ʸ�
���88�BU��$��&b,�q�Y���e��Z����<^h�\4�
��E����N�D�9�}r<��l"ΪI�77��<�+�#M��S���8�9��V�!���oV�.6�ə�xmm6�(c�_�W�kHc7��kډ��'U��߾� 3��Ŝ�	���Ù���d���E=��/��!xk���"�Ꮶ���u�X/�N���K����)��QQ}�)�y�`�\;�tzn�u���,�2�W;}"����x���� ;�_D���R�K�Զ��v���w�G�#
�J@��ݷ��3v��p�I��{+P*x2xl��e}���I�j���%����d|��Q,}���Gl�(�;"F���D*&v|�f��vQɭ�붗�P^O�Z��8����hj��wi��dǉ/1�}#��~Vu��a6�:�l�g�� �`����8t�t
\,�7�(�4hO�"2�`9��c
����.{�mzx���"]�r�)Po>a�>55�M���WKZ�]�c+����[}�E����	.73�rš5�̉�?��i0��]���}��S��Y�7�ިɯ��r���BQ�A�c,,�{�GO���2SN��W�����d,�?S�+.�T���U��K�V�!��>��]��~��R��&��H�\kưz����/�7�5���k��M9�<�8�J����.\�H`��
n�("��-���~{�2I�c��:���i�dm�R>�h��42ow<py4���c���Ȏ�E����#W���OqX�(Sۼ:��l6T�=�ή�`��Z[KX<*_�V���x���<նK{!x�d�¥��E]	4��zAm���L��x*b�\}���;�;yќ��4C�`Vl�G��6;���1ϊ#����h����*�c[���Fq��U�C`�r�k���0-�l  ���z�pA�"9�S��w��,�U\�F��ab�4�'���S���߁Nv��|�\�s�QWM?�����/O�8�7��sK��TW]ᴼ���١���w-�)����	G���G�w�s^��g��O z��!D���B9o�5��;5�i��pICe�U�'��s��D����.r ����\1��?	g�dr� v�\�/B ���aH{��k�ȼx�x,L�ϗ*���A�
�^��@�[K�fL� �M�|- O5��P��<k
�lԻ�8���γʹ��GP�7����f}Vø������IΖR�&E�D+��\�@�[ �!E���c���[n�QB��.;�*c-�O�{�[�F@e�;����&`�W�6��D�_h�Rsg1$_2ղZ1����h?(+b7R��̗Pd�f܁��_xW�<GA:q�SM�9�d����pXv:�w�|&�Ѝ���щ%ubwݖ��Xy���'S5WHh��݌�x
�N���}����e�Z���R��Q&{la;��5��T��/sN�{-�@6=�y2��s5�b�Bܴ ����4B
=#ٲ�Gj�»a�s�.�Q�%K���٭�����7 �ɉ�M	��X/����������g������*&]�����Ʃ�j\�X�Ҳy1&!�:�~��>$�z�.c7ǔ�!І���j�P�٢۲@�x�|�K��k �g�:�K��`���|��ܣ�e	*�s�K��R�xo��7=�����X�/v�X:(TEv�o��(K��5�6 �yrB(�b
ډ�k4=��`o����%��d�V�[��;��Qo��`O��&3�fq�H�ҮMBU�$��Ĥt̛;.
�-h	B�g��R*q[i~*�Yv4��H����=��Ȣ���4��@�F�ņ��%a�����M���qb����0�	A�㟘�IG�+�RE�b�x;hؿ�1�: ��ޥ/?�lq����q�;M�(�QZ]
e�NZ����4e���~1����G������L�U�e��=}����s��8d���<{��g��:������W�&^��UO-0o8��6]��Z[
���VlC]�(=��X-JFdn�^�!*���P���G��ǜ�mv�\�i�3��#8ܖ��bVp:Z�*�ZGO�Z� ��Ւ�6iPq�Ŵ'�FǼ3X���5%��qr�@j�ר��?4��bUv�NCHF-�!34p�`F��
�Te���a�X6�COEE~9���9�r������ߣһ�����ָ�=��O�I}�QJM�,��F�ͳc�ȉ�O�r�SE��Ks�lk�W�|�R�i�4ض���^f6��� _�A�� B-|��ǀ6�js��h��{�س54��C� ��>ME���;h�v��3ŷ����7�8���)>�1�T� �����cÌ&q�E�
�a�y���=�	*]!LH��Նp��#ʌ���2���!O��?MHB7T�7}���ƽS��) ���ϲިO^�~nʠ�!-�$wO��x���B�G�趼Έ�dfq�����q����~Q?	E ���2��u�*cX
�lc5�� _�4��.w�]�x]{+�i-#ԉ��'P<��Rn?3?��hŒS���x-����沏�7�d�p�r�ĩ��a�i�E켖2q2lҠϦ��1b��:-�|��}���ɂ��a���V�W��seF�XG����mk*s����{ta���!��~��7�sn���b	�Zvzak7���Y�V櫩:�����`J�b�?,�,���>J�'�.��!,�D��l1�Fd���"O���Xu�P7Sŉ�������/� Je�'Aa'���?05s�~��鶠��Ҽs��(Ƥ��'q��`�����#Βf��.ɑ��K8	�R��1%�l�T#�o������R/��7�2��Ua"N��ҿ��;k��?����C'U�:uv�a�OT�	��n TM�$��W:^�A2��%Ё��0͔��P%�>�UV�n�9�"�e?�hS��~��*5��kcԐ�=�'* ��ywq�Ҭv1ri,|2����?rd�pч,(�;��/���/I�^��� �N�0{������۳G����� p:��`��/� ۢZ8�M����3�Qv�kx��HK���e_���&�bA�K��b��j&%uE�M�q@+ ���Iaq8�9�"9=�2X����J˺=�^t�̼z�D�̩T]bѳ��� #rb�����PRD_�{��j�������eW'�
D���Uv^'��ɉ��E��}��Ɖӓ�����<���3�9��w�/�Z���|�V������K�K�'�]2�\���*�����VԘrF�=m>�Tl��2`Y��>o����ÙT#M��=S=<ڡ�ZR�/���vݵh�Xz�^xn���5
/�'d�>2�i��dI����M
eZ*����G�	Y,zx1�5������C��!�-+�
�
�.���O�1�Ɍ����.�_.��7`K@��;�#�sR�1;2t�7Q�X��z5�1�"%w+KEs�,�`������"�l�v�%ɛR�N�*� ���
뙕M�>/SA�}#����F�x��S��s>[{��TW�`�J>��AF�,�5&e%��>a>��|MMh�\�фeI�ʨ�=��3x>�Vb��0W�nHC#)���H�YN���-�{E��g�*�~�6߾S�5�
���N�gT���E) v1$ϼg7E;HD�R��4���T5i�O+�.����� ���|�e��s�n�e�ݎ�G�'��#{���Dtf��~�S �]$�}f�3�{t�h/�H'3�#�t�4Ε���ȁ��O+<�i\bkT���qP�Rֈ+���5ke\�X�q27y2R��z
D<�T�����+���l`�И���m;��������H��c3�I��Q��whV���Q?�7@�ad�0E�j����;y��Нn�=�O�+�UO�	ӆ��/���?z0~A2��9:�;�x4�Ո��3�6�Nh,�U���*�tۚ'bD������GX�����uO�-��Y�l8-�ĺZ�&nX�S�t�w~�pᇖ?3i��P�������9�%����LN��4rC�N���</yv�xº?@cO�H��"�}{2�����T��3��x37� ��{#s��SD}��»$��7�t3��Lq�- ��i63��_�������N4�#(8��z8)t���jy��u��sy��MD�@!l�����B0d	uGc��+�/ � 2��Kdy
9�[��C���'B$$�j�^g��`�Hl�ߕ%	,���YM�);���垂�7�
+���+0�|�ͤ~���� :�E.f�"���~�jY�#��Y�g0f�
r�2F��
R���ծU��d5���Ń�����ڝ��V�*����*I��s�;8`�i���α6聭xQ2�]�q-�ǎ̙��h�_���[2��A�*Y��W{0�! �'�{
�Ē�hp���4J��J�&p�;8��f�s����y?�щֻ�s�5 g�W�%�R��q_����<���#+�z��8𙷯�!$h��ǐ��a V��d2�m�K��RLB�/��Ѹ��EP>��X^���F���ɼ�
�.Վ��.�<��i�X�Y���}�L.ե;!o����n����*�禎�o��h92�o�x�X,��mi�B�����;����:�o�~-]wKIc����X3�ķ��:�L�֘q1E���d�^��뤙���Q�js7~��nF��/N��P<5'I�d7vA��gA�d�VD��&�J�B�%�M�B����C�R��/��@ש]�[�E��k����
4�U���K�ʩ������C��i�{X�_#-R��eo�������j���4�)�Pm%ú��^f�{���H~q�ȧ�:����>��Se����� �H��Oݶ��C}�]U�|�q��^3�6�8�>3b��TDcn�CfEقk�X7�VY�Qsбm.�%�r ��Y(�5Wߠ�4E�;.5�5���/��q��_%��Z�@�b�o�0Y��Q��v�j�8�o=}v��m�V��԰�Eh�*���s�ś�`���.j�o�<v��>ya���=�KOT:g>�1�+g�jR�ax��Z���1bcf�v�!֋u�U���X�s�v(g�g�*g�G��k^���e�	�Z��30��I��C)�Şv���ĝ�/��(���2z����ĚZ��va�eg�0�؜������,	y�"Mа�ֿ��/=m��e�l�}��[
A��M���b��ǈy�e\�mJ�aC��ߙ���@o�G��(컶�5������t�+�uM#cc����L��2��ӑ˫�Sos���B�ck��|0T���IQ�
Z�Ǩ�g�}���w.`�Z�-�:�z7d�Ŷ����nR�����0�L�\	{e~k����]��䴥Oܙ�?S3��#��pKbcǂ��Sf!`@��.enS��yR8Z��b�Yk@Xsʸ!Sme��l��æji.Zj,�<~��A� ��y)�����a��VYb��� �PR�Q�"�ސZ�����u���ʉ�?g�Eej����O����i_�����9�溏.<��a�����>�����ňC���e�뚳(m���) _��̉K����S���^��,K
;gX��Ĕ1��!eI�S6[�!��y�ߵ���w�т<�����
�b'`C�����H�Y驟�M�Ci��$Q-W�G<e����B��PO�Am�V$kHfbn����nq�KO�����r.{o�I��ц�7� ��ŋ�\��q\W�{�e�Q?Ҝe	4ɮ��Ψ�����@��iTs�b��%���:����|��s5�em��)��97�NdD�Wf�A�`��=�"VPp*��N��	j��%]��ݞ�J�w������!���}�@�����B�`[���WpS��Q���$��~�@ ��mf����9��z��a6�����?�p\$�hm ��ey��9��Z��02C��������d"3#M���:���ơ�������-����q~�� j�TX3�u�S������s�R��U@Z�:�
�iu�����~>����V�w���<�{�@'C�9k�P�5����IC/bD=��{}���<�q�����A����
n$p�j��c+Y��/%2�?��v�VP("���ķ4M䲰���S�dS�:�#�U�	�-PX5NDKO�����D�.���?Y+�ژhO�W�!X70�-���=����Tf9�M�
�0G��S�ȅ)��i}��"�셡����M3���C���R��ܳS�u
����P]�4'�mw����{N�J:����aQ,�G�oߥP����P�����|\UV��!����ug�G0�c�W�$ً�JQ���r���=i��(�Y�������E=���qP2����JE:Pb��h�ȷ>+%�6�����gu)c�11 �2�L�j*����I���vé�״$�ᔢH�'�	nC��(2י/!��yځx����� �A��N�5ңdsSd��\�@���2�_[}��^+z�o+MH)c�ȟ��gb�OWm#(33��hr��,�O�!��f�{��y�����7�bu��u�֓�.�5�
��Y�ܢ XOU�{��+��{���'m��#�������Iґ�G�B�u������;�$t����Vn��I��L��s�a�]sJ�<̐ED�?E��h�"�T�ntj���TLU��IC����5ߒ��G��%yvFi�d�/�¹�?m�՗��=�̉=?���a!��qyL�	`sPsi�
ΕQz< ��
�G�$��O�EB��܆���f�{�>6�`���d��|ڧ�EQ�O�9�ڃ!���/JÙy�Q��̷S��rA+(8�����J����wVS��aOuF�mfvo�ZQ�>D\ ��K{��FY��T��K3�H��:��Q�,s�PW�04p*]'�����:+����#����o{�_���9.L�:u����٥^a,*�2�� �Y��o���{��9Ff�.zJ�w%/�X�1�mǭZW�T� 2����	I�j���>�B�M�TQ6}��2N�&I�$=��;�����l:��IQ����!����>��T���A��(_i��vt�	� z
�K�((�����1�������G���?$ޅ��;f?E�a6Bg���/���&�_&��Ea��a�Hē��U���ɱ�ܣp�6������a��ΨQ�!�|J �@yQ{������Y7�<�["3�01LR���u�|���G�<�Ɏc���륞�@lK���P�D�,1W��4}9��y���R�St��X��Ƙ��Lh=�s58�L@�]�2�g�%4z���e�Ĳ\��W:�l�����o��ջ���OP���*Ar�����l@�_�a��d�U�X;�8-���-��,A����٫��g"�`��~�,�WK��z�,�V���7բ��I~�9<_G�)������>���ǽs�,'V-�Q�B�	%tI��n�q2z- �������Fo��.,�
3I�Nw·OW�9��c^L�����$��pq�R�[��$a������QwN[�C��Ǭ�Dj��F!��̻�F?\�t��>����'G�-���_t��x�9<2
��g�i�~p{��ї+��5�-��/��������,6-7��}�0���ҷ�OK,�V��Đ��\5ßex����ぞ��>M.	�=7��t����|{by��1O�.�s�W�p��#@4�T������dS�2��t�RS�(�1t|��ө]���e�¾��y�(=�ޗD;�ۅ�N����Çf%d��Y�&��/���������]�%��4�\��8�ے�fXz5��3Y�ˡ\���,��a���3_��.<�4��Hk�W��[ƴ�l��v�����|��r3ؿ��������@z�	�#WxP�E\R<N����t~{%�G��`Y��a*	da=c�/V��r�SA
��&�/�,�SꁸDU���`CMף!�w0�N>�����d
�[���̃*�[�ǅ��J�a�����D��^��/�Ț�礢Z��.�(�E0�p�@k��*`��:���^F)Tc��s�
����yX�L�O�>G�^-d�G�=]�[�N�NG6O*����w>�@�`I����bO}��<�#h�+���G4a� ��,���li�K�-4:&���-z%�/�S�<~������bfM	.o@R�2���yf���s�/���rM�o�֙�̋���d:�r	%A��W�OFd���1�v���6?`�AJ4���`
��T	b�I���V ������ �ӞC�!�O ������c	�	�l�G|o���5�)Q��Lw�r�5�h�	�"FD��%��7��q�|Al�V���0^Ϻ��*�x��A+�	���ëɆT`�އ�n�W�%=�\в^Q慛��F!NpjOf"�g� ��� |�z�p�p=���TrH��lC<�ԙ�X�wB~D�f�ę�xf��i
?_�K<h���i���p�E�Q}�p�`�Ǧ� ��JX�0��R6*����w1>@v��=1Ɔ�i��|����1~ۆ�l�ٝ�r�I����%�}]E�`d悍��f�b��1��p���y?�� Y�=����Vg�1� ��B�wĘd��զ���%�`�3�KP���h�vns'�ie!���x,޿�F�6 ��naL�
�^�N*��݃���������_� ��O�d%��̣�}Pfm�h_��
>b�Y��;�٪�%	<�1�2�P�r)�T�h�e^�U݉��.�3�y�Ъ ��:�ϯ����ͅ�D�DvsV\�o�����>�$D��������%�fcDra�ao�������]����*ΔR>	cW�~I��4ˇ5����B*+�B+H�����Aa��7��rs6������_����2�^�C3Z�K_-�EB�v�u]j٠7��T|DO����G��2����e*��#����đ>s��Y��m�R��o����{�fg�nݓT�d0C̱���h����uJ��фG< b(��d�L/	�e�Θ�QK#̨�yNՓV!�Z�^t{�\I�B�����H��jC�x�ë�N��tc��KH���w	VqG�af�ܸ+o�Č	Ȩ�յ�7�)ʬ��V���U^֦����R5cG�fp2�$���<��L���M��yO�/�g�z�ٚ[C凉=��f�0x���<���d�۾�ۃ
��M���z���'hH2���=y�ǹ��:�����Y����΁�B"�;r`t�(���/w0��@��G�gO�L5yj�g��b%1.�|G�)e?�m� ;>�_|���e W���w��	6@ַ�oKw>����4���e���� ��[R�US�V�=��j�v*	~�k�ޚar�Sm�j�_�����ňd=�(Q�;���'f�I�3Fey�u�ӚO*U�W&�mt��%�+��pڍ�Ą ��q�|��ve���������<�����s�1 ��P�ĺ��[?�"S�ܳ�vw����Y����H}�ߡ�J���rC����ģ*Љ�� �0Xz\���_<��4ą,�#��8�{w�'.�௓D3]=v0謞�[�T�-��q�fUNŪ1�B�W���O�!��p� *
�N��ֆ���׸�W��6\����nsq�D˕#�6��""z���m_*KNn���1�8��+ǈV奸q��)v�9��F��Ȝ�T���O<\Fƙ���Ʌt��8��g��x��e	Y��{OL&U	t9U�Z�����qLze���	�����5)z;���t�����'�+�y=��`ן�^G���_���Sv#��%�%u����ۥbFF��E����eSP4�(���ɈI�{"�.�в
	�����v�7\�B��o'vS�G�&{��5�)y���Iؑ @e\��lFR���y�\�4N� ���i���B*{�y� �A�8�Y��w�.��q����+yP����1���'�Z��ZB�2\��(T��J�a,:�%��  �z���3�'>� ��<t�o�7|�7ElF�V�=ch�A�F?�h�畅Qu,�*���9�3=�.�t倚J �Cc�^��D�!*eDk�������P�C�3��ؚ�������G���F3���?\0�<3ݱ-t!+@Z��現Ձ�c<��s�ݍ	���'�"��@��:��m���ݘk��<cJU\g�	�|�+����Pœ\�1�[%�@U�62���B�ik�N�ɲ�0ft]�
��M���؆��zQ��m�w]Eز�.1	hѾm�@� �@!��,Z{��.�b쭳�ӿZ�M�x��q*��?�D^��Y"�!���rg�\�U��N�N�#Ҋ���z��++ڮŜt�����p'G:�FHk�hSN_����P�I�1���J�S�"md4F�����q��w���*E��3aТ �xG6
;�!���v��LB�3n�pz��h������u������H���صP%����h�-��`2wt�u�\Vj�/�Wa�c4<C(F���'���l#�cp�h����o? Kٶ��%ϔS9�q���]�.Ь,�#�HE����(@'tr�� ��Dـ`<�+B8*�Č�5M�t�X���ld �M��d�c�ˑ��<(�baҙŀv�+o&I\G̍h(� �ȱ������+rw�k]n-�����4'7g�茣�[I��v��Ի���D�,����[�g@��$�����$;@Y4A��_E1q���V���2@��ݷ�^X(��9}�r��R�|R�����l���j�G���3�,Т������1���t0[�{LAF�6�+����!�]X���G5Ky���iH!�n�C�{G(��M��ۍ�p/�~�o�^{�H\�	�q�8�gg@��D�!nE��L�P0����C��1���{��і%L��T���a��H�u�'% ?�Z0Ǒst^�AH�,W>��l�<����%�P�!�β� T��o����S�����0[*r��!� �	��;��0��\]e��k����3��}!��V����;�CcB#��wW�J��"��=Y4�B�
�=+K��z����ׯ��'91A�
+ԣ� ҙ�۠X1ǫ�7��4�@���R�W�u��~���j%���[��כn]�b�<}��gw�;��?Q�T�0�ncTCΧ�P�S(�b����!�ڸ�=Ze����뾋�$�ʫ���tQ�f�>W�;콈�r��y�y�ʷ�Ev�t�W�۾x뺟�~5%�Y�p9JW�v=9}�˺���%����2-D�%�ZI�R�i�O��V��7��9�	���G��"А�\��2њ�J�9�+X�Go����)�(HX-Hȕ��S����!G�L�,���j���\�s��>7-+`��X��-[�HyPX�T8~�f���'��u�g3�l�0|D��&������&S�i�X&�	v��
?�X� HV�N�ĉr�	ֈ��A��"���Гby}�����;ϛ�X��^&V�8G�F��4�ʂMm/��"��l��Ɵ�a`m���(ѐjب�h�n���� ����M<0��ݲ���KؑT�X�:[^���=��A�)�A{�u���_��-J
��n��ΆǺ stM�+4�s+|�9-��ɀ2��#���L/i�c������P��'rx�����y�x�{{g��~-�RV9:WY���P�xR�X.w�g�U� �g�h�^~%^��h&���8�{�IJi�f��(L��׳2N��o��V-��h�)xz]�ٓZ7���]a;X;w����ӑ ߽J+�9�R�3W�A�qj�]F(�Й}6+�c��Gf{��6��Og��iY鷲��׀�5��!��N���0�a��pҀ"��#�3&��xi<Eq����;�.J�'�t�z����2i>P;cP� :l���Y��/5�dٻ���qG�1�x��lo��)r��x���=��o $dhm!Nǹߑ���C����!��j!�8W4�>�\f������3�h��E�Y[���¤�]:(���@�T'�!YE�1���P�i$F�^{�R�­	1��nOܛ�A8�>T�y��!i��xJ}��>�y��3�B\�yi{�Ɓ�>����Uv͔[-���t�fǣ�,������)���L
^��"����V�����WjRDv�֐'����x:]����N:tA��P�va� ����-���c�����08�͟�c:�;v] ���Y���y�Kv��Ϗ��յ�
pp���s�����V���i�LjK=nfILT ����h) �$>�)#עv0�Uq~�(Q�QČ�z��Ɠ��ͯ�w=(��p�OL߾˕v�;X���ѝ�_��a2��wt~����Me���f6k�͝�c���Z���(Z��'��
o��I�v}&�C��n�9@6���G@�@귞�U���CH���O���D�w�R�����|��ќ~���v���Ҟ/�x-���U�~ǘ�����)�q�4N4+vF�aAw;&	Z���J��� �Hok�R�N7�rGbW{΁�t��n??�_Mji(�msIA)V?���������a�[BG}�t9a瑺ڐ��dWE���ժ`�l�3^o�H0.ɶ�q'�S׹�%�k~˿�$�����oȭk�8ٸ.6=?�����se`m���MR�u�k�z��e��f������]0�@L�)��T,��僼n�8�����~�`��{~U��ێDG��%}Q�:Z(�uN��L�~��������vl�4η��aNEu�ˋEbTR''�w�.�y��;9-��%'{x3
� �ҳ�1i�i�B�>����f2�!���AX�0ϊ\��%̰��q�8{U�%�j�>�<N�b�.M:٠��ӼQZ����y��TF[��DM�⦂xV�D���g��<P�
؃�/�ؒt���/��B\Ia�EU���L��2��y�PM���sY��ww��E�<�C��*.�H[��v���Na	�p͓��h��"d�����s��~|�wkL�)�aOh����d���m�{��-�Mi�>����$�a!z�EB��?�QmF�2��Ŀ�8g��E����M��/��U@��W����`��Sm�����Ͽ�76������z�i���%;���Z"��s��a�[:R!�{v����:���"�/��uNj$j�|��Y�-�gtr1�"V��Ȁ�L:�R�/���O�t�]$�����n	������l�}>ҋhd �q���B�#�.Ǟ�8�Ž�銆�H�Ke׷*Hc_��e������"/�	n �Wj.�����!{,rIaۂ4�Z}
�M��w�S�Aq��{�V�&t�F�uk\Y!|�T�́L��]i��{B�:뉑�\�LB���|Z�HC�$3��p�P� M�U�$�(Th�F���NG��S��j��n��'��B~�K�7Xy�e�#?�'s)�"�nf�R��2*��*ɐ[m@2g+xC��߿�M�5>,t��j����ӗ����p���mt&�'T�8Q@u:Ω{�&�B��˄:	���0��0�a-��;].����
D��<�1cqo�%�&�M���^yl!�{䒄�8�A����#��I-2
��m0���B��ٻ��wos|Иr��w���b��=`B�������l�K9BC�tbo�oԢ��EĊ\>DG���w�bع+1; �]8��ʌ��t9����^`���vA*=�XlK���c�Yl����v�7�k@�˝�w���H���_ ;T���H��vR�!"܊tm���
o�_H���9�|�b���C��3=�(uq�YA9��(y��s����9OX�&����ϔ�u��3ъ=BZ�4�����6
��!
}�_;��}��`�r��c'��{f!,�<ի~�o�O�ũ�ټS�+�
�vdT��+�q��̣|
"e�j�Ao�>�͡q�>o�:��(T�3�e0�����n��vl3���Ze��F&�7K�"�r�dj���
�{s���n��7X}�������� ��W��4����I���C�ǋ�q�������#�w\NZy��K�Mc�(����d�d/FfF���d�6�qk��W6��]_#·kQ�i���Nx]���K�$���x�V��:��`�D@�� �6��98N�\���G�.1��9�Z�^�?T;pnj|%���_��:{�L���\R�+�z��	�����ءBO���xT�;gZ*O{�#o���9F#0�#d�����Br�������s||^=�҅�[�g���/��T!��$���C���d@`�s�6�Wr[�$D��s��e���v;�V��? ^���A��N�Z$IVMB�o�]�Di-{����b�S�D�P�����Qu�kj���yJ�z�$AXBb�W�����Kq�|sn=�� cAM\�g��i.�?pd�Z����fyd�h��g&t�5�Xr��4/ArWXRrD���zD���Cܩ����=�qV�Ev��y�Kc��%�����&��wF�I�n���}��	wZ��<CX�O���{u�C��*ZJ���}���\B{K�D<mNQ�e�̌��@�z42�?�99�.u�
f��Cv��+ǎhˣPb��t�{�C��4�C4ʿ?�����=��9W)��<X�o�5��"aP.��b����<��L�D
������a_��|�9�cw�-P��a�c�2�g�wJ`St��ywǃ*�
����m$�";����/ i�Ì�Q��l$}����n��,\����M�`@r+�5g:����	}��y�h"���4������H���:�
�a	 �c^�3mK��BC���ߪD��ƆjIA �B$�k�F�"ɚl�0�KbN�D���Q{Hkߞ_�I����⟁?0��ύ1�)��7��\���pr�@螮(у�H���9��ASc�%@�ߩ{��m������!E��W6$�N�5a�(���8�pv��#���3�Qo���R��a���PED�c:���`bt~j�5�yv~Ri��Q�Z�n+V����@0!��[���C�S)�HK
�qo)����q��8~�)U)1a�PX��&�'�. �
�I=��e��e�ҴyֵUy����q�I�k����}lY�}��ъ�C��Dr��V�CJ�/�5)�#Ot�a�-`�l#Lu�
�}�����EN���m�<+7h��{+ⴎ܏lﱶe�
���(��"i�t�@�,�]B��m�:I���vB�!�� R>eE9.����V����Д���)؇�L���^|������e����C 4�d�L�F��t�t�:YQ�%�r��{��l��ol�<�G�f����w+Q�|�,<�9`\�=&���WE0�f:�t1k�m��*]��;�_�>�QM_|�i6
xt�cl-2��0m_{�;\�T<�:S"��pg�9k��Iɍ��f��!��jB�:����~;�!�|�{���H7F��Jh��&μɋ�mp�z�Aq��H1�}���[��Mv��_��cL��oh8N-#�6Z����ŬV���=���i�f ޜ7��3C%��w��G'�;�cQ"k�3P����(�Y)��֭ݶ�*J�T��xƈ�_�@���|�]����&`�޻2����������֢�ԠquI$h��G�V1p��~>D��al#lK��yUI���/���?7�r�nrU��kJ���m�ӌ�cŰoϪdv�I�>�,�H�1K��IZ6PWB��t�!.�ق\e��y�������h%l���w�|����S�XF(��c�V��65��Է4L�C�?�/�=z
�h�z{�\��u2�cm%��E֏���
��'�'(V+~��-�Q����%�{'�i%k���"~�&Dخ������*3���.o��l�����U8)�Ej+Y�F/�(?��T{�?����L���Q�� <q���9����sa&2��o8�B0�ȯ���y����g�"\�yQ�>�asA�Yn{�u�
�o��jg��(�ݝ�����& ��^s�����b;�&r�͔���ؖq�FT�K$��"�������J�+.�}ƴ-´"�����4B�w\�;�n�)��!l($�v@�2{�|.�О�eX�
B�C�ˇ�����G�T��}��sU��Ў!��_�ΚE�E ��{ :�?�	����`A�;U0Pj��mo,ֹ5v_9���-�Ȗʲ�	|�T7�QS�6�	g_B�0
YX���}��j�dQ>�iAB%����p]�\�+���$Ȇo�/����0�B��$�A��>�>_G��e��]W�'�ʱ4�4$]Z�������P2�����ŷ�섏%9�j��j���i�s�~_x\��U���r�S��Yu���"�TTj"�c�7j�	�AL"�[:i9�G�1��95��D|�=[���}�� s3*ѿ���'_�p-��f,�%���ǫ���i{��F��4�'_\��F{����������4���#�	Y������v��<�����t�����կ��ZHMu�G��d��3����Wn%i��t1�zy<;��HҀM�Xx+t��gW���Kٰ�E� �֙xbҠ��шX��@%�;�t��&����r�d�H��6&b ���œ�U���O���<:����V0@.�3�Ơ���r8����Ʊ±EE�C��o�����룳�m�$��������p3ۦ��rX_�۞��q��@�	�֝�WJˏP����)/��ӡ`S�h��:�9���_#*=	��s*¬���D�b�	����~�mz4�Ao�����&���R�^"�ҵ���5�v�?ms�R�u� '�¾YIM�~�܇C�?�C=7�/��6�{�@t:�$l���o2���o,�j��h�� �/Vd�$ƶ��DO��ώo��j��7��}Eн��f�iEG\�@?�5�o���"��¿�MN=Au=��av�[��?�(H��t�bι_�u����xZ�*��^�mA�:�oF�-�7
��E�,���h��u������P���ik���a�u ���+����4F*�ӄ�P%D���͓�ob
��^�s~i�m�$�J�5}�n�����W�1��=��ߜ��화�)"$O�v�{]�/����~�*�q� %|�J�Ja_JA�&͘\a�a
�u�3^	&��?�p0�>X[�}�Ol�Boဉ%TA���ض�q6P[����_}��c�2H�@.��e%Y�� ����	���s��yRc�˶�pUsj���Y��{�C�Ks�<�8��υ�#�i�$��֜Tu/w����d���'�Aa��b���ׇ�O0�QH�m*�����O��?��=/��u��	Ϛ�7��wͲܚ*�ҢD�F�Yd���9^�%^����ɋ!܈�����[H�j��Sf^-	W�/�쇠�B��R3�^0�컃.�
%l:���(���yog5Q�찦�ieD1*U��	D��*J���B�&��Ö��e��҉;��C*G'l]��e��al�M�r�b�<k��O=` ㆊ ��>B�6�����`&���щa'��7��z�C;�)y�k<BY`v��z+$>Z�����?�4�3�[��t�J�k���KXcV1�u5,�2s ���ӯ���5��\�|B�W#�t��|�-��.n����?�������0�O6gۙ~��	���yr�q��̨
��wxZ��0��q-�h�~X�U^&�9��HP/^p�#�4����i���*�]^d)a�+۫�1��崵w�6zb$�Gz��Cz����7�d��ܛi2Q�Q��w����Ha�l�z������&{aY[Kƭ���L2���k�3`�����,�H
���Ѡ%�Ӳ�O�����Uy@�M�\R�a�c�8*̺�OS���Qh�o "ȑ�ڰ^�^�,.�~jP���.2z�����K�pp��<$#&�G�6!s-�d��(4q'H����u񻫋Y�Xb��`i��F��<�W��Aꉝ��tt!kǊn�k��Z?�/�~�b�E��1����DC?�8㙮�q'R�lH�*X���&�"#�?V�M�ڎ�F�H��d,�ae��
Ӈ�14��LF1*3xk˰$�+���nYm[����< �D��$�8��h�&�NW��r��9��� }*��jB��6��K-����m,���F�H,�uLx�Ǉ4G(s�����#C�"�>qT:�D�)6��� m��y�xߑ��%�x�-WR�(k��|�-Q��"#F�w7�%+6�3��gU����}�U,��1�V�����d��.�!���[?\Ψ�n;�e�J�F$P���N�iz}չTh��ؽ�<[�B���cVQ�|'��]�E�"��}���iaI�����Z�k�M\�W��w�׮(|�\T<��!��$Ms����I��l}xZ�g��z�F����9��5���w1�^O��p��/c�e`Eh�|~r�/����ki�6,��JF�QAz�z�l�Oÿq,%�rS���3��K��nE��:����Zs���W�M��E��(�N�l_�wa�Λ�h��:��s����cpظ�{��-����k��%UE�>j�'M�W��Si�߬�w�x힛���[���IL!���Q _�����3���^�L�'��q��@���/;?Y�wޥy��b��L"C��Nǣ�}��I�R�m�}M= �V�枪�ܼ���X<�? R�i�&A��E)�;��������jd1�0����*:�A��ƚE/���s5��J��}��f�{��$���n�p۹�JP�$��o#�T��F���ڎ���Oq՜���r�m��k�����@���v@J��Mb��HX��Q󱿹�� ���J.�hEE��_���M !��u�:��`�{1wӫ�F5k?�M�wO\Z���*x��e�u'Jk�l0���F�n�mL���+�xAEѣ�&��I��s�m���"���'!�ϫ2��-8�}�riP��$��!��<I�'���N����i�#��ɪ�D�)�VC��+�w,xR�\Z��6��s'�=�J:%�ў��K�x7�����A������A�R���,��~[a��l�d�7c�g$\5��=��j`˧��x+-���~�k}���q�	��b�u�o����*Gw9�+��5��-H����Y��$�@�����ɿ&(`��:��J>H�E�+�n,�܇����Ym�"��f�ӧ�w��զ�h�)���4RQ���f�Y�� �0�<��O��ѢpQ�uY��\�<� �:��)Q��{_�M�> oI,���߳���ք6�3�Ȕ�v%O��9��b=�"5�����s*یV��Rj��4�=L [0�s���|�EX03E4)��y�ZDԴ:/�4w/�.���	�p�����?s� f������,�?Z��W��,�z%`m�� ��ner3*G�� �C�#�>|f��-� N���	�Q�@_,��Pz<�����&�!���'��Y�dѝE6)�ĵ�Ua�j ��{��� ����f��tC��)�%������y�����J!p8�$�a9�Z3������s<��ğ'+�M��~s�����Ԩ'Ja�M�S�z�3�c�!��\�Ix[����$���Fus��8v�js!�d�졯�k�tU�<�*�Cbxc�ӎ��-^��GhOٲ�E����t����j8��}��H ˍ����{����ޑއ�{�O�C���D?�P^�!����4�w-.�*�B��[��c��mh!SF^�Ȳ�ONҊ��v��k�æ�f�o,�kOWP���:�����o���d@<%XԵ}2����ft�*DෆJF�5���h��#a*t;ѭ�>&���|��-z��xrdmᢇ�Q�7��2�%A��!1W0J�[�L/�u�*��rK	�髠���0�HMmm@Ï��A��Jsd�0S�sO��Q��I��D�fn5���B����\y>Al5!�^�m~���������Jʐ6������r2@n����[EB@���i)��*!(����܌J��x[����d��y�\�k��y�o���/��������ND�mbJ�9_�8����B|0u��/+�'�~��S2��?��Q�.�e	l	*~�}�ֶЕgL�T|u�b4�wi�e�s@�Ǻ?�~�`B���V{����$\I���~=7�^b�z-bSɴ�k��R�<�.y����X�}�h��-=�~JV#���2F�#%���:�+t�=J�`���P���2ZN��E��Lw"V،=$����P�㮫�j�q��Hh;�Cc3S�ZÞ�L�/2"Hԇ�?dvo_qV.eee)O��&J"�O�#�t	,�K
�5eT�*�p@{�Cf�����o�m�~q������Az��kDw������3���ݳ�Qq�p�>D��QO@C������q	/\�/����wX݂"�=��Ir�4�uN���
�p��τ`*��I�22p�Z��Q��8S�٘���P��w7�8�I���_��Y�<�R>l���{4Lzc��K%����r|R]���!͢�v�GG��8� ��}YV����k�)	ա�xc� ?afnT>��؝"�)��oO4͇*����+.�<+X�~�K������P��*�1�����U��Lo/��b�
+C��'(�����������p\]��E��Q�Q`6���wiu��Lq���b&"�8��`�(e�s�;HE>��g���T+��DȨ�h�1R�����-x���Ģ�1�-�GZw>��@А�Ѽ�O�N	՟v7e��gl[�eD��x��2e�947����V;��
|�z�!-G�B�(Ep�^�{�e�N�<J]�u�2�����
vy8���Q!���H⾿ۺM�4����^ Z(�ZHԱp\��)��-�r�z��W�����ǩ�%Y�];�):����w2�uN���b�Ĺ��&k�jn}�ꑜ�n�෼!9�2�fD{��NF�vخt����J͹bH����U|�3
����<$':�dR!�Fj��kls��h[08�ɾ<lR
|+&�Y�V�����~&�\Z§_@ބ����E��\�ޭ��F]Z���=�R�I\���pm��;gZ��UUQ���/�oӽ��m�\����b����� ������|�z.��=����2�I}�{ޜ�L� Z�Sw��)����:��9r5��A�=y��r�t�A	s��iPw*��:vBXR�FM.]�bU�V�JߋWe����,N�09cQ��q��� �n �8e��K㶅˯�k��T�c�z�TBf���Q��Y��n�_#P݂���4�Xa�%0L2(9���;,"T����H
jda�����y/��G��}v���m�@�ٙ#�8��d��㨲�~t�N�.l���K�X7�e��e�|�X�/y�|F���ӏ�EΒ�:H�U���'ou��^�f��hz�Koӟ���*;=�m�[K��L�lcsi�ňAB�&�/�5�h��������9&
�'xRA�xpUV~� /�zM߂護��i��˱Z�Ή�^厫����%	*��j>3��W��?��F�	�w裴�x��b������t�	iqro�͹[�BFI?�>^O���sӡ�UN�G\&��4SN�o8A�a�S��R�e.���Cݩ�i ̚GP_�_`扈��H���Mg_�q<I3�t��K��IM�G��
r	�[*��K8�G��W�Gӗ_�8�� b<Z3��WSq;��k���	��9A���B�h����]��B:�䎎Ur��bx� ��sӔu� ��6��u�K|sfo�c]i>�����]n(mO��ܺg�y����a��a#��%3���r��݋~�e��Ȯs�.�k�mn	cT9H�O�}ի¥��Mz�?�6��2��L��I�q�M�1��B��$��DT�C�$��H����	�e���$=U����CF���
��	��ȩ��>	K��/�oC�KP����Ǆ��:*>�uc>�!�y^�2�����Q��g%V�$R�h�=	��g)��4/!�M4[�[���ħ�.R>�h����ڏe�v��z��0��#��_��U�r��-}�)VYT�S�:M%��M�{���ħ������SYBC�9���Btq�# �,�S7"G�D6=?��2`�{�3�.����?A8Qhm?*�Ujl�`*��4�Z��� ��R���[or��sB���ZA	T~r�E,��2�<[j_�E�l .�p����f͝D�4�&Z��4K�vb\��q�~�����_�4�=�o�en��xIf���i�#c]�2�c]u�e���s��b����� ;9��U4�<ʂ���B ���85�z7{�=O�� m�x����k���0m<j6�9��[κ�dT�O�^�vҖ:���^�86��C3����/E27E7�5%��E6��;W{�##��K��1$�6�:��}�����h���ʤ�^����jd���~����}��́�Eu[O�|���r_r�{Dމ�TJF���@+�QjTQ����UǢu�ζ���q��_M0�����z�/"7����q��B>#�
~���h��;�te���W�	wd��B�tv�G[:�x�u��Vt�|�L�ZK�}������ƺ�6��[x�n�$�_�������$��t&�/c4٢�Hd;Y��<��A��.�șUO�m��!��}@����P-�.��-)�J(�!�	�#����d͏��E%��ȏd�l��vkK�Fﳩ�V.VX�<&�1&"��w5'��,3v��2B$���E'Y���Oy'�ۻo�~�Y�/E>�'þ$U���ϱ;�'S���Bό�����[#;�Q��6��ȳ���_ڏ����u�]��wUG�Ĥ}1T�;R���.�__Ed����C&Qw�̠�OU�0��&�� q�����3+����7���L��n�{��]��p�F�4)�f>r={���'�`�N�\Ņ_)��D����M���� ���~Dq@��hjH^-ڇ��1�W��wȔ�ٿ
���G$���=��QR&��R�"�]���vu+���jWP
��c���f����2��_ɑF*7�ޮ��Tҹ�d��QU��Yb���YM�[Qu��c�Q r���lhu�/s5c�"�\�}�"%��G�x(�`=.��q��UV�lI��N�w�(��<(�qx��⳼�"�b���;^|�u*��!��N_p�棘���V�`י�����mӊ��0C��r.�!�r�p
���;��zq' H�h�"���~n(����#�:]^�.nC���l�Ufm�q�4Z�D�M�B'̉�)ֹF���/�q�{F�+�Ss$�g�� 5�-�M&j���؝�^��ô<r�!%6i���k�U|*�hȵ���)��Z��a�n��/�::6�id�W5o��*�R�W��	AwS*���5i$z���S�Jb�9v�A����~����ೖ/ϰ��
���-�d���g��!��KG��NR���u��i���1YK�_�+z��x�m�YpV�i�8��x�>Y0rb��8�`\�(��$a��6�|.{������W�0��>�S�ܡ�%�#��Dp�v�	�7qO5E:�BJ:N.�������*8cM�	���0�[�p��&H��������]F���`���w��P��N���Tv�1M%�%��y�ĥ?U��>�i�-$Hlp�E.��'�lUޘ��J�jW۩��+[wp�P��	Y��º+kF�E�(�p:E�)�oKe�k��<�N������#�D��=u�o����ÕPM��,�]Nő��z(�]n$�D����W�{�_q�5��ژ@*����s.�K��ձ���lH�)ös��<E���H����\%z_t�0w�r�
�r�oi���5���<�*oؙ2������HiYʱD��@K��|�f\��>҃7O��J�`��\DO(�Zn���v9,c�%�vU���O7e��[wdo�q�j>i�#�/Z4�����UH.���@��ξ^ɻ�U*$��`�����j
	$�A:c=�5isq�Z���Ȼ�M�;��f[^/F[���	Ύ qݲ�F�N����1���6s.��EEZdn����w��,���_&�+�F]a�*��O�tO7��S���a	JjL%QE|���1\�H~??�p+81�5�9�A�P7HaY�y}M�+�VK�7µ�0�=������c��2l�{}7
Q��Q�1��v��ݯ�}0��l�� ҳ�Q9���mv�%�?����(�b�d�6����	�q�6{~��' l�C,��媺���
���2X��d�?���萗��8����%��0�6I�FqQw�Je��M�䩏��a�P績�ة5��5y�H��홊��	?�~����
4^�O���bG�����u]n-�U���jv����N�q'���
hS�t�2m��.{�̀ΒC�@����ɺ�MA��u�v�ֳ������em���`M2F��7���i;?��ö���,bjbN�`�O(mh���7I�tΙR�`@�����|Kס����;1�-�[�ѭ�'7���C�a9���Q��a��%��̟��z$��ɻD;*�s���Rn;�!����D����H����"���#�(p��;Z��	`"�+� �{g�2�:�m�-�����_����sYF�8�r�j�b�S�c�&UbZ��?b4 �Ù���l��:Rϭ�:\�H����j��6��B��0l^O�j��n��o�w�Ԏ����f6� V�p.�����]`y��-��rv^��u�7�|���%;��3��n�@��!�$�:�=ҫ�"�Ko�Y���'� ���ɧ#�h��!b|-���lX����N�����PP��c��"(�il�E~�����^��������Ŗ���ɬ���\���}id냙�nl鄞 <���'�Xl��������6B"S�:_��q:�X�u���>�1�H�`�J��=A��w���r{�G��J��Ȧ�3�k�����rA���8�gN��N57��Ū���&ݙg��=K�Ƹ�e�a�/�� �#;�0[M���M�ʹ{�<��Z��Nxy �@ǄUFBe����p�޲sb��-�KWʼ��-���E�_CCSfS���t=���d�K�;d������^�����d�
�(�Z��>Ϧ9*o��y����Z�NF�r���]M�}rQjS�o�3C���	� .�1��GG�_90�B���)NŘ��������"�BLr?�o�@h��L�W`Ji�Hf�ٜ���:3�P���kc	���kqa��2��xs8�6�z��в�ܞr��g��Ks/�2�~��a�������){��<��Zu2��|Z��
��_;�/�-&��