��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x������jTe�)�D�b���A����1v16�|,J6l��)~�S� �B�`q���(]�s�ˠ%��L@��z^ߴ�E����\>lt܀��|��>Y-��=��v�r@@����Q��2��^ԭ>=h��^$��f]vY� $za��"O� X��R��ȿ�u��v��\@��
��^(9������U�M4�~�&om^���O�|�;��9J0����E�{pY��W��AHgI��o(�s�����SL<�9K�	���-R��_�l�gI��9M>�5��׎m�C����E��V�e�C�FU���n%{��
]�^
;{*�>Ԣ.Q����ǿ���_�#�q�ƞEE'+E��`�H��/d?���� 1)�|鏺����$�e����-`�x��E��K[
�Q��H��n�4���� �r?say�߅�&(�p��h���P�~��2
CQ
�3��R��^!R�Lt@:"� �N�Q��_����e8aN�N_��7���b6�����%����c�E�Ի�3N�����d,K�JeAND5\�[�ў�*.�c`�$�+h�����VW�"���m�ԃzީ��G~�3t�2a8S=+=�Ys�3���ĺ����W;#�܆�2��;�v�孾0^�@�=�����i��6�ؓs��q>o�����!��r�Ѥ8Fe���-�����9�0VR�=�a_�?{=1��`�2������\$��
&�]�g)�ݥ�(��	��	x�,�,��ai

~�i�vߊ�����sYUK]��`��ؿ�㳌�_�Ӂ��m��D4h��v��uFؖ���,��ԇ���0S��tW��$�4����[t�O��cYq$��Q<j>w	��z'�+H�1�gﮚL�P��]"�oeG�^��<�/�o�mǌ3!��n{K^Yա�no�l��8�� _h�Ң��o�v9���Ա��+@z�vhz���2-���������3OB7d�r��]��@(��g�)��N�.�I���8GN�,Z>�9_q�ټN=�T*�N� p#��(Fy
��Q������a*�R�����t��F0L�TM��r;�+yWPs&����i����,��KFP���ע�������{q�f�Ӕ��\�	������	Ɂ���-5ot.�esޗ�h_y���f���r��mސu�Q��L�Vd���U��y�d�Z:��q�b���"eԇ�[�G�>��?���]���%;�Z����Y��@.��m��h�Ȇ�;�M�����j�p(5{� [�ut�ߜ�����Ll���G����n�8�)��6��C��bE	��	QM!QyK�j�������*@�%G���G΂G
�"L��&'��5�c��@��5A��N�>:��8"��R�<���/��3�Þ:�*N�A�k��Cq���Ϯ3�2u�5e�t�􏚢r�p�ho�`�����hq�ܶ���c����'!���&(H�َv�_��m�)��/ĵ9���/[��z�����W4��%fΜ�n��rSM�A1pډ�7r�:��N�@*�+���U�-�����C76*U?�����m��'��U�\��S�L�^1WQ#>Iῡ>�z2p�Tt�EÛ�,x��&�����q6{���*]k�]2S���z��j��p	"�9ݛ#���P	K\q��oCM��㤄�[#��7��w5fV��)c%7S$F7�(G�t8�*w{%��+��UgFnf�C��	�ri'CY�OV'�,�I�,��do����B>Xk�Sj�m2 �D;Ԭ"H�{~A�p���'��]՗OŖ���f�i�J�-v��<4���bXN��r}
7�����:���c(���a1B2��HN�lQ�u.:��.��%1��z��B��\���i�� ��9�gG����A�w����X�����L�A֧Ǧzhթ��Q��欚`�`l �J�bI�<�E-6�s��{)Gj����zۺ��W�U[����c�|c���2,X0~�E�O �0�w�M�����Xt�$�ԡZ�&�㼡J 71�����N��"�����l��֏8?�C�h �/���nV�Y��t�Z�,�x�P�7���u�l���R<�������j�gEw5�� ���0�M��f������%嘤(F�`_�#�$l4�8��x�%?>�mA�r�b�����@�D�}��1��wE~�1�GDy��>��?�f��K��k& Q��X�7C|"�6��N$GZ{?�צ��V+�ځC�	#GLΆ�ʷs݃�`�>��l��m���,`����R	暵q�/��co.�Eo RA�R��]�a�	����`��l�%�6�v��nz����>2�ܼ-����Nk`�S�l�u�H��P=���t��n,�=?�u�B۳*�ݏ{�H�P�C=�@6{�ĥ7��.H8� ��<B���ى��%y�\�,�wB���W�\,Q�u��;k�ݯ{��W��� ��-���.j�̦J�@��{+VԉW��}n��!�A顧���Wv����p�����5E�RnB�[R�]�C���쐙��?eG�&� �B��Y�ZK[�J7�5C]��>�
D���I���g�*����Y�ɋ�>�%�Yr�ɇ����l�� �C�2�-z:E�Z����y����y%2U�q�r�
���G	�D͡�4�O�\տL�R6�\�^�.o��N0Zyê�Ϡ���3[�6hS���#:Nv�X0M?'�7�p�lg[Fr�.�h�Y!�����~��dU�Ǻ=jUM�ʴؠk&Ǔ�j�z�(�{o���U��W5���?<@*Wv��]׉��7�s�K�}�����SuA�P�|�g9Y/ʄ+�շ��\f�~��`F�=1�+}��>��j��%��+�p�m��=u�p��<L�qٴ<��v�JO,,��^5���֘,�P�����c�M���O�@_�y�zJ��峦��X�O�~��m$[6�y�6�1���c�a�u��	�d�O�O�<|�'<�ۅX��x�ƭ���_�|#��3%�>U&6F���~��SA�����H�ґ���@��KJB�	0_c�vi�Z(C���P�kX�': �Г��h����n�VQ�㭦��[b���b�/E쪨5%�����8�*���H�,�E�j��;ܲg�߾�S�Z�烑&ԙ[bPgS��P���H����Q��L�+�ʞ#;KTqYQ��g�,d��N�嚁��
��v{|��
�~��TYt�0]�I�����Ă�uq��5i��-=��3�G�T�o�����u���'��a$�.���&9���/�
�\km秆L�)a�7Zh��E],V���U������4�����]wN�CzHAٻk62C3ٺ��(2�nƯ��`|RЁ�����&�;!;��J�S�iB�-�Ě����Ë�S��p�%+IV����v���!"k;��1eM�߭�����U�1t��
���$D���y�$���+����q,?P�ަ�JG@2�"�-]�|F]�G����_�'�7Xp�*,���+�Ӝ  �)�,�WS`y�G玊Z �ڿ��Ɔ[���1�]i�kE�'a��p��;������Sv�g��.�x��6�s�l����C����}eV�� ]�yr �b��6�	�q=k$;%�ss���l�_�4��\	e��Q/ǣ�ʸ`?j�aP��+(�Y'C�GX���n�%�FU`q����,�[��}��kHl�)�`Fnl-SE7�N�f��j|	6˖�P�=
�bI@��?�&mјR�8WF2�;����F�Dqm�qՀ�SV!Ӱ�ǰ>� C���Yr��^:�j����;io>GW�)� ���\�ty$�>Z�4�.���?(�g ��g�x�]��s�iP4S����x5�����9��� )D����KY�k��ɾ�c�w����	@��MQ���cƎ��)6��O��rJe�6���ꭴ:�aӳ�zOZ#�&�89�!3�t빸!�rt��a.N��G�JB���Y�
Ҙ��q2�́�!�b�P��q��������Ͱ,���3�I|�+����o��ک�c�@7u�`���'M����J������l��{V�-W�묙�.�,�au�p��p!(0��#	C��o��*�&	e?ϫ	z��X�8���^阦w��=��d��&��a�'�UuX8H[���&�*�4�m�\3�,}W̉hq�
���~���9	X%��e.=�}h�O��9��IUULT�߶���x#��w��aAՑ�vC�Eڹ�%�%"��J�׫�1�*�/�˫�,������CZɱ�3�J� ��)�2��X:�/	�}hl\��+c�U�,`��j�v�4�����U!�6��KL��Ql"M�$���іY�o)27t�9�G��r&19�u7=
��,U�O�)��o��ny<-��(�d�'2����W']6��n���$�&��	�Vn����䍜�ۏ����JZ���q��!�b�
����e(��v�jjL�Rc3#�C@�<�,VD�u>�K���=Y<�4i>'u��jG޲;ʊ��=��nI��9�QY��Q7�T+���im�܁�*C �����$+�V7^���3�1Z[?�h9��1ӝ���
�O��z�s`�xo2��I�M���8��/��<n�1�4������m�ƛҋ{�qud�����K��K��R�����#ttm�l}���k�����)pX�P�#�,�yNJ��o4��fa���M�=.�����E�"u� ��#L����e/��>~�GC�������$<{j%V2����t:����5��z9�'��	��X���u冷h=~�"y�������W��=� �ܭ�֕���hӱ��h���.��P/ ~٘k�SFG�n܍`?9?���x{��[!I�ױX���#X�a_��
]1�0�Jg�7tR;Lf�ҎV�U�ώ/&%B�z��B��W��gmK1��rk�Xe��5�u�W怃2��لW�g�o]A��~ʄ����O�U�#y5�(ѝz�p?AP��c�Z���귉 c��l5Jc΍��.|��$����!���:y ��;�>����[�D�f�8`���ww
~k�TG��Nl�yS�R|�#��="Yl
mu�5
�}J�ψ�剱�4� F���c	��J٢2N@�5��f��}MK�!��R���BA����q�J�T�PU �v����>y�L�\������lL�	��M�L���!��i��Ճ٢�L��?0����(�"��	�:j�RG�D4�T��PQZe�}�*>�N[`�������E0���A6Qi�+މ�����=�~Uyg뙄�f1�^a�I�c�t�zu��&���f���[8�$0٥����_z�Z��O�tm�b���$�s3䱆�L#��t,s��� ?�q[�6�7S�y������ �0�������K�U�A;n�&��2%>lO���/'�T��II���ֵ�/"����l��,ec��ik]�iL�^t�&N!�Şp?���^!�Fኑ��Z{v6��1�2k/��C��[2фV��p$p���HIߟ��(h�5U���v�2{2�0�$�Fs❂�F�B����\LQI��ɱh�OD�*��&�h֭�����~�%k�
����H.R7�P9޺���O:2��_��
 #���
.ρ���ڳ���9�wυ8d��xǻ1�MG��9|ǉ�s# �4���Y��DY�Æ"��i�C�C]D�f�-_�-�x�i��%�A�Q���H��ʿ�\gn�B�>�u���f�i��$�17pX	(s��H��;�l��Y�[Z~vg�b�e{��#n��KԴ�����J#%6��4qKg��A�C8�=�(�^en`^�{�'��4��$�,�	��cL��tW0)�-'#�*�b�^�+Z��d/�K�cW���[*D�q+�}�J��Sv{V`pWzqB�YP���3��Ž��5@0��Ȃ0T��л(n�����#��u�� ���n>�䆵K���u[�$»k��zF	!�j8s)fP�8�2��tC�h)QA�� ���pո}7�ɼL3w���J/�X5u���߷�W/>1�i�ɔ5C��V���ϵ'��� 3@�!pq�����P�o��e%�<R��i����r�i4�S "�(��4���z���gR��1�N~	�,G�w�uf�`�\_�Y4��&/��v��h<G+��H4��s��O}(��P�T����q��&�M�^(��Qh�5 �x�L{i�&=.:�;}�%z�
:�i��Y�ѱeOL�'$x�"E�e!��Uxe��#H�5E�-%��s�����{�'x��^�� ��o=��9��t:�,$b�PU�;0��c���r&�p�'�7��6tP�\�y��<O�ǫP`�Y�:}�������ʵ����D���pI����5��VC�g��R�B>p^iמ"1�B	�>��.Bݹ���nx��ޙd�fq$�E�?Q���U�u3���\�!J��;ƿ6���:�Tn�Z�׍�_�J����jyҧ|�+�Q�L0��kIwyx�@"W�&��4��/�X�׼bZ��,W��-9j̢��0T|�o�7��
+y�2�p#I�P$�6���c�v$`��И�\e� ;�������u�Pev�Kc6�h�-�B��/e��V��6��uE���	1�ض��1P̺e�?S1h���Gz�A􈩡{�_�c��!�ǘf^7���LA�-pR@���Pt �E��w�i�[�*D
������D"OX���-�e^nf�Ė�<�G`�]R|���J\�NŚ��P�l�u���`��~&�0Qy�������掫o,j:O���C�:��VWa���G�x���-�k�pe�J�h!5�dg����'*�i:�a�/�`��|��o�]nḃn�k�c�0c(Xs�"�w�i��� @h�����W�[�:H�Z��������.?��4�3	w!].����Z	<���n�iw�VÌ�}�K�4E��ő��%!	(Wr�)��nJ�X���� A�6����;
�r�W�I��G��A?�Q4�%H��&4Sh�^E?����BL��_���b٥f�:ό�����U�f9�ك��������C��U�WEQ���h��N��F��I�>�Y�����l����}są�Y�ZC��Hޔ�C�[���ͧ�j�Ĭ����8"�6cM";�t� �% ������<��/��J�	�I�cQ��5�l8l<n9%�1���3�R���|B�gJ�Ou��:��㱸-���(�`Ĵ��2����L{�Ȯ�T��	�ylq�iC��ѕ�EQ([����j8v� $_����m�ڜ�S%)w_��E'O�F(��R��=o]�W�=�	��>�W��kxto�K��E`�����\ң�][�u�V<�&1�O�+�KOb���i��{+[�M�1�X���A�@��x���߻D��e�?��]�����qJ3�Nl@��YmR��s����µ�QCP���)`O���4|at#Q��w/�/v�e�YC����G��~a�[�B��AcA �Z�g�I�v�S�+H�`^n���@kQ.�ȃꄖ3��XtW���y0;9��d�	�<7YkW7=�؈ƫ�0o�?IڃX���Z��~��By�������nkr��ԁː��y�*��\
9⏚�9�%t�١W�3����Y�����2��M	m\�R��w���u�S���f$�u����{!J/��fx�����EN"٨�޺vU E��o��t,� ���s��o�j(���^K��w�&u&�:����vl|�o;P�_�Z�tK��S����}E�a����"E������Nc)u�$x��R^Vi��G�ۙ�>ʙ�Ӻ��Ź�T��w��^v���_t��O��ᕉ�,���ԱEUJ?�YO�3QZ��c�w8W[TO���3��A�-��w����V��#��_ [���iShȋ�hxD��	Q{i��B�D	}GQsUBHx���e���9I�>�����wp%��	7�-&���du�0
�Y&�p
u��+�9��FK*凸4��:����a�/���� �e�z�N��ڙ;�6tf�<C�\�rzj/�7Wa�9�S���{����.���oE����)Q���U�a�ߏarB#-��) y���=����UrcFV�j^��a�J��=����%�J��
x��s�B]ؿ�zV2��ُ��� *y�����On}"�練�D0�36B��[�n��?> &?bp��)A��XlX,���l�r��"�>�&��!�2���Ӈ r��c��P(Ӳr�C� ع��6u&EU���c��j�Z�|e����U���D?ң�:M|�%jE@Pp��V� T��L���^�B��hΙ����>��;x�1V.s���څ��5�����,�
:/��m�g�|*q�x8�vզt8۟���%��y��w�v��I��fh�u��)����F�y;�\�_�}ũ�2�������Bp���m���p2 ���jz��"�y���-��j��C��Qj?�Gڴ_9����u�=�R�=���'��R�4�+,n��Sй�뛔�}�����p����&������7�<�0)@]����?���Ņ�j1�^��7����;,{x�$�JG�� A=��+9Py����$7�*�b��/�й ���"�����8L�덢5���J�+�o���VoA�����L�Z//�a8o��t�SY!5y�`m>L�~�c��<�jCf�h��&���b������sce�4K�_35�1�;��kFZ�o{�����Fʕ��f)y����h,:l�����0a��j/�hXq�lh��t�6炚�$�����;�RY��i��Ԑ�g�e�i-h��^|,�[���{������p-����>�sMv�I�8o�W��+��"[�� �;l��U�����R��n[P.Qku|�0#ě��	Vw�ʓ1��G��G�(Gb�[u
g.�qHLAaM~o��0�$�"�N��tn��lg�;��JS�[u��U���>nY���h1x/�)8c3t�x�}�C����w�����@[����%N�i�T��L���?OM���/���,q㮤-}��z�$"Vļk�8C��;,�߶����&)�35C�
��(8g6��Q�h��7�ͻ�Uwޗ������E�I��Is�h5pD,cu���!R�?>�6"��טV�s�6"�r߈6ڹ�G�mL�%���k�6������9��|�1a�=�Z� (������[���MZF������u�D��=�M�Iv�c�u?_�=�"�(u8`˩�1�����k�H��/dzL)g�࠳i��И�ܿ�J"��koM��]�ӡ�\]R&dq���T�H�,�u�_�j��gm�Ӥ��g�ή�W[kp�2�NT�����'f^�R���ݰ<V��$}-�����#.a�o�I��$(Ҭ�Y��審@��#M�$)4��K7�E��{�;���.1׶�a�����3^����)F^?��k�
Ƣ
��D��O{�W�ܧ��:���M��Ǖ�th��b$K\����kF���R���Z=0����8�5�4=YH��	�yl�Ջ���v�`��Vɋ�ʵ<��О�ٻ0��|�xV�� <;�ȟ�J|1�de�?�;�<?�^�R�0�,�ٖ�$��e-�>���-��gM:�zJ���.�Y\O_���/�������x5�^�nő�*�aXQj��3����3�#}���6���ϞT7
\ɬ�w����[X��5�3��G���VԄ"ɎF�i�v����p �Z�u2<�
�>�R<��2[�26�����0���p��8��pdYnk�C���18�pd]�JSVp��ĉ$"�����h�h�l�g��~�&6,A�Zt�Ӯ�q�M-r��b�*����L�]2�����^�tEXi7�Y�'�ڈ���)İ?O�A{��6#6�􋡱A�;qO:yR��(�f�O�g�"�B��l��������r��D����\�j#t�!��'f9p��j�I5Q�����v��mc9���a�;�r8a+�"��K�F$+ooIie�Vt����[��v"�9G��
Pl�g��c�69�>,[�"�g�,>�W����%JOBΪd�E(wF��.�-�6sW�36ش����QN�ucw�h~M��W4�/D�h@}��z���a���筽���%��â��-c�J��(,��*%��Υ�E��k�ڠ!T�',��9���j�`��&`��f,YdQ�J^���ؠϭ�}{�W�m��U�^L�Q�)���l2u�k|�q��~R@%/�]I���8��n{��M�:���(���D�� 3��Ԣ�� �h���<�/���Թ~>3�t�,�ъ�^ﱞ����L񙅐$0��FI�8�%t��4�;�1�?�ꇳ[�:7�}a�V�m՚�Rg�� ��u,�#�?rAk~�c�C��?geTRpO\��?���z �d���[�y�W�D99����㘚�xG	[((Ǳ�;wX�~�.�P�
�H(*X�7�_�9e`2�H"�#�H��T9�(H��J}�:/q�?�V%� ��k"�d4I�n6N����N�ŏW8��-8���ǐ��-�̟�k�����Kl
4M~�)��(�iX��SC({��Vuϙ9����zč�x�h!^���_�"B.��8u-��J7�߱U�8���mX�K�
�≖K�*�)��uy	;R�1U<w>-Y��=�j?!6�D�]��&翸��\����>��lq���猌�C���<��g�zgM�6X�h��)����|�z��)��|�5i��	Ǉ�w	�,�X���vR�*�)�3;j*���q�_]��m��X��"�g�1� s�����͟����J��%��Ι������$ǀ�$�p?�%��ɸ�����G&?M�<�~���ͨ'�@��v�2�~�o�׻M���FL��$���(�#�*�|�u�J"rfiC���Br�aMW�:u�q�u�+�!r7��4��W�=������͒�,�<��x2Z�p�%V��4^���1��&`'�	-Oa��s��<��ЕǕ6�'�M4[O�<��n��BjR�ƵS��B��4� �m���	>�����r%U�����'$ ����CV�6?����Y���Cb��6_f�V�W��sx ��U�%!0ٴQg�rV����+ch��@�S��ya��f�ړ9�CF����=J��m�Q�&�V�V��J�6�+����{��c��'�ƙ�#OD��_��I��k@GX4��pÈ�dj����y�Т��<Yc���ͩ�S	�00ȣ?O�,�zHdϛe�b���� �N�m�# �?���	H�?�HDF�Ƥ��i���g�p�d%T���!�R��̘,(Ȉ�Z��>�qDbG	��M܂���.eԪ�)���X�ia]7T`7���]#��-�NO���Q�<GP����Z'�ضH{$I�! 8'#^���~����%B7p��i��CX�*�e�K�M�  ��}+�`Qs&Z`�E���܇d�9�� َ��c?���d�j��W4@��v$dY��
��~U�!�n���\��}$�t���;IW�#�X�:���9~o_Ǆ"���[';h�ĲO>�$|�E!I.[�i@�w]bP���A�pW_���A<F�s5g��-1(_Il��D��+�9�t����) ���Og<��n������:�:ه�a� �"ư�^��G��NZC�MҹՁ��s����\?Sf����Բ �<�/�C!��W(Uҝ"Q� �%!K_�ق�7�J�1�ި"���b���9����#��g�x�T��۠��X�Ai��O�F���1�аԖixۻ��Ϯ�A�¿r����C�䡤HqU�a�3F�q�ӕgP��	Z���cʬb�A����`��P�CS孜+��21^D�U:�o����5>�g�-�y�9�����~{Ώ}��n_�,{�N_e��E���Ȗ�}�H���k�)n_��.d"�u�Z������k��9�=�i��w2~x�Ë��I��p�;��hÂ���o���|iĈ����A�y|���T¡���w-�U�%�]�Gӓe���b��n9�)d�����Ǉ����>�C5S�R2��N�L\��hw�p>�i�u� $ǅZu�+Ŋ}Ĵ����������1�
:L���(�����y�-�O>�%L��5��ɐ:���;�f�0�r,���~�CxQv������4i�y�y�v�N�m�F�֜'E�kĜZM�rWݙY0��S�NnKB�ߴӕA���s�A��q8{�M�>^����������Oॠ���g3��z��x}i����M��?Q�g��Z��H)Z깍�
�"�����]�,ae�ڍ�ʪ/���{�c��c���,�'�ٻ�����F��P�3L"��[X�1�K��� 1�� �=���R�?&g%���2��C�ʩ�T��S��Xa��oR���j�'��(��r�N)}��ΖEp�C�
k݈ϿYTj���OH$&�Ж	��Ļ��×SaI�H��/����ؾ��O�2@�[�*�T�n1^#'U�5oE�R�����"�y�jQ���l��@[F9�]G�S��ghR.�lq�Y�p�=��S��g|�yE�C5^R��ʬh�X� �������jVk�>mAT�1��B�~�vl-�c1��@S�s=�g�_��Hݳ}�����������\��U"��p!-�������3��S��4�@�V��}g�J{��f�����9�{
�Ψ7	�j�x<Dz@������w�´LR���q�GW�e�|�R�d`k��h���eZU�����ϟ��N���+W�v��oK97�����e��]�������}!�H��-{Onk�D�M�`�èa@�!^/�*��c�kb&j����B�F6��p�SO�;E�~�l+<cj���ᐌj�H��A|�[bL�������^��$)_�]]�t�NH�n�T@��/^@�J��q���vՌ�cK��2�D��6~ഩ�bg�b�I�p���0
0D�I4U9�����%u�p�E����h'��_�����C�4ƛ���F��z�V&���Wa~�{]P����}���� �EP7��;j{���&C=M��+�ʁ�8kU���6X6�@�s��Q�+N~.B��l8mq��d��Q+Z1t� �d�Ѭ8����0�ƨ�����G�0�=�7CٙcjyݘtWX|0sf��a�p.Q������s�S�5z�7,Ү�d~n1p�N?Ȫ����0����2(߬��&H0-��:1��O�ŢɃ~�Z)����y��&n��e,ԉ�'��*5����
B�V�`Z!3&�hC�����ϻL0�Ypъ��tRY�C��ݯ��(����9K���[,f�+������&HK���s�"��,4�Q_�g5�ސ�ۨ)�����8C���֎����
K�i�'lK���	/��?�Y�*Q$%@�`�s�!�!*h�����g����M�Fʄ��EU��I��*�6AS4m��eD��-a&#�o����Y���<נ���L�-�9�.�gц��Lws�n�0��S��:��*�Pf�I��L�^��Fy�C����Nv�DL�Âp��ี+��ٵ��w��̬��D^a6�V����i	��<�=A� ��lP~�ꍴb-N�f��������bΤ����я! �T]�#�n*��_�[��D�~;Z�~��C�}��G45�L�_Cg��p������/� h��"�`���C/iqSV ~^�3����Wm����m!>��n���D�� S�@�w�zlC�rC4ma�@���U�v�����<�[7-����A4K �>�ELE�S/w9^���z� 7R�
$���7��,�̔�-I�9R���Hac X� ]���:*�.�.6i?Ec�*m�x�)��27T)G���-.���퍜���)��0��C���n���NB��Q'Z�b;e�D��'c����l8�5�����$%��i�����j���6����BpT���rZ��U��޴4ʎ¨�Pڣ���tA���n婿>�1�fyQ
ޟ�Un��2ݧW���+#x9y�7[!�	�2��P�ڥ_l�$�/�u�!$�$KT�GO
����]Y� �nZG�M��y֩�&�]����x%�������iyj��&��L�B[0>�
D����̣�M~5�R����?dk���툼.0�%�{V����o�'~��,j��ݱ�?@��w栅��ا��cd��s���'��N��	��v�[�[��9��,T|?�6���^d��Sor�>�>��cg�a2SF�ԗG4x�N�#�{B��Ue�,� �՜�o�^Q�v4,�$+���^v��Z	���$	���1`!6b�2�&d������v?_H
)0�&[�v G>���j��޿�/���)j���o�;��Ы}5�~r�
\����L��Wg�Q�Oz%� ?�ێ3�3:�7#�C��﯑J=���3cֶ��`��}6o`/頣��wL����;7[&�DÓb���y� ��'�/������,��L:O������h/�;��2� K0�lGM�]�J��~�C,�uo��c�QX��|@W�ϰ0�0���$�����h�8��g�d�m�#� _>��u;NJ�Iot� r�&wT ��5�w�����/���*����I4A��;���G�Hr�������C��H~�����D�&tw��Z6t����6�0�p9������sl�z8��{��̓1M"nKv�aP�~��W� a�;^�т�����;�{�H)c���,M`�u�3q�_�y�Y�Oj��%Wʤ���C����Hx��a��?�E}܈=c:'�};(0~��!W��c��n�ڇ��研2�q�F,(���b#��V.�6��Im�xbǌ&�A5���n����C�h\�^-26��zլ�����˅Rnn#+�e�R��#l}�%��o�R��1�e�P��ԤlD��m��Q��E{5���Z�*	��U9/���?1]t��pC	��<��Z&B(���ð
}4�C+Y��)rb9?�n���k丬��ge��ZP]f��=�����G�.�(�a�۞X�'��������^9}	���U���G�c`'U�a�y@ŭ�5\.��â����g��yHb��
��{��������x�����iF��,�-��Z� 4��.#
�{���d?��QR_G-B������#�$<��^����7��h�������r����q�K�q����
E4S㥄ËJYH%:�}�h&Ƈwp�{i��K4W����оJa�&A��5��r(%�1?��"t��':{'��7)iy���g�E��`��n]r��c�!��V@���	���Aj��`�40�e�:rX[����`'C�r���������ހ��{">����#��4���M�U��|��k�f�U��%|㼸���aR*X-м���I��mɋ@1�j�ե������^�T���[��^�/����vɟ�m�FbWbm���Xn�̔0�+�����ߐ�`#�-þ���#��䪕�u��αUu�=C��v��c����mBn��p-�ux����)P��>�t���r�ˊ���Mm����Hۙv�Ÿ�A��҇>����
C 7��d�3Qq�t����s��1�Q�;��x��.���k)��E��eUЇ�X=�C�)f�xY���e(����pJhs�=d>���g��g&�{Y�R�9o���w?�鞦�ta�E�1/=�"�E��;);bFLT�%��^2s.\~���T�;d畘+ݱzo|p�?��V#��$�S�H*KRM���keJ%��O���I�+'}��9tt຺z�27�x�
�T<���UL�>]��$�?�n�&�;��Y�	j�B�a�~���t$�5�߼mJL��TD����u�Gx�% �\�����B����=INX��G,P�@���������-��B��cy��5V�����:@�0S"��k�.�`׷RٵRX�?�Ǔ��b��}(A1��l��i��DJ93�����ܞ��sx�U�z�Pʈ��¥�h���eq|j_�q�	U���� 7�l@`p�$�c�}�7�����FD�0G��H^q~b=���rV�ܼeEd�� h����m��*��Wu���$M�G���[>;���O��s��n��z?V�wl����;��]�.ɖ�ޥ ��}����܅����k��i����z�fs��.�ϋ�P���k���1x`�=i6�)����� 14Y�4��l��TO!x�-���5�1�4�D�.��K��bҰ�hD�>\e��pu�6�[rv�(p֪�b��fk<9��2 ��O`NWy_Xf9��Ɵ��:ٔT��vO8&�5�h N�VJ���WMG7�m��_v�W32n��VP�#ݽ�R�<x@+�!dT�7G�v[gQ����	\���]q��[�^��Z�;I: G�1t��U��Pz0�eYԎ�~�RE�N,�����Wٺ��Vz�ce��2�������u=�tu���[��<����c��-b%W�wemHg��`.ڵ~���R��lZD��!�^��+�(��:��#P�\�p�ψ�4�t�ީ�Q?��'͝~�W��͹Og\.��,�6�`���(�Г�����:j����4^��_ehAix85��O6a��ZqA��5xLwoU
bӒ�P��o��i3o ��vr�k{:Ԍ̕�g�9q��\uw�N�i�3&���Z+ܕ|����,Z;������ ���^oU�)𳦮Q2���e��20�DJ7��U�U�.u*�ͮ�Q�Q[{�R �	6��Ѳథ��/�CZW) ����֭��sj|DGƟT�տ�K����_�#��z:��0"w�]�AB�Y�>q��sv�5&�z��i��K�l�  RE΀K�h,�Jȟ��
�������{�x��!�Q�Di��M�j-/6�9�%�U�L����kaT������Ӻ<�f���b&ʪ�N�+H�'������)����SW ��7#�0z��4��s�lV�`����kkUqs��j�hy�cW 4��MVھ���w�
w�^u�j�#N�4�%O- 4�����p7q�$no�H���Ө,},�*Q��6��r��(���|��0�x�|[x����I8��z�%��O �x��V���UE���7�ь����mR��$i6^� �`���e��橑8��)�.�[��=92��E�<Q�s�{n.� ��ߗ����U2���.���`ҢR�-�z$��B���M\$����qg�����=/k/�M������n�~3��X���3�1;�/��`�})�c��x��y=\�pD ����	�עW��M弐�ݹı�H�+`��7��������e���~�z�N�#��~jh��7�E�}�T��u�WV������T�O݈1[�'�:�G�9���s���7PH���L5h�/}��&�T�U����	�=��j�L�gbUӇ�tc�xsWO�!w4��&�\>6�Y\����X\&�b�u�s���; &ěC��h�E���{�87�Bkg��ʿH&����{�K֝w�1���z䩈jNٯ�뒅z_G��*^�M�i�>��H��������l����:�9d)����{��H�
�t�s�*���Jt�@o`��m#Қ��� CBes�����������@�0����ޫqtY��/�_q�WE	eT*��~�k��p�N��S��
�ѹQ� [�d��׿�`v�T*�5_նs;Z�n�K����{�%�ܪ���Ě�Dw�1��!�0?j,�Z�t�Y�5�g�����A�䜗�.�ʋ�Op/�x���1ǹ/��9����U�cG��� �ļ�!�͡��퉚n���R���#��B�L���힎��ut&��w#���T�s\;x{�aN�����{�{Qq��s�f!����k�; �ܴ�ѯ���<o�(���9*\�X��"�iJ0�*�����e2G0�H�~~�c�?zY��v	m/t+�o�������I�V�������L9��O��ĲT��@%���,4YV\��S]!�iK`F��~H��� �o���n3�-��w��G_�W ��`%���V93)�q5Q2\QhS�ԣ"�4RӦuR�@���g��.�}�T�H�H�m���πL�O��t�n*-��֒4�|�r����o�%oHy�R%�$�\
v���Ә��N����E�|����ݜSv����U� ߓ�a8��L@��3����ZK��S�ĳ#�Ճn��y�|,f��VΠ(b�BR�J:�D�$kI���iwtet+Q�8<(�6���ŕ\�c_�Ɏ'��91�ľ|�K�DKC�*FQ4Ҫ��Q@Q$Kk	��w7�:���ȅ��D�b�w��U6,{���ήN%L>31z�a�Lq�$��"$(+��[��`.2��.2��O᭰S�گ��+�Zѻ:�Rʓ˨�~��NZ�s�/��C�P[��Wl�1$�ǻm,;]8�tv��y܁����m`��Y���h҉}EE��i?�:����p�ݿM��	h� ��� o��k�l���s\"��	�6O��n;Q�Z`�������N�ZE�)�b^��c���gSu�jn�@��ERu$�d.�eO���=�3!�N�CRJ��[���]�A n��d2<a��F凋�J8�(�yI�)�ah��2X���Y�>�qj��e\e��d�i���J;&���]DL6�XQ<ʜ���j�կ�����<'����+�p߳�g�"��=U��~A/d�����4�Ag��Ϡ�o~KT�[��6��2l3�|a[F��ʙY�:�ړ�[���B��X�]�����4�����(9�����h�[}';"^�����xõ��f�>"�X������4�f�����&��zD�{�d�d�E�P[D;5U,]��U�׍��k4�>�6ʒxNz�-B4avy�i�
"���3��;%_�P��N������I7�_�0��
s����P�S/���X0��O�ۤ�-��:�ߣY"R{��?�T��g���3���2�07^*�q��{|�;�%���$�w��6�2�8g/3{�a�Ox.�U�'m���s	�� �;���tZ�]<Y�ZVI��������ӧ�+F��}S$�m��*�IE�ۊ]UR������COj���7jc���j6^���QܛUQ��:�n�����E�#�_'rJp���@`/�p�J-c�`cv��r�S��]S>uC�����A)�ٟ����#��4���"F���e�0����g����5���H��9�ö�VǱ�oh{�4���)��og��)2d��y��S	��0���`� Pf����7��z	��`&���1|��Q��9gH�ZQ��E�@a�Bo,�qX5������ZI ��x����/Q�V������+����)q���}͑y����@�T��������ݱ�����(���u���i�Y�4��*u/�
�C ~�-���$}���c�VS����PA���f/)�.���mc�FX^���<ȔL��w�����{���d%8��@Q4��aϟ7�b�ڱ�(��.Mܙ��grgf�Iz5hh�D��p��sCz�� r�I�cNؖ`�Y�C_RG���=���:+�m�3�	�S�{��80����"ᥘ^Iِ�S��&�JY�Э��,"�ǋ��8�&?7���K�yI�s8��k}����J��<�������L����JƁ��Qы7��>��Q��#��7?^G�K�41��ɀ�`B�Jh�ITJ�Z�8�S�?�p��M��~�!�y1����
[�|Z��$����v]znӸ���Y������4 ���據J������*�sX�։�Я^�<����;%���n ZH/ڿ�,$�ͺ_'6ղ��z/��o�%[uͼ�2-?��-�Lb�<k����y'���65>�r��ޠE��.a9zD�{Tm�PsT*�|��{<+�;���f+ۣ§j����q@�8�L�����^u��(�p�G<i|���,�Q+�VH�TT�'n�+5���Y� �����[���Q�di(]D�Ě:�1{n��MV����<�"���l��J'n~R+��1�O�q�i)i�1��i�V��o'����)���� �L1*�V��vؓ�pm���C0]����	!A4\�����A�o�&5? "�g���$�{cI�1PnbF�D &��ZN��<T�u���c5"A"�*�N<�k=��L�~h�0x�W����Ťm	��&�B�3k^)�*b_Wր���`C�<�O�"��wU�*���Po��[(����!�V�����+��v�4YάE<ܕ��Vy�IZ�yZM���!(�2�K��.�Ӳ��H��^���5Bռs�{{���\����9���
�A�of���ȗ'�I@�����R&��r�]g�p˲���:%�Ӵm~w��җ�.n3�IU�ݡt��m�@�'���&�ĺ��T��)v�0Ȱ��%U������v�^ksJI�b-\����������!�UA�������
+��Hx�]ܢ���l��t,֖*b��us�JUZ��f����,&(& �7ǩ��JT֓��8 ��R����%ZR�`Ҩ1����z�\���y�]ڀ*�5x54�Me��ȗ�B�
p����oQԮӰ6��E�*���&���H-� U�,��RBm3@Wݮ�;���[ǧ���u�6J?p���S;�Nڹm�[�0!ϝ6��i_[��r��}��3w��a^6����i����m6���v���*p�?�SJ��i�ꋐ��N0�j�(ZW���6<�
N�����X���H�����ly�姻��m�СPj_l�4�!����-�^P�\�N=d��}Eȏ�iF'��΅n=���u�xN�D|�TR�z:p�����^X�-�V��S���<���@Cts�S*]6$�8��R}\��0ٿ��!�T'.��V픜�R6�肺�s��E��(��Bc��J����4/L��muu��ZUȶID�UOOL�M������,,�|��]���K��b1�[����4[�Z�ٓkV�>�_>a��}�?7�d*�Y�b���jSl S�ڃ���W���Q�.e��y9��TE`j'�e��q���\,=��LNuy"YNgd�O �[���d>����'1�l_��6 Q/oD������\x	Dh!�g\�.p�n����	�l��
��)���T �,�C]�Y6���Ne��\���-ͺ��K�����`j�=�Y�"Ҥ�R5�6��7k��5���]��8�~/�1�$%�0�Ohk�ɗ�C�g��E"��絓'���Ŭ�c�9�/�������PHZ�Ņ���I�$�f���R_�����͎�rFz�,`��(ԇJ�r�Ac+b�
�j�O�������u|��<��d��������>����=-�@T/`4�^|��$�Hab9Epf��:�Lw�&�R�|`��\��cJw����U4w9�r)9@�j��k\���{|1���i�������_S�`�;��)j��w�&)飜��g�C��@rd�~�%�� 7�o��ٮ�8M�� �X���_�_�p�#���ũ�A*R��5.�њ�w�N�I��'��ǽ|�����sS���ɇk��*02�$L����z�deW�{�����;Dy�@�o!�C���3��y���l�K�I��;p����ǮDȐ5%���T4�X�}t��ڒ��+�J�=B s{��Y;�TG�$�
�!���?0FS�[�%�
�|0�|��O�DF@��;j�d��6k��]�@���٧�q|�1qCa��{t:�̟�>���U�:���,3�f�C�P#���R����f+�tF̧�O�P���U�1n]�?�E���i�t�[j�1)H�f���ꧧK��Z=LC�y�֫!0�l{g��bl(��g*��Z͑
KO�{���m�!��ǝ5�=�gS�$��Ӱ�X���5�㒦r�@�f�4��+zm_ñ�
S�kzB��!�yW9��S�������ڍ��OD�6�����T�&�탅�R��S��X��wd�rrI�@D�El#Ip�u��̈́�d�m�j�?�?���%(�J��V�M����2e;���fv��O���������~55��ޡCɻ�4�=�/%�4�'x0�)�ld�fc��s.�����c�+<Yq����GwY�X��a�:��>�_�v��.�KB&�J��!L�5Ζ��6��י�'��Tp~�C�j��FyO�M��_I�������Φ������Q�}�w��Է�������+(��[��<�,]m�1���o v?�`�I=S1��$���uq��1����9��AMT���n�T�=��R�o�`(=��
ͽMĀ�o��I\�|π�I5�'���5mS�jn��l��O�A�)K!�t$�.�.���y�"H};���ΰz�A�A��b��ʞ��a��@�/��{���?�`U��0��y��iqxl�dW�QzǶ�?�㱭���z/�xw�e���S0vz�괫���ʶ�Q>�dЛ'pi��yS��N>c��˫v�CW�w;එh�;�R�'ֲ2φ�0o�
Cq/����")��_#�\C�R�\o�)N��޼�*X%j'E�;�����V���Ƭ��5�ߌ���4�ن�D�m��@Y�k.+�
N�m���[9`������_}���&.�o���Lg����*B�Ja7�⻺45���c���4H���$٫`��9M�+Hrt>ht�471d =[K��q^�U�:�r��:2!�A�i��x��2�5i�1�,O� S��(��D�X�ua���a͆�+?���v��H/=L���wqݏ��^��ZA���m~�+G�O�u�̎`��΂Ó����1m���nxg�p��h���`�C�ԁ:���Ni�
:��t��BIE�D�������qS{6��%�����ue0�e) �4���v��+�V�H����K������<�|�ۗ:Ȕ�Sɑ=�v��
�U�uLF�zWy�\�Ѭ�sF�6^:��|����}�,��O�N�n�2��F�t�JG_N.�仁Ԇ��}|"�<8!P��a�I9S
�3�[ύ�V1Hm����y!�O�bŸѹkՍKpO)x�������u�;XЯ�J�y����bώ�sx��ד��[�D��L�|�v��[�U�t�s��8gkd-��H�P��l`���Cg�W*��"�JQx�/ Sygr�7@]�d2�0 耒���:�3�um'�L����Ȧ�։.�� �8����O��f��>�uOQ襜|rƝ,yՐX��aY����KIԌ��a|���rb:5AvU��F�����1H�PVo��մ6d�����Q�� �N�ǭ�qlzy�����t_��Cq�J}�����#mBmd߷�=��.���Am7�|����3Q��q.E��޺	����{���K�7���e���̨����� �}�F���8ٮN��?��_/T��rk'`I��$5� � �Dv����+*�`�`��_��Q�Z��-7y�e�0W�h�
C�����
���8�K��`<]~ (���T���0�n�\'L����uZ�p/���L�	EK���I[� 玧�$��tG3$Կ
Z1�9�"�H�� .�H9�f���c(��P\�����B(�xg�{~�\s(����x(��x��*�&��	�5�?�[��	�q~@�R��0r�j¨d�b��{��	1eU~�#�����*��G�H����m��VXm�X���Z�Z#{.Gv~�o}�ߨ���C(˫p�B���#�E������qr(�-�����.Hhf\��P��%Yh;�W�K^�Nf%I��Չ �kE�E�s1t�m(d��*~��$��[h�jiKȜpIi�eyv�iq���8#����<<'Xa�2����^�� �����*�nH����YI�j����9�������uIg��	��ݿ��="i�}Ed�������� �X�z���^VJ�)-��V�����X�X8J{��}�pzh�B�8V쐄6��*����dE��Ǡ�}W�Q��o��,]~c/qC���)&3�{�;���-������j�%)�=;�OC�Ģ��[È6
�@��[�p>lt��#{<8S[��#f���!!w�u v�(�cߌ{�-Ŕܡ�/�����U�a�e)<�Na���g	��CEb��6�Q�s5�5�����tTl��[��G+٘' �����P�Z�M=A����:Z���EL������f��3�xqfx}�cp=Zc�r�ğ3�f~ ̿����QXs=hX3Qh����v�
�]�H#&�����
����Z�bP�#%��~��� ��-N&a(�,	���O0���ۉ�2�Q�(�.!��9�|�	��@���&����Ii�ܖ�)m��ʮ���9�e^�j����P^����J����39<�҈����Ð�yj7̧�ȵ�����^�;��tDud������Їa�|�hpG���X��{"E�˫��%���ֲ��.�#ܺ���&P�-ЗP0w4�gӴfI-ڮ��k�8�~S�P��5ĜXu�S%�3J ���Y��\�	O�L���Y�P�A�` ��%����sx7�F5{Au�呣<a�b���#
�>Ȅ�����P�v��W��;�d���a/R�e+j�h�z�m���%\��> SM/�U�b���"��r!L���\΢S��:Y��/O#Y&�[oJ;H��T���7�U�ge$���	��`��c��,���C��$�p�e��Z�kqm:MmN{Q�-,a�ܣ�e�i%�z��ߔ�A�#44 "L�`P9U�G��#za�R�PؐY���c���:Ods5����E��kk���7<ڭ5~�ZX��κ�@up��m)z��ri��EC���:o�-�L�R\��<�X[���]����I�����2n�%c~����H��/Ti�n��t<<:�!0��k��~�+�!�O�22Dtl�ϖ{%�S�l�ڗ�����i����+0{nE&���n�`�4����誱�9�󶄦�*g9y��v����E'�C~�d���j����W�m�z�����Ak��gG�K�*K�3^��\�͋ESE-Q�^��u��|y�nQ�5Z�x-�%�	oZC+��4��]]�,&���-m��	�˾����9�(l#@����x�Ќ��^��8���y����sPX*B�|*1pJz����XzZ��5��8������:�n��������\�`��<�|�n�z^]�rMX��-<�L*~��tE�n�x�Ǳ{�3��Z=��D~`�Z��J��cw��d�QE���0N���hh�R�e'0��o��i&�Y!\��.�Q3�q�y�2:��b�}$����%/DkZ��!E'9`
�+����+i���g�rR�0�#�i�镒k;�i�����~�
i7��Y�d+ip=��t̚���Ȣd�X�B�f8@'(]����U��K�+�,�.7<*Fߩ�n�J�5K�I�N��&�&�Jt+��L�Z��*�
��� x{V}Z�X�O���b����Ɉ���!�A�=���_��/q�+I��� ���U \ ��ju�;7�W;�Lu���*��U�3N��B7ٯ�e/�8��ny=�T�B�.�q��0(�	���4=�lkn�v�t<.c�5��4�PE�]ߩo��~���w&ttUz���z˘j{;9��[D�Z�`�_��}X�L���UD����4i���˻���*���D[���/�	Ж��;
6^�m	��yrG��g�dy��Id�69!I�yl/�Ov4� �y�J�|V�P����Uy��	��}&�����TC&�{����&�K�&f��c�`M,�L�X��Z��q�� �kR��[�𑔂1����r��/�~@���A�8�f7!���%��p	T(�����Ǟ"����I�t��!��YT(����⥻v�f�aǉ{���ܨj�
����E{�lU�⊶<iV"���Ƙl�2�P��==�3����fY��[��U0����4މRI��������Z� �O���f��Q?��iA�R����Ds��ƷDP��!��7�O�j5K�
���CP��EvF���>���`tK�my>Y"h����(��S�j�d���Si <H�t#��y�;��z1�Ͼ�����9kzЉ������"g8y+0��	��EKA��X��z��|�v�3�H�ҹ�N�,����C�$�+Ƀ�V�����`��RmX�[��v<�m���0�=�y�c2��G?���텞Vt�eew�+��)���7n:T~[����xJ�	C{��~d�=�t�e�[g� �3d���Q*�~��ˁ4(@r�|��*�(����?��C�DR˔iO��J�s~#=�w4�觽�{[^�\Bb�-�G�IlXe�?�p��67��F)b����6�������pb���}4�1
Ϛ��� ������`���b"-���Zf�ݩ>Yؗ����DW	ɢ2wv��� ;muM�m��:��������\"s_[D����5��E�
�*"vɡ�`c�Eb�}�����Q��M2�ٟ����/���i��3'1H�e�
��D�?��?XQa�;��.o�^�^��Z%�+��HXL[�%�>�M.����Po��3
-Ɔ�Ҍ	��A$LCo�l����塣�~g	:c]9�8}��Ǎ�Qc<���2���q*��N~*�$��_\��B�D?9Mq�S�v���� e�Y����V���O�#�2an't�����c:�UM*�|�6�*�7~�m=E8P�����b��G���CsD��^~Ib�e3��!����U~�q@���z2a�1Ѧ�'�9:]�L���U?c���w)��d����r�Ĳ״Z%$��=�@�k��j�J�A�(׽ٮ`����"�i�t�3<7���]�'�Tv ��o��T��)���m�kp������I����9�"�6��,��i���ZL�����\����6����X�kO?�S�t�Pmb6a��������\Z�4Ƌ˱�����]�Nl�Cu<ᒫXR"N��h�]��*}4,��V���@~6W�-|��8��v����T|*�4���dd^�gG� }i��ʥ�u����s
V�[��
�_�SJeGa�^#gf		T��r�k=r�]ݝh�h<�Z���pN$n'V���z������f}ԲK���)*�*Y�$��i_!�(/YD�kQU5�pd�<p��̙�8�@r��5�Օ��=9���ݓy�!�O�ۭڃs���:,b:�=r�	7#�x�9ī[��[!!�]}�h�ub]�o6�ua�����!��c����9�I(Er�J�1*e T5Ǯ���%.��W���ߐ���!ИO�cю����H���̵cZ���%��u�d�lu4��=&���LL�{&?��Ґ�<��.]����*�>�0y�<���~ �x߬�bGoa�s_t$�S9>�Y+��:���K�8]�P�������#
�8}�	�9�R�a�x�O4K8�G�@�&	��K/���`W��E�ٯy�;M�p�Uo"+�e������zf��B��o6X��L@� c�I�xV���`?�����4-~�.���p�.%H��^��E�N�Z���*Q*i.C���.u1��E�isr�W��Nk�BƮ�q$`w�:���2���$��ߤ��_~��ő��픉&��7S�ɩ,��Kq
�N��O�tYR�OKٲI�.�N�0S9${��7ۨ���W��-(K�\�4���aޱl�\���\3��8��n�n/[ 9L�s	l�U�>��o��޷�sU#}W��Ȳ��~t������<�#��}>���Kaxb����fs,m�2�}��^aa�`�(�HJd��c;T���:�L�J���1���p]؝V-_!*��1AD*�	�>�\l�c�,�3�4֐��K���H����n]�K'�������?�贅,6g��Bz�O{�Xч_.���<W�
CZQ���ߩ2]Mg0���V�h���5���(�T9��������`�P���q"�ع�="��\�A��S	��XvE�K�ph�������u�1��N
˙�O6%�@=�$��Ê>��~t�9�YLq���{��	�=!x���T<UR"M����e��h�]EZ-��T�P�As����nKp��%Y'L"3!Ӡ�W|���HU����H�T�Lh彴�)�9�x� "d)4�3���-����gU�r��a_l�{�"(��Q�{�����$�
�r������u��'y�|L���C|��a������N��6r�!%�|A�����R-�Z 1�H�\��g�I�+���t�w۪
9�����6g��	����j<?�X]���GJ{��_��I�v_��c
 >��׃����8�|u	��:����V�\�?="�5��X�%�/T-`������M���2\�
�^IN m<]~�����>�V"�	�mC�d4�q�4<���z���&��������B��q{s���1��T�z[ۄș�z������%N�G*���	X��p Y �� �C?PiZ]4��"�g}�D�l�"i8;i�'g���>D����V��O�h ��Hg{o-�"�@�3{MDޛF�~�$�y2���v]�O0\��?��?)9�� ��Bb"�����T@,��aދ��$��(�,���P@ WH���=?MQ7^\I$����^8 �j���6��54ׯm��ٯ3��[�
a$���ۛS������9|�Vp�x�\2����iL��p�P&;W¨��k	��>�-���*���^�*�e5�*�C"+[Q|��{w��#�((���+J���x�����2F"z�*�4-�A�����O�Q~Y�n�����lx�R4*�����!�W.͋� ok�њa���W��"�����4�z��L)l5�F���ぐ�~	��s�����!<a#�p��p߲N+���:�(f+_��8�3��U뜯�cQ�n�Z*���3��<ž!���W���� ڗ�x��g`{r�Y�7��
�┦�W��.����������W�9+�5�c<A+����)����{�LAM�p�,�.��QjV��n�~��sA����ښ�HD��!�p���W�pgp�P+�����U7�4�f��fǯ��&Gd�|��2������������:�V��=ќ�m�ٗq�˾V��[; �0� ��,d��I���d$f"�GF[�M�!{e�8�6%'���XΕ��
�N^i�ozs-IY4��>������������)o	�.(�1@��ł��/�*Do��{r��Ī�4��
����SpcN�V�% �� ����j�q�ڏ�/���l�O�}]�&2Gִ�VI�����`B��-�R8�f�Ϙ���ଡ଼��oy0�J�q�0��`ԕ��<߈:f%��L٩�^pe�����n�a)
b����&��r�|��S9�@��1�e������*�فb�A�6�գ
�����=�UȠd�^�1P=��O�!j>M���!H�d�.+5<��!!)�x��3oy�{h,��F��~^�`�JR�Wҕ��E�����k��_��Yg��V F��g���oJ����Oq5��ּ��r��ɽ[Qj�� �^wެD:	r�O�������)d����`m Y�d�=g���%Ýd��,�4Oh}e�(uYN�����������_�B����{�"�>�	|�-{�3`��9�g�_e;r�#�����I|����Sē�*�qb<��n�u��}�޶�jc����f�@]�g$���n�=��0����J��Pd}`ݣ"b�:�A�Ð�QZ�k���]]�b=D��|w���%��q�Eg����F�<·/=�h���<��#F~��N���ذ����d!�������,�Bi[��Y:�{�&�,�!,9�;jb�;(��%�I�<P�k_�R�7�6����:N��H�;�@����ά"�:�;��Q�{�ca�<�k^Y�5{��]�WMb��/1�A����WDNC1��n��aj"�`���M����i���ܭ�\���L��7e� և^�!o� ϓ�ų� M�* �`߹h�o��|�@�.��{�K�gb�ӻ��H$��Dss>�WS9���S�fx��r[T%��(8�X[�%�`����>�T:������xX��2�������@�k{�o��q̽���S�Fm߻�?��U���E��}��t�W���`48���f��,�'���l��W�C�C�y������$e�lk�+>0�[p����W�$:W
L��J��Lj�q&NB���9�������8��òO�O�|Ԋ>p�*����yY���,u"ɷ��H��j��z��R�Z���-�4�o�[͇�B,I)(���xh�P�ᡁ*R�Mg���+0u�Au�8�-d['\���7�ce����Q}?�Ě���J�����i�9c�iF�(,����~>�l�g�����2��7F͡���P�����D$I�ͨ����ϻ�_�+M||�C�NNQ�U�`���gP�B���^�-���h\�/3{���Υ�G�+W$���/��d�)��s�Q�.-�0O��o�>Wa���Wܢe��h��]Iͫ鿁�ou�=����*�+�{��]&�-
� �d���aNf�*zC��{���u��K��i��6R�2���G�S��~Q *���!<�,>w�C�k�OS�ɏ!�"C�o��fK�k�����]_a��P�{�l=���O�c����r�'��i�'h�c
��<A� D�leE��[�4�!������x��3�jawF>Î�����ix}Wb�������q`�iw�@9�Y����<�5���z�K�o�ܲ!�����\'���TC�̼�^�Z4Jf��'�t��)���Z4�z�m�,nV(����k��p�Ep2$#��`���GC���,�b{�NX���ϗ��V1��gz�#[�0�ƻ����w64l/5�0�������:�c~t�VAM`��aN��K�9�us�zeAMZ���d�kS���[�mi��/ʄ��pnE	'�=�Ooya�`��JқJ<�;�63x͟�G�����6�;��Q}��ԁA�Q�j0N�}���11�u��_뫿��Ѵ��(B$bTG��>����k53rb]�����E[Z�X��d���p�o�4�TU0������i!q�|��N�e��oӃ�ϫ�x��T��k�=�蓌�ΓC:��|
,�	���!쁪���*(MI����AG}ۂ5���-�<�x4������w)lL�`�F�@����¡O�%j����-KZu;�C�����6y��z��O���hS�c��ofRy�-���g[vZ��/�an�
"G ������8��[�oħ�d�0!G	�`XD=� ���� %��PL]&k��� ����>�XA�Y⹓)A�;�ܾc ����l ��t���֑�)*=��4����d�<$�
r�2΢͌�����@<��-��ý���G�&m+idxz���M�Lv{}����2����u]\b�������j{��#҈:��bÐ7q�R�2�`Wr���jmW�pDJw��
+��n� �ÏH��m(����?�]̜��7h/���9��zfZI���[/SD�`R�s1Cv�23�%Q����;dhN
PY|���`�q��{�t/�T�6��(��AP�����zq�2���m��w3�b��-/f؂y�5+��[0�oԜ���Ϲ!ָ�6K�M_�����	�V�ʢxن
:����Q����5�ut�d��ݻo�5ؼ"!��&��,2�7�iE��TG�����9��d2嗓#�A��aR�w�d��ޫ��
�
&�)�[�PK�=s��W���<+�	���0��v,���
�̇�B�xr����8����]��è�?	��9kjXn���R�o�w����8�dBmv����؛� �rVA_� �}��ItQ��.ѣQ��J;����m!�J��y�Z�-]�&�4~s�ؾ�l�=��+9�k�r�m?�RTTJ9�y��|�_�ZX�]n��
��k��q�n�nQ�;M��0]zGˉ"Ξ���la}��7���G{BLkm�IIj��J6�Y~T����*�Mt��:i��Pc�4�ay=pS�<����)T�+���E1q@�C��k�	T)#B:'3�` ���]5}��rCw�vF٧�C}����Pr$�˔�~M/Ie{�N_)����6�+A��mZ�(�W8�*�w4Ć�*����l���Hw��k;�N�>&\ ��~�WI�=yHZ���}>�@"ZkB�pqp�����4�~�;#�W�y[���m�s�m��o�о���^}�l�M��\����h�o% ш����f����M⬨|{w��X����:�^kG��c$F�i��l(�^g6&Nf1az�h;5
C�/��+�2ph{�[q����à�3��o{�O�SK���Np��@��0�̜Z^*�8��?aj�=qW�z����X��1�R�&c�Q/��y��'���<�.�6K\鎖6�N	�ay��w���Li��C�.�P�=�y��3�XlJ?@��aV��AP����9	\�W�F��`+�ʱ�an�Zu��o_�9\8?����;$	��qQ����w���c������!��ƭ="I���(H���MP��}n���M�[��HSx�@W�3��3uf�u	y�r�x'��S<`ŦO��U��lޚ�x�6�D���i��X�=� &�Pe�O�)p�(�V`i)1�{��#B?�̊{�T�	bR�?3c؁y��2
*�4�IPA�J����f���@A�
�;Vz��;���p����|�!e�z��?6x����d`����5���?Y)!�(�ÿ0�Jg��m��)O�@j��Tvl9齟1�϶��*4ٚ)�O�jC/T�R�v_O�P���j�����u謜�}l�^��?Y>P���
s��g /�W�����~��fCvL"7�Ix�������v��$���f.���w�4�G�(R{J�Td�A�pC���7�߅��ӯ��H�Ψ�u]d�S��"gܨ�扈�>���ܺ]1d�^YL/�}ì��$"W�J��Qv׎���0��B��{�
��D��B�đV#�=���*2��,�p�)��O�m׃�\0�����溸:�@/DmJut�4��3�=����M��`�;x�H���Ch ��$d0���ޠ��#7���8�df�-0�E�h+�*K�T2����I�?�Q}��T��d+	mb�E��2$�v
VqQ�'���)�����C�_ d�TH�J�����I�L�k�P�l�^٥�b��076=�m��ӝvi�2���M���=?>�hX	��'0�f��5���d��P�Eȯa�*��B,`]#�<Ø�'@4�
/�Z� j݃-WWؾ?"�?ʃ	���}q�X�D���p5~��=f��,���Ʒ��+|! 0�e�yIX����A'��{�����l��;
�ې}����/����F�O��@��ڿ� �'��fY�&nO�������Uk�+L�����P���n�$$Q̍��f,����`_��䁼Ie��w��$*�P¡k�4�#!�TA��da��p&�?��;'���S�jL�~�d����Uk�ŤI���ݐΪ�Q�d��LNr���/���P�ه�.s���3B�!�BR�#�^^�I&�:|A���榢YΗ��:���E�'� �2��c��J_��K�ԋ����<]�uW�<qPV�C��۝0���kO:�f�wG5�5�F2��
4@�cy�Ța��Mڳ�ί<�[n��0����j�X�	�B�|<jI��Ñs	*�T~0g���Ҥ�IM�$�K�%������% ����Kf���&��mŞ�T`�g :���Y��h)
��+¸�1Aj8���p����n/A���E�{
W���$g��S"�%E��^L�(2o�3�~-Q���Hٓ2-��\��"��V7�r�;m�q���$5�k����;&���གྷJйT�l���%�,�*(����j*���@�� v.0��֊���D��Tw ���	�cGi���
�?��JG`+�
��\q8d��ZQ�a%�आP���OZ��Q��e�\��Fӵ��=TyP�@�L�s"�/B�O��4o
ǒ�ǃ��Ž��_1Y��Œ��F����\���}���(�=���(�W3�����In�J���؆�
���,�9�C5�5?nT�iݑ��������=�f<�#n�����s|DF���Sd{5� ��aR�4��w���y�{�T��=k\t�f/�(t�!ƎT��w0cj��П�G17,��n���L�^:�e�H��޴����^FN�Vq��с��=жɚ+�3g����V"�?v�v�0�[	�Oxu���ih��(E���A��i�v��Bd�!$=b��4&ޤ[E^�ڌΐ��AtM�꽊�>;��Q� ��ȴ<o-�����)��t�/nFN��Ʌ���bY�L�|�^��6-*G_��_���X	�(���K��(%*=�tSD
G�����+�z�e��g��k^#Gf�WrQ^V�7�ex�&��{��k��M������4��e ��p4������"� U�g[�/9����D$��%�d�h�P�j��+e����� ��5�xp�x����w��-ɺA0���py%���x��}���)F2kb�=�[�w����M��JB�ƣ>s4�,�؅��Q�>��s��A��vV�f��7�u��	>Qg�5�����l����=f^���B0���i"�Z)N@�::�ˀ���~WPנ~�k�_��34�H����@X���ƨ�� �%�_�p�;IЂ�`6ӟЉ����%�ϡ�����F���<'��.T��2ش�hN��&-)}�9뽿��E4P+I6꘷��{���h��J���qh�D����_�g^�f�k-�� �Shf�hP��l�Bܲ�d�=�o+�u�Q�B�p �
t���w�������!}�Gɸ�&iXy\o�q��z 1��� ��2w��"ܐ��m�J?�A�&y6K�X-��lޮX��RFO��Wr�7M��7O����?�e( ����7��D���A8$[�ok�oЪ�M���S�_}<Y z�I�ƚ����FV�^��%蝛��!Yxiیֵd�j��W֘�d`���t�=��;�R���!N
�Γ;�ǈs�KV+�H	Ѫ^�".�����B�����:Wn�sH|}�;����)N�k鯦"��_�Ά����jD���3=�ҟ5�K�m�Cw�F!wD�5�BI���	����� �*ŝT�߼�~(�X��!+B,�9�r���U/k��7b4�x+ɰПA�^�����g��`B)/kY7�c �8`S�e���͘({�Һ��̹��7;�˵�D��7p�p�5�>�b�`������N�z�M�Դ��\���FT���ê��hfK+�$"��������2���<�t8��N���Hc��;�o�Ҙ�������0$3%�s�t`��ҧ	_�,�
F����`�㛀�ͮ��D�+�Ǌ��,:qȭsb/�9��4��EQ�4�G����{= �:��2��YRN(�[b�[�"Qm��l��7ݖs�Ub�d1�	T��s�q�-��K� q�H�h.@S�U�(D?vX�w�c����kԒ�w�n��O�'��.���������_�#�T�в�^/'��& �{�#�k��P�S�������^)A�@��P#���$=\������58V��l/q�oݴQ[V�/�];&7$�ύ�G���mT�Gd0�U�!W���h�	��=�D�9��vLoU_����u�7�k�k�<�H�L�0��Ytɮ8Gs����D��%�C��l(7��0��Վ��~�3%q�rju�1�-(�{������B*~����_�]^�QQ:_��V>����^����qa��⊃ct�$�ݜ/d��R����cq�{���O�,Qs��q��Z��lɂ��=�F]�%5����o_̾Ho��"
S�����51T�$�|�q@�G���������0c��0�2i�N��0�ywh�I.aI	�X��m��Zً�Ƙ��[������J����2�N>�8�<f������H�ۈA�i�ڂ��@!�`U��HaLE7���
.��I�
�E<�n���X � #�����
��T��y2_ʴ��r���i� !���2��+ǎ�m�L��v��	�<�QCA�c�����8u��RxMK��K/����W�7;2�;AR���إyAH�w}T1E?�$ɨ��^��ǐi�U�p���#ۮTM��n�����\�QyH|��f���x=;�Ә�9��SA Ʊ)����"T�j-�|�eVð�Ղ����m��}b��h�|BBO��ڕN�n��t��?�nՏg'��t��ވ��^\:�s�����%a���hS������e�?`����f���Uݿ�.+
i^4��Gek,�����u�����	�g�W'j3�2ӈ2F�4�OG>�ڜ;¾��b��ä����Q��������f����Iw�UU�U�Q����+�/��_�L��	i$�沸@�kh4�=�+T�΅	�A|���W��|KBjl�z�7�(�X��
_�ߚ7��&]�����U?S
ڑ4�;������5a���4yU8Q�I���!vJגf/.g�L�	q�����"��+;����%�V�geۢ��^���,�B̕�@�q��b��u���H�z�me�d'�G�&�Ar����6ˮS^�f7@������n�P���V���]�e20��Y�۞֋���y`"E��Qo��v�)���v�%;P2��<N7ysx.����ˡ�ݝ����5D/�+�K)w�ߒ�%b�'���0�I���%��!��$�����]u74��OPq\��D�x!�$r8ے&���:G_K������D�A.R��n�k��77�+DS��0�"����GN��z �r��b�	�ňI���+O�n]D|Re�1ŷ��+D?4T3h�����;8n���{9����Pm��l4t�J�#�� p�zSrv�p���(j��R�AГ�:�����`П��'�^�k �� LqbSN��T;� ���������^S��h���j��-7�)�>�#��5�D��ߚn���W�Am@%�����p�t����'Z	X�4-������T�*+����̕\�dv� stp�d���@g:;����K�5;��b��3��?�x��M�#Q�:OJ���1����W'W��H����ϸ/6�C~H�q �V�����u{,xf�X��x����m�t�������ھ'����8�h=���+��6���R�/>�D�*n)��22.�y7x�����7�^A����|-�LyH�O�O��o�c�'��W������"g)g(�EM���0�y$W4# 1+�Eɺ�v�iĨa-���R��]g�S����q�,!GN�zd�mƗ����$��N�6�V޽�[������ I�?�"�?jO��|$�j�@��&$�<�Zlߧڍ��R���J��x/,�:���)�����"hgO�	�B��r��؜�d��SУ`�. �J�z��v�z[���,x���>F=2�, �q�Y���R>^,����p[�I��~]!�TC���ڏ�#��/��0Z�L�a�*�R9�f+';��Lx�1�������^3��$6Yl��LFr��5��n�hnlm��~�`*��7D�i��:Swd���V:�%(���v��c�a�M����#[զ�n�.��;Y�阬���>��T �z�z�,Mp�tGo:&~mn�ts�9N���`ľ
9�MyR����a:������J�$ø����D�q�oɪ��+���AI���_��R�$���P*��R^��?bڡ��(�Z��3��A�#u��""�b`Xx��![:ѱ��<ή�_	��~����*��2 ���o�]��H"��z�7{�������?����;q{�{�r��>оg�6�Lm7��?e�	v�Y`�_��G�SG1ɜetX04�ͅU#�����`�P���#Z��y��'��>�񳲸+��9�y�ea*X�$ٕ롴��i�Fw,��p�)Q}�}�h�.������I5���AM�l�*D~ߐf�{��y<!�0�\�JwGp���E�Q��U���.h!���#�Mf�[�I4�L����$��햞 ���W��H��;t(�d��n��ƛ`@�� ��Pv=4Ϣ#'��/'�!8,�e��FZY��)��og@��0t��"�IK6��4�<9�,[��er8�����G�w7�հl�#��P��{��ь���Q3�}�6�R���3ZVA*��m��G��o�ԥ����'�>@S߳��!i*^T�߁���"u� ɟ�d#��6~���ڹn��g>X����}vU���*�A"U���{��vA%W���~�uݩ�?���	�'q����f>�*l���M��OӔ��}��z��b��t�<5
���e�׊���x��)i���uv/P�߭�l������Z�e�[��,��4e�K���~����nxap����~*Z	��������v%Q{��;p���CgH ^���e�,R�%��&��,�*���~A��)j�=ePHWG�#%�I$W�zȂ��ue��I.�h���6�|=&G�m�6�bB���Ur���Bd�g�ǝ
�]<*�N�2�[��^C�ꓘ�tE��ϒ�G���tA�m�;�������	 �D�"�<�F���aKrC�V.�0Ԣ�b#�N�Gq��T�vG����[�й8�[{�
Z&O��C�R���3�$��`p��缃�}��@w�`f�wik�=�I���h���g�<�S�]�z"pЊ $��h��O�pB��x5�T����B�\j6��)<1���4/���{wf��:���:IH�7�ӣǌ;N-���&�k���V�)�~��*�dI��-\#��ш�0���`��5��W��11�,S��ja<�u�Ԅ��ӔpMu8���7�`RtR�d&�0D{k������K�4Sa��<�����o�ʪ"ZM/�EB˂ﲰ�H��J<�t�G��i{���}�p+16?���X [���Ѵ�^�8����Q1>�
9��yvW#�U%�<s��X"��jԶ��>*m�n��^r����)q/|)�$GO�4\ ���A�����'�*���?f�V{�[ʉ>Z�*8(x�t3�����oZ#]u5��$:��Gv�%@
#̄� �#O���&oH��.;�{��w��4$�!k�ٵ&���Vh��򍽿�.+��p���٨��d���^�7�t��-��Y9J������
2��{��޶U���w��mန3��_]k��r>��f9�f�������S+!�Gq��y,���Q��R^�kA  ŷIHe�x����L,�Տ=�$a�zQ��&9 �="2(R���f{8.���) Oe��C�`Ϻ!�Ej�z�+Ԝ�U��Mm��W� �D���O�V�i0�����\Y�C�v�o�a/�
5'�����d��͵�%36�|��)�uF���3�B����b۞����6L�d�yI,#=f���yc�o������^��o�<	m3L�s�H����_��>ј����]i�����Z	�/�����ARÅ��\H�-e�Phъ��"�d�f[h�td�`��(q0��r�#6��kRT�N�w,��,���2�Ag�[~'�*w!G�+��h@�è����b\sg���m%��\�䵨�
���,����rG�~�n�(��f��7@�Xp�fS�H���|.-#Y�h��,���&Zo��d�S-���Y(ɦ���!a��� �L�q/6	e�P���3���6��������gFexz�m��h�>�O�a�c�?OX��Ì�ٮ>5����\���?�~x�N)�glrܷ�gF�x�`�cFg( 2�	!�nNPԷ�ԍJT#�B3�T�#eY6��v�[�!@��
,�#��4�38����20n��p�W�y�<̈���3JG�T��:c����F����ƈmu�j1�7�*�I��8��7�9�Z���x�w��D#F*9r�����mD�Q����K��CKˍ(�3�9I�)(H�	��˜xo��6R�N�R9�3e7�}ٜK�����F�6:t.�رZ����J�&uW�Ir����nt!li�-���ئ�A������=�$E���#�N��a"a���5�c��b�I��Ѡ�cޅ�.>r�s���8>�D+V֑��\I�;%�@ �4�V���5^(���J��_���9�ऋyI4�ُ�-|�.�i�.EI$�����O��Z]J ��'�qr˿A�h
�����[i $y��'9s�ٸe+}F�Jw=�Q�^0��;�/9��-�Cnyͱ�<$Z��@�؀��ưj�6�n���Wtb��c�g\������'��u:G$����7'��Π��
R�@�ֻ������:�j��Ǳ�`:<:aQ2d2}4�}j�5U`a�Sn��zܞl,w1ό��ɏ����(I�-c?i $N�Q-Ȍ����\i�}���^~����'	���I�,�#DD�K�I
���Isғ���c�p��W&X�Ps���=�]����mT�f�Z�	����k�����ǚL�E��Ճ�@�,����z��3y&"BH��z�3�1	��q�����y��P_�h�Z݊�*7E�̲���<G���7�P���W��џ�o�������:>s�:�P�fzq7f�<��;�9�{��ǚ߈�����=�5/fu�<O�<;�M�	�x����� F�����Eq�)}O��U����=u۪�C�$�h��IT8�M
�U����l�>��b�=:�?�0��(��≵9O2p�����6O4+���:s��S�7�"�|�-��`'��2�+ (� >y���UQ����$��F���ħ]Ư ����\�������#��n����r0:�)EQ|g�Ƃ���:���5���V��6��_9 A���Pq�4�(�ʭ�9�R4�>���[�X�'�����m�B�G 0�*B�eڵE���'�A�%��;)�Ö�Ӳ��?+N�k~a C/���Dw$�^J_1�R�v5�Z.���,a����ZB;�=�iZ^xVK(h�*�Z]Gu����D~�g�΅
x���-�{YB��\�1�Js��t�eo�,8n�����B�@K�╼�k������� B����8���xQt	�.TL�]�ԑ�7�6�j��~�wD�ް����` �KD��.��5��i����f<�fm
�v�Bߒ�sQ�[���y_ƙ�=bC��]����?�E�k�����4b��&����(Qo�;E8��+�p��]����`�o����a�5Jr ��wG;x���5�Ӈ��V�rK��'�̆��%T;lj��J�����_���*XM�İ*���;O2��J�ƾPG�М�j�>$����t��0	 ��jҿ�~�@�e<0�g���[b��sN��j������Ŭ�M�	M���ǤE}(Ia|T���˼o0<$���fIG��C�Ȭ˯���8'{E[_���s��']�nβ��p�gc�lZ�����|cv�r��Ǆ����/aVy�q���k(/��"8�i2IX+�,|��Z7�k��r3J$��/p�nb,�ϓD*z�T�b�T�k�C����6��8j��̿�b]���^�/�-��f,��TY�eTO��4��`y�ŀ���&$�=C�&/Έ$�ژ���*{�]������<�ܭ6mk�Tm�p� 0�UBl]��k-�ϙC�j	;�W�:�ό�~�s�;��_��u9��� '6v��5l�9owO=Cא��붉�?/(�I�3�����f^��^.�{�;��B-1�͋� ��CgA���P����?G ]��)���6��Y�0<�'x�O��	g�����*�S����yo��2N#�x�frT��0<���Tq��n�d{��$�Օ��_&��נ�07��7A�u�oqFۋ��/k�T���TT���F�zޓ��Ű�q�Ca�8<�^���fc��N��y�p?.�>ĀD����QvZȘ�0!�5{����՝�����)�?������㦒�i���P�f6�{^�gb,n�Z/�Ȭ��x�+��w��Ȯ;��rXZ#Y��'�2���Zu�Rie,�n7�8�c��=6�U0[�#�� �Sk�����D>3w8�y	Q��^p��Fu�^�������
���x�����`�UQ��ǐGf�q��N�j��J��K�/�cD)W�Խ������
k��!���~��|1�!�hjG�E.'��թ�6~�P����2��w귀���O���RgKe�}֧WH}"��z���T	�=\�`�Z߸�#acd �v���\�(hϬ��ǵ!;��^t�^��x��Nv�WhN��мk�Rͳ�y�p�^�x�Az�S'�:!��ĺ��U{����z	�)�7�!@?.]�#�lOpP�&�xe�ͲNȉ��4�s��`5:X�v�%�~lo7�h�Ư�����_v����5�0��9@�y��Q���ߣɋnU$�On�ц#����qnW)��i��.�?6-�SI.I?A��>{z a90�f�v�<��W��A�ך�=�}![�ty ��D<��_����Y7������w^8���։dQM���A������!h�]��xH�����⃡�� ����$IA]9=�)��x�Z��K��e̞b�K�z�jU�4GjQPK���#^6�<�>�l ����pX�Q�C�����fW���TO�0O4�����A@Q�/�*�,ӭ�V�B���/-�r�.y�Y"׸T1�|��_�/pl9����5��.]����m���b1kS��$��o2����D���^"Th2Fw[������<�y��]��%�_E�K��Z�T~��uΓ�pQn+$��gtt#`�,#t۽�����M�u��+��i;�.xmX�p���s�a��@P�dm���G�e��*��r�r֊Lh��,>Tq�XN9��½-�40ݣ<���1���=RٔIf������6}QO��n[��|�Dqȑv�e4KU*�|W�.���D��Td`EV����V)�����GG�}-�/�B��	99��/�s��P�K<�YG����d"Wi���=~�V�U����0~�`�Y��`�@����S��/�;T=���=^v��3��7\)��g�tR�L�DM�<ܑRj�$VL�P-�L����f�*yM�\������}���� i�p��QxB�eԅ����Ic��R߻N�U��+���X��� ��]��o.��$�&�S���)T��'���*�,�7��`G�2<!i�c�������g:7�`�s0Y�s��}�e6T��|ꧽp��bcs$��!ai�{����F����� �.�6!��6�#��T���D!t����z1�D�97m#��hS�O�.b�����iA�ʋ�V��!� �1��9��b#I�Ј⟺f��)�7e�Z����+3tSno�S(e[/� �X��/���`�}�җ~o����FH�SL{�Vİk3�ӝ6b%�KKc��"�l���j�J���� ��.=�ɑ� .�k�u&|�k���z`�O��eMˀ��Jl>���p��-��n(���a�Ѯ�^E	k�&\S�Vz��n��Q�]���H�O�(���xz�9g�������7�n��{�S-�%낓�l�6�����@ ��q�B�J�@8�v�@����(���_��+`fbfȝ�Lk�	��q_-G�՟Ȕe<��NS�`�.�Ź��-u�u e���mlp�b�������)��IV�}�i�B�~hu
�bl?Y�|�Iј
6?�/v"S�)�v�$�g���z���QD�E9ۡ����Z22.u#�~Z��up�22�?4~"|��7VVh�9=|o\z��źs���ʆ(�Z�і,c��?�PB	��rl�^��6VO,%�
�Usاs�t��f�������f�υq��U���n��E+���j�5S"��`�X2��
$8�$���OeJE6,G3����v�������������]���e����ӨMQ6�G��U�K�%��w��V�U�b�%��W�e
&��X"TX�����|�8d.��!G�w�/�m
������b�O�n�mTܭ���C'�v�	㶃Y��kM� {�t��k徺�ٜ��'�������mk}=��۸�X����3HG����L\B:_"܍�*���gP�;�~��������-�B5����͘��Ἔ�!�?��H���<�b�
r�1H�ٕi��U"^�SԘ�Z9�����d)^Μ�6���-�Đ�|��Q���4��8�ÜW�F���4%�ȥ�������rй�qXt��DM�� ��-0l�<�N|mK�	�-8Ֆrg`#�U�#0�(��zu��D���èA�U��:��E�H���@�3��T��<	�4$���]���5=h�o�A��z�d����}�<�ӇŖ)t 9Cݹ9�be�)T\[vX9���j{�B��w!����Y.��,��[�3�ߗ!��	ز۶m�6��e��8��CL��-һr��)1֊���#�^�8�,��R�䤟:�u �xZ��_<�"LR�5�A�!}UA����a�ɐ��$dK+3N�����Ʋ�H�4j��\`?�P������Dƥ��%��V֕���i`Ķ����4�"��,q��W��� ��$S5��<𾻟��<oh��9�ۅ�I�.֠�F�l����^b�D ߓv
L����s-�eN�4�ٙ}l���8'� ����X�+@2'l�����>@��9�pJp��`2���V�n�ʕi=-��SG��5/{�[�Q�c���F�(���[���I=���2;B%�ؓ)�3yzXG�3M	ڃ}�:�"�(7���S�T�(kXB���@��Q�l�����J��SJ�V\{琣�c|n�q�gXD��J�	�W���NÅ�g�O���.��W&?�F*ͅy����� z9�D=���LҡR�� ��gy	#�
=x�}bknS=�_�)a�������i��B� b���x���hK¹4w���s�8��HлV\�B�>�*f����� �ˌ��;�o�c�Xj��W��p�����֨���sa����M���&�r�H�fv�6Irnp2�iݜdJ�������,,z���
���X2�Rr���jUoc@�]̞������G�7���$����췧���&�ka�P\�e��<���}�> ����Rw8��.z�QP_Ⅳ�<��-�:;Ȼ��
�*�^	 �{�d�s���$�R��	ꮉ��UEV��7��5�"6:���|�`��yvE����z 7y��s��j�L�u*�m���b`h���F��g&CJ?["�sWp�`���ۈ���������ͽ�k�9��AB�A�+eG�T��
����-��H�=t����-f�؄��f�R�7�j�8s�����\�����W�Qe�񐄢S�"� �[��5��<�;����,�E� ���Y��������*_���o��[�iR	��>`7�~�`"��,K"u�_^�f�BJ��I�]4.�{h؜�.�H`�N��Sk��u����*䝚$r�H���
2V|��Y��� �-I�O�z��tb��/(4��D
�,��MfzB	�AY���	�5L�*�&����w�ڲlv#����Q�`�����������j���jgV��D���FV+��U�Zy�;$ ��\p��B���Sg (;�&�p�l�ɓ��>nB��S*^#��*C'��xƹߥ@�N
���<>ܘR����� �F���e#����P�����"�WI1#�N�3��%�� ⓲��+a��5��
x��s��NTt4+��R�4�;.��QҊȡd���C�IyQ�]��=����d�S<{����,&7i���m�J=5�/-���&R�9�<`�H��.3,�;������m���ߝ�|c/���E�����[��iR.������;v�.�2	�`&��q�]�3����?�L�5h�<f�8N�����Q�#�����3�+���&���?Th�{��0�Ͷ#K[B���V��'��+H��^�+T�����%�o��5~�Y�i[\�h5�A�2~@�?R%��4x�)�c��l�A���U/x�����ŋ�ᔤ�R�K������a���c�L{�PeD����AزL`9s��� ?qO7�y��b�Ң��T�#M�0�P�TE�A@k\�Y����:�E�����j�?��-t]u�:��.k��x�C5�F�w��v`�'��}$��ly��F�"x�t�P���YN��5�������ZZ^'��,l� �=Myi�9��SU�#��c��F>$dGb��-@F����Æh����Pӏ��AC�¼�E����$�G�bR�k�<�?Bn:˻'ۛ)ERd���ٶ�uwۯ������	v229���C�RBݤKF�vY�V*�<$}7򣞬pۛQ���^¶63ؗ�_*"s#(tg<m,[f��Jq;�!~n�f0=�Bu��c��m����M�ʈj�; �4�9g�~.�����x�pv�����C��Xe�O�c���3�D.+�X� '"B%�mD�#�?@̸/���}���}�ѓ�zP��ݞ�C�]�x�TDe��p��QAF�G�$Z!M��IE�:����ӑB��**��>��³�:�49�;'��rgA���U�Ĩ�{|��8����]����a9~oMsWd7 �TE`�<��6ksk���޼[�m��V~n���ju#˶Z,�ShsE���ZPP�̔o��4pQ�)�V��VPL6�lKO�2=&3�,��apx{e.4m�F~
����(���)��H,⑒ݿ0�}Peʓ7��+C�UK��{τ8��p��Sƫn?�~�X90/ �=��Ezҕ��e'Lh㟃a߬�V��P�b��߁4	��������E�i�W�N0��O��HV��*i�=ۡ�u��i�U*��?�x��x�#�$&X!!d���.11�Om��A^烩/ք92?�5��j��wL7W��E2�%�2�c��o��X9g\�G� �j�Zy�a��#&�xX��q|�~�,��hY�!��]�P�+�����3��ۂ��z��<V�xD�=߸��@��+�?�����|��FD����0���S_�|X9$-h�42hy�5
�I�W;Y	�J؟��!T�K�ry�����L�Id���~�����_1['Wo��'�֪"K��;vѡ�/8qX3�N�����s�`�8�����G�kFZ�ia����vt��
�v��N�/1=ȃuʐd�ҎΗC���9�6yq�Ő5M� pJ��.X5��
}�~�3'���x,���w̬/>�H��'O���,�p&3�PV0%,��\�#�S��N�y+��y^�Zn�Aa}_�xڧ���F��`���m��8��f�����""@u���@F��h��m�d�$��=�F�����n��X)k��z-��|���>��r�$�r�`@��hX���{"�j�p�r�ޣ�d%o�%���3E3�n����,F��X����G�C��!іr����r�����f%Z��b� �d�����Z7�A�.�q�C̴
�mǎZ	X�tcs ���'�r<��]��Z��$`�p��\m����Y�W`��w����2֢]�o����?�JT���x�I��k���PF��g��
9�ů�U.�ٛ���zB������q���\���ڎ&6{�P�W�X�Aw���$�h��+��N�S�u,�d�#5�/h�g;��}7�S�D�;0�O?�+\��]Zn�Q���!$Ij,��A��$L�V��1��������Ш]�-P�RB�Ν��sL�
��$KY��i�[�C=���W��Q�>B����J���Ꮃ�H��C̃/W�5ݕ^���`�!�H�f��A(l�%����-i��"E����U/AH��Z$�(Iג�JA��k[9a�B�a�STg�e�|��<�ї��=��}�.������8����)��&��p�QBgX.q�m�4�����F�˪1������~)����R���5	�Pޱ���<hҩ�\ӑq�����EbL�ҙߓ3I{M����R>.�'Wτ{�r��B͇�GQU�[��x�TW[����G�@��첢9�H$K@��k��-��w�^Q$�7�|X5�Ȭu.ҧv/���1Bq��Hde�{���b�u�_��YA!��P�r�1͘�ک�!G���o�F��@9ȭ�/a�6"�/5��sGŰ�}����+H�2w�Cr�/ʇ���Q6�;��ʺ�o����lÉj��t{�-]�
YNRo�,�*-ҕ� ��-�LO��H�V���^%��җ@CB��UO��$����1Lpԉ��'�Yf�Zֺ���41%u�ڒm��Ki*r����B���Q��ʁeAh�������h�����-A��c���`��5�*O�AD|f���u6iB(���wZ�|��C�?j�i�0/���0�Y�����@�L�w���j��H>���S6��E#>��Jp���_�����A�)=M�H��gpb@��<�[=+��^.yc�&��̆���O%��f�����Ě%�a�	\csx���3�撞��J84m�9/�u֛N	a}��z6I��VR��q]�g�(�-md1!��c�Uz�O�o.ߒj�0Lz�::���Y�����b����w�*�q_���R(�h��Ih~��2*\�-24&-���GlV���6c=�7�ש���Ps*S@4qj�Ob�&����m -zr�����a��O|W�M'ה]��;s��#���k&�����AeY�D�e����M�ߩkj<�]
M>Y���uda�fgUbcʪ��a��3�$!�(�k,$)�a;�����4���Ki3��R҃͝I�����}�h�lc���oH�2ϔ���B?���h�o%h���Ā\�$��p�ˤ�ױ�v�_=�8�L(A��8 ���*5�P��j�t��+U�>^.����D
8)�$+�p� �~D"�9�9W���n�<� ���������!)��B��
�}�M���u���ِU4�q}��=����Gy%ͅ��Hn��&MU�`z Owy�����0K��k���8��V̯���}
E>�~�>�n9���ŏlRv���-D�����@a�^a�B�b�5����x*���͞y���<\wӒ`�����.�m�("-��ыyR����6��vΠlx`h֮b�P����9$hD5$8b=��"ݕ��Q��ȑ���᰸F� 6��}����N4k�Q��2`�}�J���y���ξAh9I�T��%�j��,��Қ��_��>e��N��4�����t�ݔ�O���kX��iT�<��7�(2�*e'n׾��oI�M��s�v#�>*�a�DFѾ�u|� ^W�>/Ň��~wu��}c!�������L$��A<��_���.T�MR	Z�+{��[r���O�}�*�����W�x��C��n�xn�$��"�� ���.!B{�M�E� ~Vk�ymN�-DW:�?��q��u�z������k �]�ŭ��ȯ�ܡl1.,�)0��f�ꚁ<�� =��}:�M6OP;�-/�z���A�'���A���'���4�y\��G���Ld��,��m��$�T�]�9�S]��ґA1�W��-�^�k�BIr��p��S��x8q�.����(-|�u�޲��Ȁe1�a}��{���$�Q�#�z�;�����X)���)a��y5�ޣt��0�pª�������