��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J��R��g�p3����Apǜ��p�~��!�XZ�1 ��z���dl��Ѿc՗{����
5�H��=/{�bi�Æ���4��㊢���W��rzBћ);C֦x�&��O�@� j�;E���`l�h�[DIaģ��0r]�M��m��_[Lc���>��4�AZ�uN�Bn�TSh����/��w�T�ZKL�jE�C�@#1���kE� Rfw�&t�Y�0�^i�9�)��5��9��g�$��/�<���������s��aT�>�If�{�!�}q���/��f��!�ߨ�.�\.R�W�nU���Jͱ]�-����-Wn~�3�U]�AT�mtOۨ��@k���U,�U^s*��n̜���}:{�3*Iro�#�q��|ˌ*��^p$��Ȅ׬ �f_`��S�޹�"�K�u�X@y���1�h�m��VY]��{��Z�� 0����	��MH>���`���L��&��^}U�v�pj &�E��!�0��>�}�'��t�n+	���&Ɤ��gѳ����W�t��8)�tȚ��Z.�`���w+�S����,~�_�-(�M��E퍻�`措���IԊ��΅��R��g͆\=��O�l�3��"$~I�Bt|���c2k�b!�|���J�Gc��� 2	:����U%��&C�'���k[�^3㤃3����c���
�8ltQa�R�������5&�=���K̽(�`k���n`u;�\K��!sZ�Q1�@4��5r� y2dfR�;H���犴�f,�@����ãZ��V�����5P�&f�S�M�6s.L�9�����:໾�tq����HW��w��Wꨝ�~F���(�_>�u��7ʇ�2(K��u�*���6�~0�"�ӡU��@�Uދ������P���dh6�kBU��bT��ӳOs���n�c��{�@ƭ�� `�*�����>�yA%*+�lu��3�b�+^�9�%:Gv�MQ�T�Ɍ��Sƣڳ(�Q���?�|��h�#��7�M?r��KJ�O��^j;�P��Ύ���b�H�f�m��y�"	�����xy���wŎ{��}c8l��$[Ƅ�e���7��1���TITG���WKkhˣ_���ã�q*s}�p�5�^9İ�U����\�Ęx�8i�_M ��%��@\9�O�U�j9��M=�v$��]3�K[B�){��v�0I]�D��ݥ��OmMd�)��a�|zL~S��cX?W����B�!HW�w�'�?��pz̀�]�i���x��cn]Y�I�=�T/���hD�u�M�u��*��̛X�x�NM�����Q�<�6L�8��~�|��4Ʉ��Q�Bs�<x�kaR-�����o�Wp-�*�,��u������/��~����^����{y!�6wx����L�0x pƂ�(�48ķ$mM���k�\h�p
ߍ6�`'�#�k�1�_[!;��h�5;u������)>���y����f�8[-r��|�*V�M�~UV�\��Q�U�Zi��E��^�YR���s��cn�Y6İa�(*p�D�/Š�)�R~9Һi�	X٢ѴxI����j��E)�%������a`R�::�z&��=}�=5�U���0#��T�M���I;eM��4��b��8���-�U��Ta�,���j�m8{R�k��#j7�	�,(zA6�r8s��/� |E��Ün������}����ag�ёITo���s�
������]�zYC�+k�-����L�p6����(.q
}�݃3v��-wf����ϚY�D��:5��Y��$����J�#!�kR\縷!�HQ/���E�X�fp��<N�$3:x�C�C��G���6��d���[�0���"%�c5�A褑"�-�P��Y���HP�1ŗ�]��~����X��C��]�c��ˮ1���݃D�\ِ~��x`.U�:�Qo��itM'HJ$B�u�(���n�������R�;ǀ�cZ������ak2������,�؆�1�oy�"R4�v�Q�]�Ƈ^�h9���"��lu��+��Ky؞,��+&{�^�E�q瓏pr_/�p���"�0}��@�%����ȟ
��&�#� <t�e�Aè����@���K4�h�ECn��+\�I?x��?��[[M=]`���2�Jͩ9�����y���a�h�EꟂZ:�CES'Y��8��� �`���5:FF.E�#�c��8j��i�Dv�kA��Q+�HM�i���p�6�X���{Rۯ����:���,.OA��^'Y-+ꈪ��S[HJ�$�����x��5Γ���'�ElF��N�:`X|�>"��C%�:�k�e�N?"������tA� 5���^����G���W=��g&��u`ZV�މ�i02W�yPhEB��	�Ee#��Fl��p���8�`M7���E�Z�159+)������4.����7��?�������­`*����?}
:�٨��\�̒E��9/�n<��㷥'f;��[CC�m/M�H�Z�Yi���ߩ7��B�v�OB��M��'�0�Ԍd�k�΃�;�aR��u�b��Zh7Y�0-��T�  G���&�Y����Ҹ4&��eg�6��K��"�3%�h�Tǵ!
!�+��<�[��w���� S����"�F6�&�\l��v���Q�4(�^C;��RC	:�.!�M��y��|�q>���	�B����C�_��R��=_�r
�]B�	�0z�S)H($�G<ϼĥ]��/�~`L� ��2%q��HIo��!#xT�ػ ab`��Ssճd�|�h�o��	I����
�������c�Ţ\,����i�:��d�uN�vol��M�x`�mf֯٦�y��=C�ؠ��
����� �6�	�F�0�U.�#�e��;�z�Y�Z5&_�S4)�(b��\%�D�n�r��ծ]�v�W$W!�_��a��}�g�>�s������(�^x9��>����W�x`NON@�1;˰#»>���@w��� {�Ҁ����|����D2/���
g�ƖC/����62�p�H��8���Y��G��,4SS�L�Sj�E��-W�J������3�޺7lxF�#Ȍ�x���~(g�h�+��/畹�x$zz�gY�r�[��/����"ҹWI@rI�IK��Ā�G���9%M�4T��Os6��:��,j	���iL8�dlMZTq�(i��a֩��Ӵ�P3#��OP�L���D�y��4����6<l��dze�M"�K<#`?�2LB���Ψ#m\b�JY�M����jW�&�&�k��=�8�-Ž,N]9TI	��jy��[��=��׼�я+m+��0��A����=Za��-o x��0>�0���S4M8��~<L����\��#À��H<DL*C�������(=�����9�㴿(m��B!~xR��]�%���Et��!/Td�´6��uxF/c���<g�l�W��?����.2T������H?+�O(�Jqދ��1�M+��e�$���v��������\�hr�]v��n��f���C�;���l�ݻ�y�M��r��a4mQ��A�[�T����ڝ�@�"#T�%hO���eSV����x�4�:V3 �'4����ǽ_#�CQ����p��,M�UY���dG�ЛLs5���Gk��X'�:��?4�D�J�^��e1};!B���:0b�!���:y��4��"���<�bC�z�{�N�)%1i����
�Ѥс���.�E��"+I�� q�-���vȾ�i���7��	}5��r@����A���L�*�ʶf�"m{4ז��L�O� F=�W�:A�eV�<�D��WpJÞ|��&�l�P����7`�SI�ϕ�Mf�J��N�n�Ӫ�q�4�Q�B �]�=�33י��|���W�dN,��'zѲ)�h�ץkQ&sD"�I���` �`�[ق��&}K�S����wE�_�g�?x)4���C޾hII�c/9!֜bϭ��8W�Km
n��Bk4�(�:�����`���9��f4+^W]�~�uW�(�J�E�ڐ�P��QnA�#��h�~�Ak�	����2�r�^;Q4քin�i��J�����9eC�}ݗs�s'v�?8��Anp'�6}��֨��,��c���b$�>��"�>�
�ܴͨq��ӻ�q��s0�q��c˚����k�lwL!V�sA���&�V�S��+w!�+�J?<��Ӑ3���Ǆ��⁢,��`�C���dD*�&U,�0)�S�̲w
���u����	�/��(ϵ�_�`�2���Ԙw98���u����=�8�DoS�gؼ�y�d4S�<Y|T2cg]{�BƛRWǢ��J�h�D �V�B�yu-k!`��Hq%8+����`�ަ+��W�ˠ}�3��)��8a?���!҈�Q��)I� p�j%b���o��-��H�Xiaw����jk�r��_�9����ʊu8$��H2~�w_ܩp�swZx���92����Vݪ0.��~]S��ov�J������:(Ǡ[dM�V�	��*�p�����,Ì�ϯK6id�[�&k�g:�
���p���X�bK���_s�s{��j�p�'��RBKGqH�sBj�q���n��ɀ�/�*܎!�D��2uH���GQ/D��نw���6&;�
��٘E{HcjI�
g\z!�,9�rh3�cR�ìN�hUh�d����ݛ�|�8(�fx��F}%>�;���˕�e���ߞ����fk-^�v ��l�d/C�b��U�v����bES�c^96��s��)YtT��P�l�Sr����~A[yh��f84)y8� >����(l 5�as�+z��B. -��ѫ��5Ҭ����K���6gqz�9�r�����ٽ(���	!���pS����H�x���<9�JW��m{rDi�_,����Uߋ�-^Y��6�45O+��zKf1����`N#�_��ei�,���OX%�FtV��I�m�@>x��1ݤ��St�͙Vֹ,�����Q����� �+�f,��Nʯی��ֽ���f�$�� 6����@G$�/�fԾ�5{&Վ7��5��3*�Nj��.2���g�>��X�O�ۆv{���<�o�L�.E����ԏ�5\R{�����Q�b��J�0���c-�i��L�nG���q�!M��21��0͑r��+8l^?�x����BS$��I�΍�j�� 7�R;^U�)�p�%m�Z��("!WvYe�3����{�α��bpb�����)�a>��i��*�~����Q�c��۠Te�fׇ��J�7����I�_1�U�TB���t�&���u!�MI��&�yk�g��������VR���*����>��3������V��f�N���6��i��{���� Z�U''�j�i`>��q[�z�&5k����N�i�b/OΑ��=,�ߞ+3��#����!�Xκ<ϯ�� �ߵ�éʴd�X}��.˜�T�W߇uY2���/��(D�x�K�`��mp�������fט��(}ޒw!�*])����� ��wpC\�o�_Gx�{�lo>�ن�&�̛�*�o�oe�|�_>���ikJ<f��>�����2B���hn�mnx��S��z�!4�A��y�VJ���c���O8���&)��H�-���%�VЫ����J�+l^^��7�w���^�|�a��T�F;�v{]7�|��o��}m-�?W1n�tZ�Y��F��6)�慐jv*sJ�)�������#��|{�{_�n���uh2�@�s9�����7<Q��.��!��ӥzX@��X�.���`x�.��0�T���#�����ю�j���b���&�f���q �qX|VVv�l8�BGB1)����Ł�jh�M|d|�B��>�S�iLS�l���PNWG#���8�t�}�,#�[N�b?��ȯ����}S&a������,�c+��M#U2�}����ʔ���_�O*n�^q���p,?�i3��(��$��[��t�]��#��b�d�V��҆�7��l��h�J��p�;~�o�7�(���?���y��A���U�"+��\��3���f����OD��,R���x+��=�B�`�?v��#�>�܃h��ľ�.O�2��统�"�e��6�S���)xGJ1b�����>W�:XYj�N��E�jF��h�_C����3�5��in´	����E�T-������-?��J�I�l=��ۚ7:����5���X����,j���f�]��go�1�\ZPy)��z����*;b����sꟹ�z�!��~luO W��m(ۤ�д���npwZ��/��m�ݨ1IS�x0�!r�J���Mʔ��n}g';]v2ܺ٬ �ck��!9aՀ�Hh�S{���<G⻴���:���y�	!���L�-T1w-DPR-�Dl2#�Q	/h������q �ա�� aT�ׄ{������L%e���4�[	"�Z����;$�6Y[z.yܲ��,���<u3/n��0�Z3 J?M�{��ǽRV����n���x�)s�o��+��
�Z�B.|���\�E.|���	o ���z��W72B:`�Uꏽ]����DD�I�"}@1G�!g���ҵη�R�#B�|���7-�C�n�H�`j[�z��$�bZ-���칰*�Z4ug�Q�D<�-tq��a &%S�'�-!���2�������y3�M'���*4"��&"�C�#Xq����z�ɾ�oӕ���H��U�v��/}à����£��yd�t��%F/�<�Y�5��8�����U�Ҫ�`-��}���PKE�ҫ^�	�[�j�+e��̢�����#'��U�~��j��zc��Gt
'E�(^�n�-�$�m��j
��O�wy��(<���]�˶)�)���O��fa�h�T�m�����o���(�y�v�_�p}��[6�QL�&8-�N����mx��{UP#�i�� ��$-o�l�����G��{��ߪ���I^^��3-e{&�m�5�QZ����U�5���;?��p>O����|���L�򜰩�~�j	?>]1ƘfB;����~��Yj�xA��k��?����L[�&H7�M&$B�D��R�0}���c��A��� �O�H�|u,�eyY�<�1|�������2�zrG��oKXe/3̐�p��B�CQ�S��v{�h�ySv�X�;������V�|�zβ�4oT����iȝ�i���E16G����˯��|����E�������>��e�ϣp�U���4kE��"a���/�}� ��?��ŲQ�b�K+>A��7�����Bu��'���ΈD�_� p�b��K��>�a?/��@�X���)���B��>�����,H��v��2FiTx�]��r�*�W����H[^Of�!��
�����ril���9���"��XAz	[��2�{�H@ ����45��4 7x����I��i+λ&'Z2y/���W����_`O��>����pƿ�i	��"h3�����҈8����4.,Hg��������Gl�p����o�W^��Q깱��:��^~A�΁��@MREx?�_�q�m�̢=��9�|�]RƲ�a����n����2`
(&IQ)KQ���o�O���KuV?Ũ�\��<��f������rC1��ﭻ���+|��v��	�\��{}-|z�e$���rE��NFPf#��B	����?~�޳?�Џ\�n´@M��2��5�cH��k��)���@����IH�z�!ݵ�$đ�@2c�
-�1.�{l5�h�t(��)ӢJB��t-�b#O����bڗխ����߷L�&rs,� -It�_�ؑ��)���â�|AěB�h!��6�o��k��0���'��Y�k����A}��w���	�ڸQ�a��Ibqy3h)�?2Qom�����5/�kh����/S�֬�(�ב����r;�rX��"����O��W��)4�V��{�3y�^_���NCH�U�D�=6�u��:���&vt����V�� ����������1U�z��=��-Rfp�t������=��-���Q/t\sS��D�~E$�s6x0�Z�������V6!�a���W���t�m��T:j-� L�S��&i�^�0<�UK�8��B{�z;U�Dcl��sV���k�x�yf��I�-��N�Bˎ޸iyaS�ŉiS%��I�� �s8����}����u�*$>j6e����JM�
�4����z��~W.8-�;?�哄����Eh�+��ܗ�Pi����m����7
Je�����(�d�;���ub��h[7q ���g��*��6�AP���Z��*`���|�繳���d�n�p�T��3Iz�K��{�,"O�Z�(��|�H�?b�A)+��Q�m��	)�,�KkY���0W�v���\8	uZ
�̌�p�_��i��ڟBD+=�a����G�<�8CY�-���H5\��H�fHP�u3�-���1X� �<��L�*Jי�%Ma�G��u�R���1	�!]RUlb8�%N��H?3'�bG�ѭ%�2�ۡ �r�hq>P�oY�HZe�<j��
 ����F�����"���U�)��*���)+'j�.���%�-����B�B��p ��B��V���YZ1-��[�e�5z�	���5ac��rXI���}���|��H���]W;�S�	j��&gA�0$��f�u�At �Yfx���%R�����]{��}z�,�O����J�
�Dj��PW{��L���6�d��i���~}��\kFs0�c%f�nI��zŦ��*�!ׇ.�ʸ�C	E�r6f��Y���xSsNE�� ��j[�q�zC�w˅�r�½ԤR"�}c��`�ȸU��Cb�v����f+�p|�`�m,Ǫo��� 9�VA���x�!F�vI)�l<n"s��g3{gOø�ƞ|���V�4#]�Y <N�1�n�T>Ș>D!�f�S�c�?�+j�dd	��e��D�C����Bw��r ���=$�Q_a�L�u�y51�%�=.����ޢq���G��ɝ�����J)�%�3g�I���
P�8�Y6	�n�[D.3�U��}�!�	^�v�s�
��3&���{\��0�8elցD��+�O��L�G��?,�PP)]����V�濉X:�e�E�Z�q��D�c.����s
���QϾ�g%�v��&��1c��J}\��V�� -�&V��lk��8C��Ӗa4^㶽����6�!��� \�V�2�Kv���t�t-��3��ъ��d���ը��E�{��Y#0�$���sbQ�ф"�7|�<!��Ъ�bf-oQ>�'���L�a��$�#*+&C�Kz/�vV��?��O�,�����U�E��N�Y���PKl��Ak�a��q���x����l&��b�m �1�$?g���w��6R6��Q������X�)����O�?�SB��6�B�X�q���$ɀ�wT����~��r�:���pY88�IH=}O�7_F4�KY��;W�R- ��� #��7��Q��,�ïH.k]8�3b�s	�����o��O7��ݬ�9w�	�,ξ �}�r��L�Ԥ`<��������;H$e����`�a�A�����'Y_�)�VdK�C��S,� %�(�NZ�°ԊD���DLd̵߉]-�k%K��Q�4�K�U�$�3t%��]A�����q�5��@?��"ܲ� r�!!��Z����
p*��nBۦ�tX�b�8��	�"`~v8<2�f��I[ ���;�L�Ӛd���%�<N��o�Y��z8G������81�<�g��ѳ�M���#��$)�nw�n�]R�t/0���_�N�%x�:����&C�G��W�����E�8��͟�C�q����A�Q�G�$�*���gҦbE���Ϯ&�5%Z,�8�O�&��r.q�?��#X�&R����О� �Z"�׬���_
Ug����f]�Y����$�N�k_w�;�5��ʌ*8�H6�i�F���I���^���X��߷�-c�h�[7�f�A�Z����u�x���@$ќ�R��?�g�ѴCf�r8����{�����	���<�E���Rqyf�1s�7��?�#�B6��d=�U��h�l�����˛�x�s��o�����X�Q���cٽ�<8	6,{��S�G(]�.�|
#����)�Z��C�Qb�P��s�'S�ё��E�nE�a���Y4���K%���'Y6VB~���g�Z�	�0�ݥ4$k�6��9��"��Հ�dPXM%���g1��43XM��a㋿��U���?{�$X��׎2��5���'6-�x�N7�"��8%K���3D��_�<�?u*�}�<2�������(�����٭/ �v��U�j��a����a��H��~c{�M�>b+J&��-)_Ƣ	�����%h�lvwwX5���9��z��N�v9�6H�V^w��X�B����YV�WĻ��t&��t�TS����N|u�����Hn���v���^]�5K]H�̨�黒�8{=i2%�7�Zm�[���X�*;T��[�X�Z��Ճ�,P�����e��Rm���˻mU�uW��Ѿ.�x�k�?����^�u�;���[��̈́{�ذ^��x�O�g+.u�� Tv�����ѐ/�Z�áN���9����vZC+�a<�0�T�1`J��&�@�v����)����:��҉�2w��#l'N�X�$(��z�A3	{���c�6W���2�\����kv��'�8���`��*"'�/�ӑ�B��̘O�1`c��=�� v�"K��Iᶿ�����"�l��Um��U%ϸ{�'E�ac2���94�*��n�D�������KU�[::��i�Z@6�G�a�uR��j����ԖP�C`��<��f`������e�����rY[��!Ȯ�� �;*��bx`�x��B��OZ1�?�<P&�9"�pU�.�ʩ�Q���-�=��񊖰��� 0�I��ʄ���pfOe��Kh����h�%�v3����}���g��#/����Ե3�l���ʮp�/�
���_�Nߏ�;`�S�賙�gݏ��g�I>����zU�`8O2�P���z����KQT�-@'�M�]��6a�E�`���wT?�����k9!з#V��/(`���<���e���=�e�l���h�'s���r���yߒh+_�t,���r���6�ՉET�Rp(�N�c{O*�G�Y�U��m;���b�����h���Jʫ�q�J����Xa�����|`�zvE㪔@I2�<�w�<����T��0�
<���T�	v$�f�G�#���:���6U�k�l���0�1�L�=�|q&	t�Q�'V0�� u�l6E�����V��0�b�b,��:
j��sL���;c��vS��U�ՂbG�`��g���&#����f����NU���ߑo��숇H�ڄq)]|��/#Ζ� }�D\�y%���)��_7�G�n\9���G�\�31���.�]�2	���\t������2 �ŭ���6;��<8���:3�7Ww�&��?����<&9:��X����r�"���PL�Zo��iB�??���_Nx�Ez�_�#%�J��&\@��=��'��ИK+�A�k�l��cT�����9����5ݢ�w"���^��Vsr2F�����;5������wN2~�Ŏ<d��^Vf�Y����v��$�B@&��qN�
D;1���/MU�8t;q���lm�����e�P��E�;�=�~�� ��m�A^ƫ��������'%��g!9��Ril��0�c�3l�|3��*]�l��CяA#���M���l|N��4��oD���f�L�d���Yrj0��b|t4��r�܄�!Q ���m�/���*��mA�
q�4�W��WS�;���	�+8*,@A>Y���gM|���#�o2��u6�$Q�j��Z�ͅ^�]g�?{�b��E{oS�����u���oΧ_���-H�kU�H:��@�ns,�yq�8Q2)�+,SF=V�p=*��!� d��Z`�Q��=�x��w��Z�*a���|U�%,�[�����e�*锳�QM���1R
ԑP#�q�B�m��d-g��֢�������t�3�+����8�:@N2��LN�$垐�s^�(�� χ'�.~,�痰�C��H�ٝ��1w�q8��"��Gp2)�����%�
��]�:���}r1)��������}_��}g���F�Kjޫ�+l�Ql�s◽�y%��*e�G���ϙ�<�N���x?X��6HU�v���+[���i,O�(n������j�E}�r���l���_�(��w�c-�I�휩h�=T'P��1��ۧ��&(��}�� D5���Ī��)�k�^�"���C&�f�� �Y-�uv�H_#<� �%#��&T`Q{g0�'8o��oaH>ڇ�
�v����%X��B_i��1u�0��WU��ׄ6�o�;�{�8:_���g�E���B�8���s��@��Ǵ@?��oh/��(T]�b�������e�?�\3.O��G*i�U��'l��+��ᚈ7�`���G�~Х� $�B�Qg�$� L���o!�P���3R}�Wz`�b1�٦�,���t'd�bZ��n��Ro�.�vC.��)F^0�L�2&"�;����V�m�=�z��J��ͬ�mC����&y9�K���È_��KQ@����L>rU��[�z�?&�О���F��>"+t��X���X8��nX�
���0O�̊+۪�-�,������� �Uن�sK�����F�kh�1XG����H��e\���-T&1$��ޗ/��A�~�y?�A=��]k��V����sb'��l��ʃ'-�0!��/�|��@ډ��2����4y{�YW�����/RJ�*���ݭ�B��� �P0��<κ��G����г|��8A3mYZ�?�L(��p,x;f��7��'��!;��z�Ko%�b�����m�8iN�^Z�\-�p����(3\�̐>�Y�2N¬�&�?!�?����D��Q"ߎ���^�M�B��E����p$\p�bg�Z��D�,����`��G��Q�3�M0P?������%����gqB8��Ր3�b7@U�Z�7j���6�����I�x�����͌���=�8��K�BeΞ�:�e	g>7\)�+]�Sl�[�㎽�IXU��lh��3O��6\������(��K^���rpm?�?sE�Me�{\��hjl/=�w8�"&� ��1Rz�wӪi�`�M%c �!�޴V�(ng��!!�����$)_d���>b��n�	��',�%�?�i�A�B�~7��j�#y�&�	�q���c��o�>�dє����	niH�UJ�Y,r>ޜԶ���?���ar�k�j��y�9/�w!�?��oB���_���YZ�"|K�Xr��W� �t�y	�"F�(H�� H�O1�M�oc)ow��3��� ��m�AO$�C�@�s���� ����s�E_�Cg�cO2�:�&8}��G����MGz�t��*�O�w���FZ�(2V�z��5��u�42�����ye4�`�}*�+�!��B��S�##�Y��t�9��%}S��`�C���=�\��C3cu�!6��@����:��Mt�rD�i���!	5�֊�+�E}u=�
�!<~FAjn��a���-ކ(��vj��uI9��.!��&�+��Cj �\1>�8�	�G�ڸ�R5W���Y��O�Lu�Ԭ�����v����PO3xO%���b�}�g���E�P����jЇr�ؾ�������{�#hw�&����	�qa,���Dj��f��v)7[�v>�I�La��M���n8<));�����O-�xE8vSZ��syt�s"�����7h�1,�R�����W_���Jڭ����JN�%{�;8��Kyp%LSA�;�,4H�:j{��a��p��ϬṯcA��]�{�r���ag����-޸�V�r�`IC�&�|�m���d��#�?�T��p��/����D��<��m&��bg��N(�P�zsGԧ�7U�;�/��\}����F��?���n)
����w:)떃�EX }.<��ĉ&fY�&^8N#��8q��I:�+��b"	^�P��߹G����ỗ�]du�?b��\͐+`_��ڐ�|ZJ�X�y��% �o���l# �:����}�򐋮c(��ث�A�k����<�q9�:�����ot¥��
��s}�dȷK�߇�[�6�­��B�~p���X6�m�@F-�A���B�u:�>��b� ��I�2�V��@8:%�C��Xr�����=��J����.U�q�G�.7rm:bp������u���f�(�j�1������!`,G���+#�s����1�4�}�����9|6:W2U��=1�D��6t��D.��V�n���#^��h��&؇��2�X��ܥ��@�x�m�e�r���>�2Ne�prTP��(�s7ot97��\�c'�����^��RC��Z���t�O�t�Hk�ԡ�)ύ��j\��͑��_�c�W�-3��(��/�Z����a��f�-��1��%?9Z��^T�2�s�O�#);�\"NZr���Ȏ*(H�"�������� *�&Λ����k�Û�$�������/R9��٘?#}��7���R�sb�t0lE��F�,"L��XZ��KS� )A�@���x�#����d�*���'�~	b�M	��|�Ŧ�
y�'`kq*�*��~/��/a�"��$8Z��I-g���ׅoû�*�(߅�Gm�ݠߤu�p*0�E�I��2��zG&8ܓ�����-b^,��#�������l����
�0iCz�T�ľ�������^iQ.�-`j�w!�G�}N\����+���'�CK���WU��l����^�4΂ܔ&����:o�mf�-'T�����������JsTJd7t�jkb�$۽ڟ�y0��Eљ����~E�?�FSIk쫣Ҡ�kH��]�+=җGvr�K���ߒ1�A>F���������Km��1z��]�z��{1�L�9��k��DD�'����Cy��i; ���A��g�G�4�F-Iw
�_U�����tdm�Ÿx�/$�#�Z��	�[�}}�dS�<�18��:��� ۀ���j-o[�IiD&��̃�dUe_��ƕitG�}<��E�Y�]�yD�R�����T����§śn�\_����u�;��L��5�ȼ<��_8�rE��+��,�E�`T����Ɇ�s��6:�.Mt�<r:Աi�Y
��|�����Vr��ķ�д�y��\1��}L�
O��`��'����J.��
G^n.�hI/���_�l���0LՓD���*�.�&X�U�~�B�<��z�#�`w��I��\�)���ʓ+x��������>kA3Di��灛�"9�}�Qە�g���f4-	�n��zV���퓚p�k^��_�A$��0��d���"a�%�f���	\��ȭ�_I���~��fC�V�������=)LE�*�W7��b@4���T���W4�s:��c��F�)aQ��N��m
�?z�����F�2VS��(Z�L�y����ͼ��g������:�i�lc�٦׹����t쐺2��&xv���B���m����k5��]��� ���{z��ƛ\?*"4b��]&?�q]	���ظ?�@�F�}�-R:���ѧ9Ц�xg��D����X1�5�[��u� h�}9�Z)�+!� "D`U��,2]=��Iq�o�9��[��B�����q���ЉZggSN*�Q��N?�x4��hW�e L�
J�Udm(�RO
��h�����_����r=ɴ��B$@d!a�Pt'<���-q�uU�F�z.�0��: �l�+g�����"�1�d;t�q���"��TY��=\>=����=^�C��ζh(O�/�΄�R�uR��zd��n�,>4˶���П��A6N�87k�������3`���SCeyʍ�E O��!ԋ��.�Y�'Eq��($��/ut��7�;~�\�N 򪪦Ya�1�zn������yt���������.}wh
}AN�UH��>q�q�iᨗ\�B��'s�?�=�h>_I�KH=t~�駊�'�t��)�)Ϡ��xQP��}�����`N��*Q���q�C�A%<G���~���3sq"G4_G1f�������9i���!�D��u�:�rW,(9A�|&���5�m���L�Voᗚ:��DiѾ��b)u��W�0K��Hc����`�W}V��u'	.�`F���M8kH�#�W�iv��Ǡ�U.K�J?l��� ��[K^L�Ԩ�͞$7�1'�y�9Y�l�э�8�ӛ�?xi�4������&����%���S͉#�T���U~_������w��}���04f�� ��q06�53M��8I�vqφ��-�d�KX�{�
�fꟌ֎u�
Ռ1f�+��M%��%?���>���	| �mF!����k?`�З�"�Wq���ɼ#M�D�듈��EP�;�L�Y��[��X2p)�����6�.\�I/��f^��.��(:"Y)��3=�~}THK1aq��Э�\-ѧE��6�]�M�r�~��lJ5z�c�Զ�d2B������%�L%S�@�C�j�5�Y+d�zu�>�d�������o��R�ԧB��դ� ����z��w$����-��I؂K'��4;-_+)A�2.Om�pc<��b-g��#���ا��A���E�o.����]]b�"�=�L�K��pj�L!���X>�Ӝ|a�l��뿆 ZA�;�N�o�H ������m����pUt.DI��� ��t��:V�?�DAi�d���aN��\�`�Y�r��nY��{��m���L`"��~��6��Nexb��ST_NN0C���/L��.��2t���R��F9�Q�̱1�Ԯ�3�H��ːb#r��l�=�QT߱�X�Z�/"�|$�X%�L0녷�[�հ�IdP�]� ���<%A=!-Z�]#�=|qR�%)֫�����䁠	P��� �9\�+l��/ҕr���$��3���:Hh7���gp`T��8�)M��E��I*|�,pW�	�2�`�yt�Ӆp�yGc}��_=o5�:��ߔ��$�@�氂��;��_괄�g���S*���34�����qvm3
�6Sְ,����a>e���p7�+KY���j�����y�����}i?��>��hq�D�R�����5����;�=��j/���i6�(���#,�CRd�Iժ2����ȡ��$��C��@�EnԿ������PRaؚ:�ߺ�X�9���~c���+��,�@sU��{�)�u~k}�
/TW7j�F�c��r��loG��K:���*�i����Q���o��L�lNO��f�������`�շ�1�U4
x]XH�[	X�B�D�~���-�E���k4w.�A���.%(��
L{�85�2{b�jN��5��mw~޵$�edV����Ad�Rý���G��ֻ���]���j����2���tL9O�4�s�W�5��z���P�&\��PH]ͩ���օ��x�z�'��#@L�����������O�����O���N�*#0a�-��NBI]����r��5�H�w�ej�k��~��?�9J��z,�����9\n�����I��X�y,�W����$��lU#we���S�Щ����O��Ӎ̊��� @�*�6�P܂�}�6����ic��2�ç��J��S��{7���kGA��*�l��XJC�\hT4^^�����V632;����C%�/�Z?�y�'�X�uPx����l�M�j�����@���
V	qM���y
�MҩHV�.��9Qr���Z��x(�נ^�iiї�O�	Ϧ�� ��K�Zi��F���7�n��7���)���Z���'m�}�Õ�@!�i*6@IT'{���O��d�=��U��=(���M�~��^�e`=�>��c���mn
��Q�:!��<J��Y�N�!B��'��P�B����}�7:Z{������E�����xR�5�Z�3���s�D�(��4�P�yn��ohz�{$8�0�@[ϙ#%�_�NȾ#V���@HE�	|����z���� Ḣ8MIB�R��
��C��v�-ݴ�z�+D�[�x�_�i �Ԣ&���O�k<G����+q>�p@�X|��7�y�Ǩ���rgZK�(e��S��E�6���Jj�j|��O�;���V�6����t'W��5��7�yn����V!f�+0poi{V$��2-�R���_0�N�@+ڃ��kޛ����*e8Im2a��M���U'��n�	#ذJ{K\r����M����1�S_/X����R���Z!�>s�9T����6��m���+����q2�\_��I���5~��[�\�3%́�x�9�O���T4�1�t���z���:�!J<\�M���gA_@0�#�'�ᗵ�ׄ�h&ꅽM�����L.EV�٬���#C@7^'��S̰���ݟ,�ڸ�D�/�}0+&�Fd,�}H����E-B�$ͩ�5L���U�:�����Z.�TT�y.���ܭƎ�r����F�6��x����5�aآ�O��Ҭ��C��8ѻR��Wl�m��*cR*lB�	����$�i�YfF;�T��n��0�ѫe? {�[|]������_�1���L?��<�7b�t �d�rkr���B,D\7̀K�_�Ob��܇���>Nt7n/Āܳ�Yٻ,WjG�X�q_ʒ��ax���(�\&3C�*�"|�����U�y��D��@u���m���!��zO�
^��	�&D�qv_i �lm�ڲ�_Wph�?��i0x�R�	�?�c�?�Y\n��=o㚓����E��:�:E���y�m�N�C()>)��܆y�^_b��? w[�a�~��.�=`WV�d��S�������0�w�ү�r}��+����7jJU��;�*���!}��z�-�ËRbce#���L=y6��Y	-��"�4|q��ϐ���l��<eǶh5ǫ�̵�ۻ�
��6����R�x
�xq0[��=ֽ�(�t���RU�N�_⑔�SD�l�~$��U��6�\;�jQgJ�G8�<��;?#��c�5V��ӛ�����{q]��<�xXKZ�X���y}�x���`g�ۉ�����C�&E��&�/�ʁ��p�:ŉ*%���{H�� N���8�"c(^��F��oێ����u�4( �tԖ:c� �گ�rI75��wk�~2_�1J���nῘ"���<t���vo��� �ab���Mh߸M�iE�6d��B���]
z��yK�b"aEH��t< ���h|5֗� �{�s�Ƒ����̒R����,CB�y���E�63�A�J^���| �@�Z=0ݓ��iJ��m��O���]z�5�1� #Kz^ O)��G�io��*j�W�r�F�����z:��${�I��w�t�<I��!�K>�U���q�y�QҊ�quջ���*�>GE��ƫ�_'�&Zy��I3$W^�`��29���e��2�\4�Q\L�N�`��'8a�􎠗"4vTdz��␂���NB�&Tq����?߲/%F�.��V�o�*?M����E@�Sr�9��(;N���Q�j�H��!�Q8�Y���&,�A8�>�ٗ7T�N�9&~'V2w�4�T��`[�;�(s����'����Ţ�H�嶽�AFNn��=�RT3c5Sܭ�oN�3˾l�K�����S��.�B6�PQe���?Z��-�	O�[���b�JK�{�@ZT�:wg_ȉٯ*r��'/�\T	�f�"Sԏ
aD�
�0��%��Y�]��ț�ے4���d�����*�/��}1���Z���c���w����Da2��F����h��;2:����m���+ff�i:,�t�Yр�	�F,z���07�.��Ò�k����� �@֯�?��Fr�>�DC�yW�Q���8Plp
���wx̸�^lo.T�\��J8�$v��Z�Q�5������X���H���d�	zQ��g�?�ЀH���~��a�H����"Ě��R�h�4_���Nt�
OAx�M�p(��O�yqX�&Ie=gN����>���ϊq��J"hy����xZ�w��M$���c��x��q�FM�Ǉ���V�FsTx���3˿�`:������5�p��S�Vv��2T�F���_�p��t���G�F2��jL�̛�O��D��L�����ݤfbq��)��6��Q����n�M�f��dP66?AS��i�d	��Vτ�xe�k�E�v��(ޔ���+���F�r�w��\���Uc5,���>�􂜥�p��ˌp!�Lt�t*hf�/B־�{<o�[$�!w�1>bI&䶠[�d�������>B�D�� Fo<�����J���N;>q\��ᆂ��A�T'J]^�u��(���*͑'i��nEFeT�/V��a|wY�+�WA�g��G�vs3����vĄ,�mZ� �؏p���	/FlS���fؤ�L��N*��7�YgLD����]^�e"�J�G�3�?*�?ȍ��sx�$�!=C�7K����{)Cr����?(wx�SN&ϠR��	Mp+�"Ԩ� R�� ց��o�e$�/���pl#:yw�4�w�����iZ�����И�̌�B�DCt\�+=�$��K��(�mM�bs��#�$y�������.kԆF#�ʘ0-@�s��{�en��>� ���\P�=�W����j�&&�/0�(eO�5�o����+s5ԁ�e'�Ɲ�������L�>�۱��I�Urڂ������s�WZ_J��Q�~i���!��˖��1:���z{Y�����Io��1�S��#�!�P����̆[nc�4i[����T�`��ʰ��+�YB�U48�ցɔx�ʓE��t`J��J�X�H����� �k<z�/�NCw��n��"��,�cZF�Z@��Shߝ���hj�`P�|2?r�PԨ` �)���S��i��;��t�s;\��R��j�;�ҥ�)���.����zl <��"�:3Px�D��،�*��ɘ��-�����o�=�E����#��Z�&؈��Pn��r��R.�X�4\E����K��mu@%���3	�E^��mgq�RI���[�����M����ܼ�����/��]�L��휋�@˨*��jZ��5���O�㗅I8':�i�z�<��N0��!��+t��)���g���+��-%��F�6s�(��+��h��ʤ�Sٻl�`�'J}��K�v:�y�Zez�$�a(>4q,�"��XZdGRs��I*f����h�ϫ&�=���`�>��+��#�`�E�x�l�irU��y*��p|Y���y1c�!޾����f+�X�=m���C�r�,���Ls����{ I~��	�����8�a2� $��Cħ,��ڜ�
d
uTŷK_��1���`)����s��YB���"t8	�������6�;������>~GTBǦY=�L�{��=-����W!�"E2�E�V��~��IS����\0hs$eb��A��\,�E���L��.�z�8��.M��`��#�\�i.EV|�e��J���,&�YD����R��t�����Tuq�l�fi��M�Qm%T������>�U~�5��Z̬��t^�+�`����i���"��i"���p\��c�%���5vL�Jtp�	��e��%w�.1DFqR�M;l�(�sb͇(?�ӊ�6(�p�F5�w���rQw&�Χ�<��WVg�?�-�w���t�Fh奸��~92��(�gB{�w�1�A@�i>^�V��U��y��X����D��Og�0ES{����y�R}��g_�M��~��Y|�㾓7���<