��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]Ϭ�1��@V��gDa�~� ��jǈ�0I��#S�('�p|C�Q���S�jF�^���=#s�ZW,����;��fQ5[3D�!�s��R�����d�F�yKd�H�l��t4��x�^��G�WX��$	��B46�wn����Y�nLXr��Zr�Q������xvPҋ����U��c�G��7�7�
���*��rH�>'�5���B�-��:�p��i.f�;���%�߈w24	�ϲ�P"�䃠OT��#z� k�֪��N��;�.�D�L��p�l���1��Wp�- /�J���"�� h_	���$F6(a𬣭�՚75tet��mq�f�
�rhڈ6b�	�dMqi۶z!�do�����V�z�h�"��t�TD_�h�MʜP�f����;M�r��)B��b4g��E��A>B;af��U}���򨚐JK���VJP�w�b�N#iH�	��� �7��e�)��������O(��#�%`�8P&_~�_�6D��۱��bw<׽9{RQ�,esn�%'W�8f�l4�.P:���у3��v`h_?o\�G>	a� Y)'�%�iH>[:)?,o�ϲ,c
�ڽ%�����4D��+�E�(B�����V���o�"�r���I�i �������=���+����������SZ?�0ׁ�n��w��j.�züo4�����̳���#��MBD��};*S=A�q������q9���hIa�����qye"�8m���^��:�	�70W�����l����LLA9�E��������,%u]po]U=�K�8B&=��4�D�P��b���P
|e�s�2Չ�d�Zs�k^�OY��0�Ύ������v ���?k5e���}҃@Ĳ�Llc��ܜ�$=y�}�`u���A��(��	{z� W$���R<����Y��N�|�%#Z�ځ>&���o����䪥˧��q
��ʆ�-��G
��	HL�_v�g.=�@�R"�4��6e7 7�MQ�zGWn�����
�E�Y�;F�U�pc4ؔp�ɒ�>��B�$w�@y��/�����S�CTd�=�5��T����:��Y�����L�Mf��? ��m��9��7#U�:
�݌>�.	O���ϙS�L�h��[IX'a�LDx�ȹ�e��u�W[`IO�/��E
��m!���~�`��M����nΠ�&��)��X�r�a��,��	�8��GL"���Ի�T^]�"�1��,��_+��{�]�f�r6�l�wo�?Y��bw&8�>>krb�f�El���ն�r��Q����^ �_.�B�k�M)C!̈:s���p�g!��S�)���R	��</��}�}���}����ƒj@8Y�&p#Qh{��d���̴4GEY�5w�i�B�{$���_��y�/�81��8�����;7�mИ�|�3�4.~O!DÆ��#���O)7���<(Wnp���ͷib�a+�r�`�С2)�.���FRȆ	'��uQ�e0�}�v�#�~뛀�d	���a�ga�u�֡8zuk)�u����f�k� �~��0�J���ܐ�aGr���S�r��RT�ɂ>�l�Ơ�A�Tl��SO灖e :�ht��&B��fy���3���x�� YI(���	����No�O��1��B�D� ��I=�z��=׈]#���,��g��^b�t2��r�S'%Q#��C�M�VI5O@K�Z��ԯ�>�4�N��	�i�>�w���W��0�` 9�:���F+�(��U�vD��zTЃFHSi����g��Y�ե[P���؟�æ�	: Ͱ,闽Tp)L��s.���mJ��](no��kH+_�Ov=,���W���BS'<�Ü����~�t�)�+4A�Ʈ�.��1�c�/�˺�����3/���f��!�l\Z��e�{��%��K�߰yV($W�	�T���U�?���Ū��Q�bJ�*�.��><%�q��E���r�(�IK���ZM�����>�V��j���B�x�YV�l&��y�n7�WC�muO��π�J5��>l��v>9.w&�bt���?.xۍ*�cQÐ ��ՉSCw7]��ٴ��
k{_��B��HZ���rG��SH��B˼/u$t��D��չU����l�����Į+��!Ƅ�t����'G�{3Nv\��];���r�%ܽ���.n�Y���[�N{�X�a�0�d�9Ǿ�e$��%sw�9�"T;��l�V�����t���U�x'�6o�� �޶Xj0�����*6UoJ���M���:bqO]���?J�È�(�y��,�������H�)��ak(���<#A���7�Y���\�'(^����kq<A`CW?s���A�ɹyR���C�l� ���6�"�="1����y}�:-�
�=g(N�+ڡ��:|b11k;�#�I��#-n]�zVI�f�
\�4�6X�(c�/iȀ������;W�����4��2���A�4�C�X���b>~�Q�%�����>���zT)��{З���!��[��.q�m���6�����y�}1a4�x�a-W�`F:|��,J�/���h����I0�*u�!WlU����L=�z��i����yԌC�?����|��$&s��@ҏvO��B�,���I���,9a�v38���DР$j߿���OU
�$� 5�H�;|�\b���P��0"Cs�x����bL�0�������x	���$A���6�?wm��~	d�!���<�_��I��c�Bؐ����DPL��h� �r���'��Q\�L�@u�.2�j�vx-�#�=ٜ�ȡ�'\�C��9,�9���^��A��Ήj�}��@�8]%�OId�CVȆޭ�]3�n��כ��ܢ��d@�0�;����^��+͈� 	`�胙`�
en���lTM�����6D�	a=��,��"�'���7Q�F�X�_D� 3��D+߫��W+�������܀އ�
`��,�D�m�y�s�{�m+���g�'`)f�,Ӧ�'���6<	w@�85P�r0�, �/�In�f<骭[r1S�qd�VWD�i����B!c�|9W�$�M�ǶyC��C�h�Q�3)g�����]i����c������0���T-���c�v0�L�&�S��w�;�f��攰�'�\sM`Pxa��9O��C�)�<�Xze%���ؤ��W��U�{ö�#�6����H�rt%|U��;�}{�y�_�+�1�~H~��;<6�(-���)c�x?BP��f��%����x�oLn%���T?;&��0�ⷖ�P+�}6T�Ac/p.��)B��p=O_�޷
���+�'/�7��6�� B�b8s^L�{�2BH�gh���R�
��"�!mI���� ��m���>;2V9C��N�
Ð8 ���뜔%�#AF(��ט�K{t&�:ׁ�vB�:(G �؞w�����kK��&7��!%Ř�/-]o����V���h��`���_�olFitUc���%"�MVДI�J�5/����/�s���ܻ�)��
+�2�)���G�F����O����G�%���2�s��������DnPu��Ҵ�~n�
-٠��Iq �ژ��B�I�RyK�h�Kט��o�@>��DB	f�BҜص\o�l^9߀��+�A�Ϣ�h��C#���Fx Q5������X���n*j���D ��0yv�"w*��� j�%4-�t�SD���w�\���vT�;���U�9��vV�`���5(f����"6��8�q����Dl�S�%D2�Q~2�‡�/B�2�z��DJ�.s���hg|*\��M|�"M`u������F����e-ɍ����	<5�8��o���T
K)g�V�ln�\?v>^|
�� R�`�K^��g �z{����8J5�%�;ᱽzwJ~�eZ��J��"�*�/:��.)'��c.�� ׾�����F�wd9�+�	�{l�z4�xHhÍi��9v�,��kG@�P�0�;��Ǳ���j��c>�4�v7�as�#��[�|��O��f�e��uj~;��x�̨�J�M/�B4��ڟ��>�	�S�?�^��27�La���L�$�7ߩ<@�zx�砬�Cԡ(��{.�/��'�`H+�=6 �%�O~"L^Q����fm;�+�TOH�3�X&�K�ӛ}��3���.iB�������$�y��V��gD�˕g}�n�N�.���Ab�<���4��$���п��ٚ0$�t������#5��K��^hT�um���"�f�����ZE���(�����
϶��R����sҀ�Wȿ�n�',#���F���5���T8s�H�����s���c�=$KHn�U�t��@$�m�Ï�"Qò��v���}nT�2/���"�39q@�R���s��l	ȝ�����KC8�<q���݅(���Q����HC�[}��dr��~�"
�lI��"�Q��v8E7�/�y3�o�Iqϯ�:�U�e��r��{W̳w+���
�JЪ����T�{�[Z6h��`���1�����Dm=��P�h*.�)Mla���5�T���n�p�w��)�S�1z{ �<L����aߖJR@���\_#Y�P,;J"c"�Yo6.怨7q;?:��=#h5��8�$ѱN���Y��.�3���������~9o�̃��77x`�q��v�F������2�ʦ�[��᭗�u�0&.�@ĉ��Y�7n���nw+-�T#i��I�0TN9���ۆ��-̾e!&� ˂�s�5=!�{[]A�4,谶Z��O���{t8;��i��ʹ�SҶ��(�k4
Rm4)��墕�}gƏ<5}�x����"�ξ�;Uohc �$Ty��h&ox~�	=���M���pX�#&WIǙ��f ؼ�I;����BA�Q��զ�JN^N�
�S毼�)h��NV�Au���=���0QG��ѻ��t����Ẵp�8S��7�Y��KT��9��ѪZ�@�"�i>��`��l˜�?m�:��Si��������	x�%���A6#{m��Z��]���k����왂^ǝc��OSV&a,�,�{���$,@�(�6}7W�������^�tk<���J��G����}�­��2�X5S��y�~���\�
��m1��O�Z�.�<љ�f�����xF��u���eK�L��r[e��-�S|'J��Վ��+7t�0@R��ln�̍�YŮ�6N�enG��u��l@��&��-����� rM祪��Z*�_�;����z�H G��A��7J/��7� ���ɍ^�����#!yŞ��7�>��/ܚ]�훏��=2VK�n��1(@��J�b�A���n�\������g"�D.��?��d;�Y���p��Q�q�6����;��5��`B���e��}�'go�V�&��O����*d:�|N���6��y뚨LY�y��x�\��J�����/)8I:�2j�O��J��L7�q%=&�0G�	�,:�&\�~ǖ�_��R]ڴ\����E�u�n~���ׁ�2r�%��-G:��Le���t�p��$3�>gh2P��>�bB/�x_��_��:a��9p]N7�ҡ)� S��L��a��dZD�I%���Y���'t ❩ ��Oe{�7��S:��^�8��xV��� ��L��d�%�1��}(��|M��Bz� �����(˗62���vΘVI�^��hm���-/�3tG�nZ	�MN���s�,ŕ����:�S?�K�P�$3f
j�5-�k���E_|j�����j�[��*UD��~�w�Xλ�8
��n�c]!��v��T�SPW��=��]]��$� *�q��S��`�L�J#M<�S)�n�M�*�@�x�۩��x��4Ko��ɨj���� ������%�C���������P���e@�	J��@7Q�#��b�����H�n��G�F�Gu\�iėr����
O�I�ш����֭p��A�G��3�B��lo���qU"�K���r"t�����Z�~,�T�V>}t��k/���x�8ȡ�Hb�|q�*�:ȕ�?m=�*��{Nw�a���ٌ�m	�;X��yr)`p	�+��/7�(ǽJ`�%��="��ɱ�^��@���?�ͫJ\�K���"3�� �������M����s?^ͤ�Հ��1�H�0ԅ��]��S�uT��K6�����s$Mo<-�gDF�SỮ�u�U�BD���їM#�g/��fnp� qޒ�\F�V�z�x#Bٱ�Y#�����@z��-���0�(�K�ZS%���� ���V%A�=x���H��W��߮-�="cJ�x�׋$d���bђ�@����6����`b�ty��ϱ�Ꮄ�����T�k�i݀��D7�a��Њ� O�i@��t�;���;Ye��RF[N�j��$�]neo�3����ξ����x%Pe�D"��g	�f'��/R˶�R�8�̈́C�Ԙk��Sd0|�`a���z�!��,1����p�Շ ����8t�(������$#a������@��E��a�Wܢ��7��զ?	p$�
�&b��D���ED��F��P,����j!n�X�|���������4 ����3��+�u��!��.@����N�X� �Q摃i�nj��L���2����e�~��YMp��!W���Z����q���g�^=��U�!��e���q��[m��<h�n=͟uO'��,��G�|Բ�s�F���?H�YO���Rm���b�~Ns^=vtJ��
�R16ϧE�5NO˸|�_���;���bc|5{����Ch��@bf��p>/�ۉ�o��Q��r�mU�jn���Nb �_�o:-
��ܠf\B��%���ͩnwm+���(����^�oT4^BDF=�ȹ�':	W�ҁq{|�[ehò;ם�_\�&�K��=�&�=B%�*˪n_eo�bn�N�˪��jB�m9��arR�<K(�e��~��3]�d"W��GS=\�l/��S��~'%.%y�w��m�%����n��o�$@��HF�3`r��#�Ո� ��$�x���>��h_BFB�M��1-�W?@+��Z��\����7ͅD����;��~BZ��Nu�v^5�[ǁ�b�����b�����������KU|N�����5�
�٥�r�\�d(c����V��^!��~��9��5���c��O���o��`@�Z��x�?�؉��:R���=�+�I��3��wD��l����jNI|���R6A�<b���	�� qW�vȚ�qL���ۗ�KH��p
���B��X�A��L�K�q�#Q%os�p���$��0��1���`�o�A�Ǣ��h)��cb+�|�]������@�����Ev7�y�q�`,���o=�z�AV�����l�� �^M V��u�W���ws�ֆûy��I���*�vr�H��$+��U�������u�%h��^��w����(:�'/q�� �C�+���J��`9�U�`A�o�O��7	��*F����<L���@GC��!o�<�3+�N�BO#�+�Ë�R�r�-��[�:�y��I,0�A"x(�t%5Z��-���T�t�ƾ��Dj��