��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6�s��4��q2��P����s�j�Ӑ�u��b��m͹ 4�yR�tC���7�w��g�ū�O����ٟؒ&�
��-���WP�Q�Q-Xy����q���/����&��4�hH�� ��[8��<�W������"�"CBF����fxw�{琯&=�(���#�LͿB4��o�`p�!�ݳ��Q+�+�xY��uqeol� �{�K��?�,���.K1��͹����S�?�r����$��(�i����VZ�N��rSΐ�o���wLH�7�a[J���&=y�>)�^�0���/�wO�W��T��G��S��{��X�)q �r���ɲ� 	*�|ԴR���GA�I��]�l`��M�!������D_�J���F��/q�(�j�(��P��{��0���.|����>%�( Pk��M�����*�_��.l%��˩ߒ�fˍ��b�$X���5
�2`��a�V���g�Ik�D.��'ōv��\`� T(�b�@���Uv��$���BTM�k��1�����毪���a��ln=N�)�̟�g���{�ak�^����ε����2����L��HT�䢝F�Y+�	�7%�J6$K�z,mZ3�H��et�e	w����vd�����a��r�A$���0 ��=��2�bZ�Wa����F�2����.�+�ƇOO��YF�`d=0>9�lAb���'.w�.��
p����=��/�Q���MK�|�D�^	��8ݠFRXg�o��YB����v�n6GsB29\70T�&\c���<������yh�S��믴v��F��38R����Vņ0=`tW8�LON��a�������yZX�r]��I]��ϙ�_Qр�z���JwͲb�ԥgzh����8y�N��{�G?�ז#��hл�Їz�"�"�6ؼ����[�Q�^�1A7�F?M������V��8��J˹�w{�uG �Nҷ���/�Q8	�?�%�\��AeG�Ic�Ѥo:�33���vT{o���h���+����%�f�I�++CI�З�}�m݌�=���8���I� .Xu�V�4�|�0)c��Ę�ل!�צ{Z�ײ��iN^uh�!�n�RI0�$锆�|^@�GA���R���'󀬘���E�������b �Q�Hy���@��|���J����c��:*cFRLjwPN�sܒ�P�6����3�`\�o�N����yܓ1��1��d�/~涸Ƌe�&�f�Ep�����t�3�X��>G,�E-<{ZD����+��zq�uQځ�js�{"����Tb����vT��X���|�H�~�&|�2��q7EG��kf�ݞ.��s�	?��3:VvE����L��6Y���T�`qp5�Pl����|Ps�d	h^
/���h ���a8�F�#`ƅ4�؛]WZ��z]_�Nk���I�|s�2���ש�_�������G~�-����*si|6ނ�%U�z��J}k�� 9,�rNj�a�H-�6�h���M	�Jf�����*�*�3�d>��Q�z���8#%bwbA�c�JsL�%��Q��.��4�
<��C�V|��'��vJ�WD�Fߧ�
М�"�����ذ^��:i=	rc��z�s�-^w3W5U�V���7��4dYv��X��b�u��\P]f�e��D��2�}X��(�.����SZo��S]�	y���O1�nK�i	30�i�w�C+����}Vg���o'��{Ҿ<xR���es���g�ߧB�R����Z�# �A��h,� �u�"�,Q�W��)~�n�&�dk7;L�3g?6�65@QT��7�u���#���� 5�>�#�9xf�����%�Čb|Ry���3�i��"}:+����><�Qp�W%�-�*����4�� ���}TN<7F+�6��<�1��@�f<|T�{A!�N�����]li1�8p�Nvo�	��Á9o����?{���[&��Z��J�yǨ��lX��8>5�{�7T���L<�%�$�&��/���t*�^���mg�����<644����pŻ�M��5�/7@O��.�{�#��u�YjRR����S����Q~(\��aJ>�����y>>�A�oO�/����u�pe+�z���Z���U�(��?�� d�n�=�GE�d^��:e̫��3޹���7�zt`?���?A�f�|}��B�lB8�":��+3�Hk�kL%���o5f�́���2��<��04�����7Q�N�	豴vH��`_Xp[��i⹧�Àxf���u�9Zn�����ņat�SA꛱�50����\�Jw�r�΋b����8f�?�n`U�^�iVcSݜW�P3�][��Į\�G���4�a����ڴﾻφ~+����u6��+�v�9�3|�Ux��`��'�\�qi�@�E�	�и$E�d����$5s�`	��6|��,6������"����ag�@��ey���U�D������U��P@�B�ԓ�GP��VJBFge���m+\����WÂu�{��l����"sӢ0�]MWZ��۳Ou��sJF��QF�eƞ3�#��qd*^@6�Q����,��Z�.�,~�?ile�١>�E-���Q�O�د�z��S���-;.y�|/�D����$���O}�6���<)m��B��ͤ���Z�z�a^l��{5��]av���Wrݻ�&m���[D�����Xo�2�>._� �N-u�QH˝z��Г�y��l�����7'���O��\fCN��~}�#_7�D6���c��7��Tտ�N��s�o8W1{�O��#?/\�c^���DR63�����hF{̨֬l� b8-=��|P@rhX�BFstm�L�Q�7�t��y��˄V��w��D��1�[�T|�W���$�͑�
��e����c��^wr��,=��{�ez�^�>�-y�7��8=A��"}@�_�ME5~]n�5�Q'�)��E�{�#&�����<���)F�n]T���k�b&����3��Φs=q@����GC���M���l��t)'���f�M�_yfHk��(�> ���_�!�y�[�}�9�%t�6��k4m@���qߪ�ə�4W�.ew�.Z�i�Nl+�!��x�u����p����'H�0U��i�S�Y ��̛�$ye<����Dj���MF[S"΂�=�6�&τx%8H���h�
���T���7��l���y�ff�$O�zs��m>��Π.%1;�c�n��\��=6��~&qI�)
��/�x�t'B���w}Q������xcr:x�]z#TlV���Uy�F�����i��i��P��o}o3�����9����U��>:��A�o�z��Ꞃ����F�C���r�9���M߫|��ظ�G<�$��4���D�~��&��4sC:h�!�_�|�]Rl�ƭ��D���b�C��R�nn� .y��qi�Q������>6�7�=|�J����
��Mn�6�%�1*��z�*�C �C�N~U�o�v���u�q<�n��a�/C���c<������ʸ
�.��~���������cjE��jtt�����@<7M�w��T�M���bo��@g�<�+��[�8��h�mԙ�<�_�0%�"@�C�H���}����GV�����\�n�U��"��q;9�)��F�?��Ev��w�-&n�cUM�@m�Ox B૧��h�;�d��]�h'��V�#�PŒⳙ%K�\��/�u�SH 6�y`U������"�{��o�P��X)��V��V��]謯_�V�i���:e�����h����>a�*o���O��z:��Ж��^��J���˪�l����V��B:.�;�1�-`��)�:���g{uv�0���۰��H��H�.�w���!�yw�{�����x肷�|�����+����2���5EV��r���J����R�ͺ�"�`�
�� ��ϓ
m׆�bF�>���c;�n�0�^P�^����~|��V����e�-�=䁏mk�n~����� =hY�c�="�%j�i��`�4��ߨ��m�28&y��t��L��5M�Ƨ{1)(J��eu�q�� 	Rʏd;����~Y:��;���&D��k��\��
�|���W��opDׯ?���-������n&�C�"Ǵ�Y�~ҹ�X���r.�j;H���ʼ�vz��A�ݤ��5���ʠ[E�aO�;�́6�����O��Ԇ���Cf��9jW���(��ж�vH�"D�����l���0MT�"�`�U�2� ׎1�?��û��[���D!�P����h*�r9�?[�}Wk�C���Kˑ�]0G}i^�0&)Em�I���4��8���ـU�����l�o�9ő0�Mq<�'�N�~�%�LC&�;}Ú�l7��,�rq��8&u-hp#�g~�p�k^o���"
��>de���/q�ρs�G��q4��U�BL�$�,ܰ#���;������rP�KI����!��wgc�x���J�<v�4D.�yrQ�p���i�9T�����Ɲ���%������_���6�+&X��=UlCz^��2��\��D�|&oe9ۃG���J��wUB#�.e%��*P���A6܈>8�
���ޱ *�3��أd�-f�7��uP<j�}�?M:��\��p���6�T�I��%����Z�r���C�䲆ap!f�r��5ѡ��a�b;`J��Aڎ���-��ԎSY�/������7W��6`�~��o���G��E�����Iid�b@����Ɨ-����w�̶�����'H�V�w����|!�������n��7d	�,�̟It<zծ5F�HJL�Me�}�֛����T!
3i���ꭖ���ڻ`��2�+�V��B�t��9��F��7�?�=Eqo6��=~M���0�˸{f<!�>��q`%n+E�+�U٭�Z��Tj'��B�*�w�͠��S5����3��6P��>��|��Ѭu�M��>�{���ҿy�����F�����a�w+�
Kp��뚸p��<�����
���Y;7	d�#-zR�jpN�௧u�%�Ԋ��X	%/��*�l�gv�C��s�oZU[9�
w����V⚦�HN�l��F������������:��l����Ul�4�iQ7��)vO�~�5�*7 �ym�ރ2a�$��X!���[D~B�h�F���n�R������J^ee��ҍQ�W�yj�6$�~��.8=t� "u�i�h�;څ?��� ȶx��]�<���:oV%vf<h;���GWf����Cd��h�4x������E�o�ՙc�f��� N��F���u�@��\}e(*+�|>�n�X�S�����ȏ�ǆKV�nP��Hj$�"�W�E�g#�M_�
q�����DBF�L|q�DdH�	�ɝ�~�`
c V�/��_r�`րȩ
�,�C q�5�u�*R��F���#�!��웒�Y�[M�G�D�q�f��@�s����n4i�1��Bf	��z@7����D�2��$wb*Pl�ڢ)U�+#�K˿[U�g�{��Q^����>���w��k�mιp彐���r���zb�'p&ܗ٩fGx�����D�H�/�{b
��?s��I�ֳ9�[�1VrY��D�m�M�+F�Ur��w�C����\譍3Iz;���q�y3�KdD��8�0�#�vے/�u���7c�=
��N�Z��w~��1����S�n�J��ot�Z8��oB��}���6H����� �s�]�b�1��gd׃D6h���,����@��tnQ�Y+���Ir��G�e��B\m���f�ː�Gc蠻�����؋ �7��+ڋEv�#p܉��I2��}��_/lI�d[�-�W���n'\����Xfb�FP2)��Ta	{Lh� ��U6���`?�7Tv?h@�/?侂�&�82~�>�Fl׏{��^-o�-��͜���Yk��10�^V��<�&���h[���%�>Sײ�"GSI�k;9	v�٪c�V/�O`�Vբ�F�)`U�V'��~�=��E� �b���gOQI-�Ma���5�iN�����R����8jY�'>f��;���mĉ囷�A�'T�8�N3�P����'Y�b���W�ݵ�qs��a��β�i��r��R�{^���.D��n�V�C��䬝Y�r��g��/�H�#
�d�q6�>��11Tz&�4l%�j�u���u�z}��HФ�t_�4�K�"PT��"���<�ͳ�����uz��H�Gp�,�!q�h�nP�N<	x��!ĭ^o.�@�)D��OI��>S���ܟ���z���9'��-��Z=� 4tF�c��"��G��~(��%��E'],��CI!�>[�w8?�"�"���]M洎QxmU����6k0f��y���uVܢ ���
��uMwQ�|� �Fz���m�Uc��i_��ĕp�+�(cޚ�b�1�_��_�qd����0�:�]�BD��� ������p��	{*-d��5�oG ~D���U�d�w�wĥ�b�@k�5#�{Z|zy�e�q�:pSv8�D|�JW�z�H]{���tO�9��Wa���G� ]@�^�>?��Y�g���Nof6��	�: �����vOW�>����>:C��&�k�PdP���Fb8j)}q߭ʁ������)H��4��_ن����J��:�9�.Z�5ގ!,��5��aj��{��&=I��1Ҡ��AS�7Nb��y������7��!��n뾳rJ! �^�k��۪������֨:7�v�����>s�j�SA|� �m�b3�b�w�����lZ�����_�5P�t��h����H
B��� �z ��o~
�)7z�
&�}ݢ$�����a_yf�M��8c\�'Κ��l�M$ͫ��P)	�L�h��롟��t���;w����Z�?��D��p��s������+�hhx{v&շ,#��9Ԯ���S��
;��{�Hi����@�wM�ej�����+�"�P����b2LO�-h��K�O��/i4jL�[�%$�X*�`��9���[Y�}KT
��-Sz�Q ��B�\B^Q�OTV��h',���m�rT��a��-{ ��0��b���Ͱ'K��.��>)�,�Q�W҇�Jz��ƥ����68kI�N	�:�鹛���$�H{x�����ϲ]Q(���T��`�nD����ec*{F��U��\� �K<*��NJ��'؏m�iz�;o���Oj?����\���`$ʗ�|��=�_��Bɾ������׃���Q�;v���"@[E��(�T��w㜯�>�zME�$u�/��dA⥹tҜ݌���N���_��'�b�T:^��d��p=�f�T��/���<��sq\]a46�>��d�?�����|L�L��z��3�{���u,���@�#%0�Y-���őZ�9ͤ��2\	�(ʖ�U�y�����3B���[K��>�aM�п]��e��fz��Y��5�X=;�ZG�1�����/�
^4��������\vX�&�������`���_��� c�ܐ��CL�R���1]��*�*!Z��J޷���jy����u�6��o�s��l�S����-�zl��?1_e�A�0�651r���e̗$�����-)�k<�1hӁә�R���F3+�8�ⶈ|�w��h��rK�46=�ȫ`�R������t�M��bj�Y������;�oVxr��+WP�A�9WV��D�$�h��oxS��Il+�A�����x���˗�=!���В�U��f,#�o	�
�~�B���9�yA�$�n�Z�3�)߽)�X�T��4y��>h�w[�����}$�Oa$ѻaC����+��E�q2��d�杬+0ɲq��Ppk�l�~cA��b�T��=)�9:kQ([m���C���ì 3�Q�����H���q*YQz�)$��B������y��Z+̃�(b���^��I9ptdd�VJp�#o?���F��6�5!�a��@ ��^��u\I�#O�B�{�U4������5LgG/���x����K�0���@�gK�9
)U\ګaڳ8�	^��Q&��Ț+b� @�2;^�ɫ@��S�"OmK]����tP�B^Gn��~T�d
����U�M��>y͵����ۓ�1N���x\���+ ����r`$D�`�c���,��&"R�K^���uX���"��<�(U/��B�BV�,�!�O�y^'��eX-l�G�x��zVª�ͭ�+�k�r�A�U�� ue��x]piz²K�A� Ʈ��zg� ���f��UTw(k�7��IN��A����C�)�n���!P�6j����o~��Ǝ����aKp������G|���>O6�K�}e���.*Ҏ,�����#KH���|����ϔ��Q��݃��}-�]�71r�#��y���~����l���o��H%81n0~��#	��C��D��B��_����nmd7�,��Z��a�Z*��)I�𳘞���7W^o�+�\���v�Vë��|��l�)E���ށF�W��a�dZ�K���8jE���q&�H���MZr�#���C��[�y����J�N���b��/tшe�"E1
�ր�FҞ���m�BK$���y�����b����5��vҗ�BMGhsث�Y(���X1���0�.���D�n{A���0�W�ͻ��ɧq�Ls�J���>�3���� ca/��]�l�/~����V�U19$~Q�o�vwd
:�dKU�2�[�v�L
��~��@5L�.RxV�ɻ�xOPY�}��#�cjs��})�W���W�1�)R ��/�>���2o��Ho�3�����hr��^��ih(̟*ۡ��!��V@���z/��=kDN����o��O�Y��5I�Hv�\`Ű-��iTk:���� ��NGi�5q}�����qC�:D���
n�R�4���M���4��������Z"��ak���Rd�9V[��=c��weČŮ����<y�c�jH���vC' Fi�z��2W�@���D��c�-,�?�-J� Ж܇)��穸�'r���J��9�j����=�^!�YE����	ZS�~��;B�3�M��Fը&L(���]"�9P"\p��{"�V�5��N���)�B#��4��u�%DY{�F�oC�g�V}�kG�Г�ӌ�mvE��d��a_�+��t����й��Nh�7�Z��	wֹ�rS�pq|���t�8=6����g�o�ߏ�|�~O�׆�i)������RG��&��D�#M�8�ɀ��ޱ���wAKm?y	F���g`4K�=���8%YG��1���&+�5��3�S�/[*���9P���=>9P���|��o�3��²��sD���#�
ӝU��@բ���G���n#����U�����HAB>\_8m��	4Teh���k�3����M+�Q3������ ���!no�Q�]AFo��¦'�|d�fsY���a��ٜ���z�ܶ��8�ئ�K��:���������jҼ��a]���.������S�r���n�j��@�L�jL�M;�72�پ4�7)|�+��'� ��x���>VTab3[Th�hbG��ն�����p�q^oL�=�\��/���5��W�J���3[�y?�f��J�Ϝ��z>|�\�#e=8;c�ZN<���I����`��i���"f �#�C�j5!���f&��"��I���&�^������Ԫ���g�Lϧ}*�e�-�`PQ�֜��#�<5���d�y(�/L�8���
Z���I�":�Ru��R�k�ֶ��O|j?48����E?����c: !pk��GO��u|Z�����j����޻���R���0�[V�u� �J%�x0b2��f[jplF������������������L�AR���
V&|-��w��jҽ�O<�N��_KCA��F����;!�'���#��c������ʁ�{�]���K�:�1��㔄��꟒HOmD|���w-o�}���52��!�ȱKW�_�!�I�y0"��!�!�W�����$RW�͒z6����q4RG[�@ɖ��08Ģ}�b=��]�?�=A�rÍ�V���e�eرW�KKz�:G�����̂�N������/�kBt��c��1"�F��K'������1	�l�1��6*�]��bk�ž�Hh>9�%vI����Q��D�V��k�\����ѭ\����jg�����Vo
�#�}l�`s�Q6O�"�𴘉m8F�·^�V�!,�\&y��.ʦ��f�&h���/���u?3�W#\0�����7���5E��yf=�K)_{^۶�����I �+��D�%�d/�AS_(��(x���<:x웧B�+T��	=�!S8����!�ܙ/ߩҕqY�h�${$#9���nG��y��o�2~�ت��${��+-lY+A�Jӳ.1Y���d�j��M�	@���ܽ�1
���^E;�HM�a�a�h�%�*����&�D���ϫ U��M�]��#���w�ȴ7P�~��ű3�:�T��"��fRcR���������ťu����Դ��ʳ�Wdv�g��,����H�]�rI��FO3X���(�8��|�BQgc��GN[�%�<nQ�]�|!"�j>����e㤵��X�oqQ}�pZ8E���W���5���Lh��#.�{��c� ZS����i��h��'��{����.?����ac�E���:EK�A�j�0o���z	�V�c���C��'U����F�Go�զ?�`���6��V>z�EF�B�>������s8mF��5����%���9�*�|\	���T����f��h�7?dY�>����rW�u	��s��`��z��r ����5� ��$��g���רC�x�j1O��P{6vfʱ���/�%��-�p�z���u[�[6N��������_nG�(�7����?,O��ŷ��n�D\��#�g&�0F�L�̻O^��O�+��z���y;�o� @��%l�9��,�� �s,N�J65�^���!tx_U��Y�KӸi��k�v^fv���:�):��
��*ĕ,��7\O(Ob}�-~���%O��5��y��
��!&�|�|�ˉ��?^�gյ}0Sl���w`��zJKS8/1[;�%�Mȯ���o�6�9�u�\�^�͝	�m�#��z�G�7�X�A�'�BF�V�3W��[���E0񨷶�jʀj�.�jr߶Gѽ�X� ~Zm���2������=Ը��5����!�MZoAS��lê~?����<@�Lꌭ�
ȗ����n�$JO&+^��z��Uy "&E�<51ү+�W}F�GF��"�r�Y���v�䲬>k'�d�-ELZ�l�=`�_W�w��`��c3t	��[xdK���zoDxѻ!��*��[�|�_�^ː��5��d��DbJt�J�*Bv���Y
~���dwn$Pu�'�}a1�x����7I��yۡ�ti,�zT���k>�Hw�O�u4.׻2M��
;P�>ZC�5�\H$�a�Z�z���V���㐧�oA&0����2�s��\�`8l~��U]<�.��{!��+\ur����ߠ{���I}�>����(�u�k��u�4RѤA�$U/`q��yV�@���=
��O��LO~P�{)s��-���ϴ#g�E	�
�L!��J@��"ù�tl�z^�����C������Sܞ�(�b�v"xta���pZ�}-�Ј��!JZ'�vҿ`�9�Ij��ٜ���������˵B�O��_e����njQǯ����2�(,������¤Ԫ�}�ĽF�A+l���|3���:�8q�Yhbk���_����b{L�/y�@�&�dj��^�']ie�"�b�KC0 �dcF��$#���V��� �1�fU�� ��Q�X��s0z$�{�)WbK6�i��Ȅj��v�ٟ�
���D����,o�q�/WϖZ�i\��a��/R����r�����=l���:��
�e�^5yn [�|���*κ�;����&z��r�i9I�\����͓��#��#� Ċ�!�4S�e���$�Z�D��OX�ܔ&������r��.�'S�m64?���3"��/ \���)�h�"�DxRf�_�N�bJ{d� �^tݩI��W�yH������ �bi"Jb��ن�xj:����s��o
�^�ŕk��ʌ@"����ߎ�+S���L�	��E��"�k�jW¦%d$���	����Yڳ�PJ+�ՓL�xV�`�v�lX��K9��7���yX����u�s8��S�f�;t�R>��߳�ORR��@Y%��곉��՜�pZX���<�)<-
�����u����3�p���zp�E�j��%Í�����E�4���gJ�=K�BQ�?zz�\�g����/�~�EC:��@�K��5\��T�`ҍd��C䧂�~I-A�]	�X����e/��t+:�s�ɋ���W�}��!]Yg�EfA����N��{yZ��U����S�k�m\.�K�����=�O\9}5����R���	L?�$<�5,��5K'P��̇�I&t��Q�[#�yw�U���Jw�T���%Ǯ����YJ�]�k��lI6�@�N�i����w��z	�(��L1i��q���*����'��}�x�+�x�I�1O�vr2v����G��J�xt��q�mYꪟ�5q-s���a#�Z�z?�KY�;�O��	� ��9:q�؄�Jl'��~�x������H����z@|�{�,#�1�C\���䣱K��z�Y����@���}��i��t�4aA<���̆���&?h��Q�ޓ�A�u^	�˽jc
w�K�DmMmo�o�<��'QX�%���J�0d���m�����B&c�\Ia��xW+�����'��'sYR�J���3�bn��g���K�ʝ��BB��`V�}D*��n����*�37��p�A ��Y����������K]Zx-�Gy�I�<�yi��FK�J���F��}iWcBV���^�u�rX�БlY����{�6��8��=ywW�2�z���^�J;�����CD�r,y2F(�i{Ӣ ��ݽ����Wv�D~�F����r	���1{VJ뼮��J�ָ�fw��= tT������$��z�5���p?e�[�3�|M�_�����]����'���H�N3&\F��"�'Ū(4p�f��3�jl�<v<��.i�@Ţ;̍ܘmi����<:�6'�E�j]Ӭ|w)�d����_=��C ��^��9���#,���Z2��u��=3-ʁ.}�d�����%�����Z�
�H�O��Q �@�&�]��U�dE?�TU1�w�@W�Μ#Q��*�4-���Glg�`5U��A7У�)ع<����=F����XIѳզ)�%+�� �����w�v1�x��髹;7`'���E��tE����&4�e��n�ET���=>�qu��#�TE�A����O���28�����'�[��̥�6����#+��J�hZF��px~��>O�R�ې����>��
��KP�z��u�UN�(�rb#�kUG��x�`W���B��E�+�`A�@6�U��b�?��Y��lr�k��"��CR��䄱i�+�
w�-�7iN=�Kk͂4᮶^GS!�',<L�MKȨ�Sv��'�\���h����K
Y{��(�N�9�VhcG���h�$|�A���}���r����P�b3:V��T�4ı��EY�m�S9��C����
�)�CD��?�D��7���ߠ>U�}��_U�J76�n=m�3��w�Tl�i����s��s'�����8eI].�0��ʺ[ez���ąc$�y���Q[�Ze�}�d�_�KC�"��p
����;���EM��R���++^���T�����x�b��$�;��w��78���^�-�o8�2�=i���D�7{W�'G�5ǟH����wzQ�:���]�˳�^3�?�\`���ѻ#��ܘ^�]��/���ڵ����	p���A���y�)�E�`�S���-��4��Os�K�N�ˤ֜�
�y�20�[KX�K]N_I��ղ�mYR���ؼ��|g�RѾ�<j5~<��������������58��2�{��E���˔�"\�.��re�n�u����4�K��L�`^�h��fc��si+�9�`��sc�Q�ħ��ba_}�:��fJ��%F���9|@��Z�ƀ��/vch�8Sʸx�&��cTn�Q}Pg@D5��rs7�SFdW�HrG(i�̸/kf��±��˔�l{��􄘌"&N���pGᚁ
h��(� ��}��"d�P�%���2����п"�a�`!k��`�+ �<���<[�����*u���C��uUl`m�]��݌� ��*�>'TFe4�&�"U|+нVR�P��6�%Z|!�N�F�{��zc&6�!�5{i������뛾~��3�$M���I	{? % �e=���dr����Z���T��|7���f�;|j���D
��y�@,�t�׃��B�!���_�)KT��sH=��E������T�@&8o��hş�0�<]H��"��un�&9U.r��(�V�����ְCo87��28m��܅��a_�=����4@��q�͍nfC��� ������c���5ԃ[�����G�r���c��wH$�������!���g��^w�ۺ��i[�����k�2�#jK�o0 h�T����0��x-��C���TU�l��+����D!,x��h�v�� w,�=>k�^���|پ��L��%e���~�]U�~YkI!>��p�a�^�{�S�u�D��DpST���]#��$U�88����N��r�����9�t0�q`�@���8UW'y�X��q�P4�Q7���&v
��:Q��%xN�aP{�gs�����Æh�6l����@���EvX?;=n�c)���0Q�%'�(݊��Gy�q�6`���e��Ym��k�U��Cj���aE(�T����}�=D�D�cG��!!��7-[o�u f�=BF[�6�q?4p��	E?.�b�	i�J *Z�]�~<��?�kI�ុ�`�NlI��P�D�L =c� �C��`�z>�Z�RDK�hD��&��.|!�Tw�
�^W��2���4D8F���zC;Rv=�2���������BhJ����ŴDTŊ�� �Gp�a���ud�r*�CKk�j�j���c��p'F���ܓ�䖆�JP�4>P�e9I���o�Y��շw!/�h�/$�׹)�-�W"�-�&��=�X7$j��[�98�<o�VuY�Sd�Ba[x�*\:�U��_6U{{E[�i�Z1CJP	L^���"Y]Kz\D�!���9��i��֒�h��du���\���T/?�.gg��k��X~AN�K�-�V<nX�-1L7#9iqY'���=�d�����²�v,�7+�r�7�O��
v_��#��5�kq� ��x3P�$J�� Xv�����*�cp�2����ߏ�+uF�sd}��p迹)Rkn��� jnJ�v)�-Zu{I�����LD��W��\
wp�ү/��'���ş��N軅|Vm^&q{̅�q ������i`��dK������A��粿�IjN�:�4����JӔ�hE���e/#I�E�ɀ�у5��o|4��홈��KCͮyi� &�������fg��J���z��t����T��8�,Bj��1��������
���������_\K�ե�;�Tu�
*a�!��EK���M}��tQ��1���ƵQ�+�Kg؋f��-�GR�����2 �����%�c	�`�W��"t�>�oogO�;��p),^s�Tv��o����tbd��y���us�n�i$�R�Ox�<3Nyr��?S�>�	FJ���gh��2�NOV6�%Y��oͥ�
oΚwR�#6���q����B��X�:i
�VD��*��I��"�����(�+l��02��?������)�dm"#X��z�p!{�ǹ�����#�~bfz�rO�.��UҥD�P����a@�T���T޻kR���'��d`gG!��g����0�:��UVJ
{�a0(��.���3%��8�9Xz�n���r k�,g��9�ᗃ*�q�i����q��qWj>:�>���v�(є��F�K(�*�*����`��Ŝ��*۾�aG���탞}�����?�h�� �c�͹�tʛ�[r�x�#T��>����� �>�O�Y9H�����h<n\��<��U�1���c<`4���w��D�Y�U��Vt!Ꞩ����Ӵ��&��+��1�/�r�J�x�[����7�S
��i�.Q��0��m��4���-�	��^P'V7S8��<���Uٯ��P��:�<e[��L���+�<y���&�Cݮՙ�t+!��'���S��E�c�W��DS@$��(W�Ϋ�8�XsP;���Md�1�.�#BT�N��P�B�ک���˻��R�]4R	}�1^� ���_����Ɯ�����-��eX+(&�&R���~�����e;<��uB53�RnZ���'��Y�(�ɇٖ���XKn�L�T����Y��x�(�|�WN ��@'y�F<����3\�\+ZОeXV��"���O���I�ʨ�}4i�e|����M �G[X~��⮰����O�O��b�Y�md�������ܖM͊ױm��,m8},/�
L���5���Q�Z4��Q�W�Қ�ha�p���Ŋ3�f��8���U�iP�^��b��B�A�ZA�4z.��zy�3,!mֺ�6a��k���K����ȝ�5ۓ-Gt�>7ᔤk'�2��pO�I~���o��,��(m�&�B1���m��'�(��H>��6�1v����UVS��hռ	=�X(��>��9��^E��gL�^�I���BS�Gb���¹[���U�v���P�-�r���Yй��r�~.un������+� �QH�Q�w�A2�.��P,)��RJ�$(�,6�FB�n����q{�B^�}��mK~31��i����(S������������34��~�����'�Y���:��#�9mfJ��sg�VЈͶZ���;��8�!彡��N���^�\|f��Ġ)S�u*�\���rL;R�1�ls��}%��
6~б2�� r,��K��~g��)tHa>*V�IcX�P�)|3'��g�B��/S�����K���ϔfޚ�c~1/{+"�C1�=�v��I�3VKT0c�=����J��Z��{/E�v�ëCB{�OE��T�횇M`��3]l�-���ˢz�<�_�z�6K}o�f��Y�l�&ٰC�p�:I�O5� �����F�]�/sJ9 `�9�*�6�h�+w�ٗl,�$D+���E;�9f%q��Q����oR�aV�B�F�#ݳm��U�惀���0��qS��nv@�:n��{�^i�p��^��rF���䭋mS���Qb�W@��j��ׅ��ݸv���:"f0��AS:�1׸�x�r�3�Tц���H��R����`�ϑU0s57�ş�S3cA�<�i�����f���W�nI_��h!��r^Y����"r>�6:��+���h�ݷc�uJ����!V�o��p=	b��8Zәyr"�ewG0��
��\cd�*��>)ݻW�-�����e�^��2�N<r��A&Lr}�J35�tM` �t����?�)�cR���n;T�Q�hz����0�����Ƣg�A=h8?�<%&<rz���1j�1}��,�~��r:P���:�\�n��ݓ������ ��!��8ȗ�4�=nޠ����K'��G���'Z��So��_�K�뱄����	 �������Ib+8:�u�<���g�n�ḟZH��*���AG�ՠ9p!)�, �~���af7��v&ҕ�8���} 2�mw�۸�694�i��
�5�QZ��I�+���wy�O��t�(ґ�ژ��P�$�B7�,�n:�m�L	���0���3���~�2��05NU&����
��Յp����|*;u�8*�
��4�޽�m�晤���v\�#>�Z��O���{C������3�U�27P�-��f֨+��|�>P��B��OPq�e�P��b�$#���F]�>0�\��G������Z� <����}V�ϸ�,�lu[
m*���Ň?Kc�~/6.�շN�I���w

2��)�.���n.����E@�8To�Bdm���hM��i��>n]�����L!��Ϡ��e{�"�¦��H=/1Z�hO=U�iO�K���R���s���g��;�1�*g�2�)W��t�|�S�
%֕��an��ܨ»�S���4�>��3