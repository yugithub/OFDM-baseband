��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�a�_[�c>p�6��?R�e0&��>;ٮ�.;�w��1)�ɶ	�!���<�-ED���_��Bu*��t=��3;(�����f�X��`��@���yh̻wd��~ȎT� ��s�me� B���`�?D3��s�L9�C��\�yka4	L�?N���
�']�fɛ"Y4�?�z�M�z�m�H��1���4�؃e/{����u1"��i����ďƦq �9��=��|TDc��y����%��4�0#�'o
(@Q��*-���X�ut�E]�ت��9VWߗ�����ɖ�%�T�f/L��}�3��`֜b������^2w��C���1s��DT����By�X��4���(Q`m��� ��H����X`��P�:�6�ӣ��.��60C:�34S�?��e�,\R�'S�q���+J��a���P��F�M�G�+�"`DN?��eSs"-�烶P�-E�dw��UT�
B�f}�H���F�	�����d�T!	,@��V���q��xXl�p�A���i2mз4�RI�^��{yy/3��8j+�K�����H�3��L��@��B)t���h����y���\�a�+��UX��(2�s��Y��D��R���i9ݍ�H����ũU�:C�Z���R�V�;�BKf��C�}�Κ��ҨУܞV
�	�;=��>���P����	)?/"}�]�/�5���~FO�^<�"��F��Y�A?̥/!�]�]�MYՑ�r2�#��?Ɲ�<�\p&����a_��rl����_�?e�z�6<.bZ^%�Qۢ�<K��k+u�e�M4h�=�=>	�@w����p\d$�@�X�AT��eKw]~X\X�wH͖mP��h�$��&$a.6+��n�l�8U�����Kz>@�/�x�w�H��7ЯT��t)��Z��c��������Í����G�(m'cr�-1hn����jQ{sA��Ar���f�C�RT�[f�����-�$P��'��l�~Ȱ�Y�4�=�	EF2�t'�p����d�5�u���1�Tw��^3�ѩe$l�A���/J"�-��+�i���5DG��EـO".7�L��Zn����
��p�'M�  ;�U����-������Z�V��6▽���;�yշ)H�0o���z�%g����=,�����v��E�̾����&7�2s8�e���a��(rŎ����� ���V�\i]��'_^R���iXP3��h���;.裯I#�Q4�(�C��t�|cq=�5f��Y�YV�J>mAYt�t��R���bh�Q5����5	$�7���-��娔���j�s����a��8z�ё����9bK1�Im����.�fȕ�\��z�Ĥ쁟���(�W���� �=�+�f���˥����>(�g.-$��?$ػ/!(�(�\@��帞X�"�v��	��x�[�n��k���V��<5ՠ�����YFAT��a�p�Zo��2 Ѭ�n�~��1Ѵ:sV�9k�p��
������C��J��k~�]5n��uM+�y1��B�f�q��f$�,o9�#�5j\mU_��X�"5s����p/�t�����ܢs"?@�����$�hW�X� ��� ⼭T[)ϻ�w����--���4c648~���ԉ��@^2t�W��7�H���Ģ�����;~�#��Y�p`�{�? �����H�1T�*j3�J7��F����#t�8w�#ɼY����Я�����(�Ȁ�/\\��V�w��[6O�� tz�V*r|M^!\S�+AV~o�q<�����<�����'�bN��~hz<u�QM;=�|��x��s�sD.`���yV�r@�U���!~�wm�IW��������ˉ�P؝��A�
�S�Ŏ8�b���3�< NLQ	i�z�!߄|^�~:(��S��)��ׇ�"��'G�ӧ�a�?���W^sK�
�;�1V��%Aػ������!��+wq7\"2�E:iR���� N�;/a��	������i�T����z�WS�[CD`���;|���ZxN����!�zv� �K"�s����[��v���]����E��9�_�i����v�p�Pz�X_�����ʣo��q>�0��#���L�q>E�t��I;������a�B��Y�F�3�{�7���̈́�P�W��f�):|N���.��Nw=�c0,!��;��L3�l�=��V�`\��x���?f��&��{Y�v�~�Y:t{_[*'�h�򏱶ay��8��T�����Qk�P�w�3��IA�9u���|�;/8�pjQ�_�L���!�܌�9�p�8����Pp�j���?�w�a�v�e=mN�0��25g����c	��Ϫ���uF�)�H���^Kv�z��H.��{i��@��\���f��)���hC)!�1��!ĭ(�Կbɖ��\���}�%7ΕI�b��S�od�cu�iH����N�l�5�ǀ��|�Dyڀr�1fQ0|�S6w��nT^���!���:�`t�T��K��1�P���-%D���j���VQ^:5 ݸ�ֳ%�2 ��
ǘU-^QS���τƆ��
ߩ��+}6WĂX�p)�>d����I�ROdȖ���B5h�P�FҰ!!~&�<�q4�~��/�]6��c;Ґ[�j_��oE�"���rLץr� x�c��y��f��jdِa�~o%O���ˍt���f���X��=�aG��;~Fߙf&����!�fC7�^}�%�- �=�W�:x�I��2 ��]���K��,7���f�0���jw�4.�<ϴ�r¥��<O��B�O�ut�j�!M�\'TjG�I����o 5�^ �w�o�κ��}&(T1��+9�њ�ؕ,�T����Ӈ�H�DL��|����Ag���Oԥ���Z��T;Ҳ�D��L ���ՎH���(ϊ��#!����ΰ�h8����s�~�1����>7�Rۧ��H�C_}�=���%	������^��I���T��	Z�&MJ�t���u/�Y�#�W���1�;R�bl"=�O`�y��:;@�Y0�J/��7���B�Q9#4�����Q�:p�f�����N�[|+?��s�؎�����0�V�&\n����9�jRD0/���	~��.�W@�������P���u5�����7�wW�LbCm�j�.�Ї�.R�9����xx�'�.�"Ok�o��R���q ޽*uO��O����v���y/W4	BHM����G�$	�6�l2��.!%̕>H)��� ��.�����=*CR��&�X�V��Ϡ�����1(]�����������l��"[����EsS�$%#���_�|��	�R!�(�鉑�\��>w#�6��$���6�i�l 6{E�A���\D��1Tc6�X8 o��f'˔��?2�O�%������˲0m��"�ue}����\+Y�>C����~����M��'�
p���J�wMw��Ts�P\�\۝��Gv��Jx= �`��I2z�J���t�����+rԷ��w�����XȲ���!RU�%_iي�Eq�T�4VTW�Y���X���W�I"����]�b|������9�h��>���ص�/�x��G5�i�r;�w���IZ�����Χ����U���e�����>Xz���F�!�Ym����Dm�{j�cf齳қ�!��-�Zh�c����蝝�x����2����VA��H�w��t�ߦ�Jl�2ĄrC��
� +��	>�٬�8��!��χ3�&��l*]�Źsth�Tщ��!�h/isޫY�v�x���m[�!�j�AY;C�<!7���_�8�oD	�?�ţ�Á���t�Y~Z_,a�J�W~���X�X*�i!!��u�����|ӑ���Ë����}x�13@ȔbA�M!��k�QK�Yߎ��ni�+�:O���?ݽF>e���I���NA�}2~���~5�bX�5ȭ��UՀ�;ȵ[i5j�RL��]��1e�v'k��Cv)Ԙ܅sP�fQDn��
�{ �
;k�4KR#��d���� 괼H�!��E��H-Ӕ�Ñ�Гo2��u�9�d�"���>S�� ']���W�\t��@&h������C.\E�i���Ձ%s=��#�5ϳVZ�3K�U�lv\��[mD��r��X��Yc]/�*��:�ފ)����Л�����/L8���s�.����iB�㘥�򔜑cS~?b�����94�{2�vG�����@n�)S�<9��ӯq����N�b2�Bco8���Vl��_�c�<l=�@�z^ߣ�h����?��T�c��ɨ��6��>
���.B�����*��N�{���C����qsd�9-��奄.>�Y��l	ا�h���j�fY�D����:S����Z��ٰ��X���/pJ����Z��������š�y��H�����	)���Tz\B�4ItI�R^_�
�� ��\-_2 +��>�@#
^<(��g �G-��1�� �뫠�\�������1��ٲ�8B�`��!�N����Ӆ���t@0/�8���\LOc$%.��zAq�Q���y�������(����RvH�O��n�igB�a=��=���K�bN���2�"1�Шnj�j����uDn���K@)�$L���y�����X�''O��kly#�#��ʹ���<0������:-�Ε�����(i���Q��o��d~NR�i &�uJE��>�Q���
����K�4�rKsJE���f�P�B��J9��=1aj(}M�)fV/�nE�^H]��6���Bk{�?B}�Uf��u^��u�B���^��!�|P�_gcq1��K��J5�`H��M?�j=��`�,rُ�����᧴��d)����C�ɥD����"G )pZ���8�0���2h���+��)�pjA��ZL��3�z�v<w�lzzy�ūT����A��2��]�x} �0!�TkQ����a ���+i��?R�<R+�_��U䮆^Zu8�A����Ν:��n�=��(����ې�Ü{b�N#X����V����d� ��2�'�5e� ��_�3��2.D�7>������� &3�x�g�ؒ�]�\��[qo�����x�nC��������?`���o
��LY��灠���C`�.$�\g�����7�iC��)����h��)�����ȹj ���fD��\�����gcM�Q��յ��3��O&�����DST׭�\��'`�.8+a��g	�IpL�������T�����wI��e�+X<�ۘ�A��2��z*�gb�(�HCu#�c-`����jxع<�|<@�-��?��)2 gJ&���<�^įަ�h��a�u�Bc��w� ��4҉��V�,J�6N��Q+w��a��O �p��k/w�D+x:u��j85���o�<.q�-i�_�7��J���8!�)
��t�n���7WU��Ʀ����ǲ��� d��Kq�\��Ɋ�CU2�SR�r��fD�%�|<&��
��d����vA)0C���������jm�kWY�J%���m��'8�L�jYYJ�Q���0ma��}�F�}�CM����5�cWT?�9='?���3���jI]?��q��
��ڽs$𰁂�����+~.��
C�b�JZq���dfʇ,-�&Ѣ�m
}��X	�5�#�P9Y�~Jm����A��J���g��/X&�|��̭,���Ҟ�S����Oj>QR�O ^��{�`B�Y��y[\F�`�*}�-�("_�CS�+�Z���L���Q`~���K�	6-�m��Z�O[H�L�%�a��o���ԡj�zʹ����?�#��y/�+�օ�yao<��LWퟛuiz1�Ӹy����c�	��(e���q�`�'9�DL.���N���sўz�R��3��������)Z`N��Oأ��y{8�I`���� �J�3�� �{l�2��~��W����ī1��?�ژkb��!��cE�Ne"�*���5.L����
�!���ld�1&��D1]jZ�Qx�M���Wh�|�ʌn� k����/l����%�Y��w4�+r&ۄ��/xpN� 3��� �^"eǖ-�J����8%暝��*]=I��+NA��Pg�$��L�ߗ�1�H�Z��}*��c�ߣ����.� �v�.CƋ屉�0A �ղr�l�#����:R\�I�X��%Wp|�E{��@�7�'�q`��b�"\ۿ����%����]�<z ����ddf��Z����WB(�ܬug���qΓ���K�=�y�q��,��)*��v~uM�����xԠw�3�	ޯ��a��7�?�1��S�����㐎2of����$��f "�)���#M�M�Ub)|��Ied��D�jk:T�Ĝ�U�l�������U���B�"��vr�-�9���8�{3��;|�W6���z����8�w~^V]{��6Ve,��{�ΓHelc
��ؤX
�J��%��I��'t���S���(�߰��,L�'7�4�+!�A;:'6>!��!��@AT����B�n�؛!��/y�9,���l�H�����`J>�8��m(��������*rxGa��[HG���m��5�\��1jW�uD�(�g�W|�0%h�8�t���a庰)��%��� ̟�g�Ӆ�bnܦs��<B�?�ۚ���S��V�����ҁ ڨ?�i�����N0b�R��O�?���m���=�&�S�]4�q~��d�5q��ܒ�R/w��Є��?w�/�ƴ�+�;��S�����|t��t���!��9�!U��o9�'��O׻e�VH�DLO�<t���w��.�{��P�W��M��O/�����1��UY�4>	�n��[e�m5%����A��kɏ�V�E#B�R�a�l{�o]K�[�<�k#\V�c�o���T�8�7~�B�s{.]ftw�����p�	�'3P�{�8!K�Wg�$��?�d+G5�K����o��b�!��mk�ep+d�a�)�}|Vd��(]�n�Ӄ�j��lM�Վ��f�/a��9��]�i�4,ʻ�W}�;8��n�툱�8\;�}0Y0�~�e�0V
gֲ�}@�}�t�i����h?�i'v�=�޿��db`���[�T�w�,��0k*���n��]rd��a:t�����W}��x}��ҵvo���F�S�_��\!��z�ټ��Fx	���N$
t��=6ªI�P�%4���w����6�Nη-+�~e�mx�Z�+?*V�a�0g�ɵ�o�w�h���ך�rW�z��U�V�����s��˱�)��Y����}5>�Y��n A��|b�y;�lC𚨟�����47����b�΄p�f)D��h�g�ei�/��g$���p/ƀG��%� R��=��55�	NlD�����J�m��BUթ[���>
8�ũ���Cpժ�Ur�HwU%�)#×lΛ�qM�D�4��L׭L�E�=�W-��m��g`�.����r"�Ҿ�ƥ�h�k"���{�w�W�c�9Z��{Q�@��q�M�cH(�#<	[�޸�N�"�p�=��>gA6}��h��D����U�m\���NCޔ��w�u쉷���`Iι��yj�,�
2��5􈣃������{8�0K`�sb�V.�A�m#�`B��Vd	��ϒ��+�Cɧ���7�:���i��~k�Vޖ�>��eLvO���?����ِ���d�]Az�Q�-A홡�7t_1i����Vuo�S�a84�%��<ei�˽L��\���ǋ&"pŗ���g ����Lz�b<vM(�~��O��|i�)�H�7Ot/����R-��tk�נ��[���8�Vi�Rx�p�_@��6V�B�4#�2�{�Ss�6�=���,B�8�I�o���y/�1Ueоda�}$9�j1R"��ᭊ>�~=J7Zs�2� ��@B�E9�.��,�P�E�]�'�R�����F�;M&t�͐���H�2���cxV�J��L�!/�$!H�ʘ�>Н ��iB��p-�)���2��HY	l�v�H�������5�;�-���Ɲ�(��%<��1MPT͠�b�8t�YҷT5�vm�al�7�Y-��T���+.�����@7L��糫n��8u���d��H��Z0��I�(����¨�S�Mȝ���nQ�[ǯ�����?6u��aM��t�^�M��X;&b`�v^�{4�F�kuJ��B���@�����[��{����-%��͗,��"�S}r_x�p�aeژ�c�M�\hۂ�䤻�Rb2�,�*1�d� ���F��*�eҴC�2����i"�'��C\�������lt�K�Q`�μ����
F��2ȝi�@�N�GZ���'a���H�������cD`ͬ���0��}r�,`2O,��#W4�t�P��e�-�uM���f��&-αyHJ��oB.�$3�"����I&�EK%3M�l�&S�O m�ޚ8H<��x��
6X;?�y�)`�v�ܜ�-Qj��֡%&�<�F�����<�� �N��i~Vpu��JI�޻��z��(�Gz���;��ѠWe��`Ȗ����1�����$��C��?tآ�0�ͼ��Vq��e�!�#���s����$вU>T��q4~k�������ž^K��lWK8��ˊ�����W���fAq��w��4�(D��P�����ЭxPx�����I�/�-��N�fMB�C��2��Y���Y�]Gm�����+	�3n�_E#GK�5���m���*"���rhA�4*��� FJn [����.cg8�a�a�.�CJ�O�>�e�7��4ߞ.�^�7 �1���Nظ�|k��g&�_��.#��7�~"��J�YͮC��Td�o�p��h���`N1�H���uY�L@����dN��q\+��7lE��*�Lׯ*sk����塩X�G��NdG�p�%rb�(a�,� ^��OO��C�i�[�I�=/���wV�����`g֬,g��zO���f.M|~O�/���G!ډ��3*��_����Ţ��)K~��je�����(~�r*~x�"uZ1��l�"-;���T��n
PB��Z��t�Ӥ�ʙd��^Q2O�a���氏Ճ;�eޓ�*`�X�[�ۤ�Ԟ�7l�l�"��%��#n��W��(��h��'RtZ$w=��HmS�2��A���4�3�u��n�a/���Ի�)@�7�~��Q��$ �|e���	d��5�Z�ol��N��*�b`�^|�E�-g��ڑ�#�г;�^㪧^/�W�'��عG����{Ft�K��y��JD{���G0S���Mv���Bgr���FH����G�}
�q�ċv�{�uԡ�W��/t�m�L���� wc�q��`8:��Q�v�>壷�z�w��~)�w[���=�/0�� ��L6�Q�� e��=���Y����nf2����΀�� �o<�J#���;GR�agZjVК{�w�Ts��E��7��B�8��6׶�����3���6��8�����L^&���D|����A?�A�n�_L"���>�����5t_v�q�;�N�%�$�b����i�N�H�~R:kJ�tтYן��I-�q
�P�FJ.f� [�⺵m�},����XXn�K�X�f����x�����wdф�����2�n��I���R9��Jc[���/���z#%V���q!���ƻc�a-��[w��8��D�ug�_��XϋR��?��j&s̳o쮡��awQ�_�X['Q������j�k�H�N���7MY@���<y��>K�1�������%>��%��S:|V�F����q�|�t ��X@�h���������c]�5�$�����:���TO���`��_����,�֊ߟR;��B�w��ͷ�}����x_�$�5�9�:2e��J&B^��w,�x��k�kȁ7si�8�� �["x�m2Y.��3��c�#�&�I���Pdj۠f�(�,6��f�֐M2��Ǡ:�:� ZV��1\�BS�({��)��ItyC*Z�� ~K��؎e��/cw�ۭ���H��s�������Of�'Zbe�!5�,ŷ�A��ŞM�(n��2�q?;k�������&������Q�7�ج|�6�9y����l'�\���άx�����
g�Z��8���Yt����Isű�?;���Ɛn����d]����Ld�Ɂ��d�q�y}���Y��������y,:�M]��/ �z�����'�}JyxG܉�n�ֶ�r�֛`h�>Q��Yb�����r�h��F�K(Mm�N�$!��4��N-���rSRGnB�,�V��<��*w��E���4횝���N�2��!��$�=��i�J(Zٴ`P���D��B1��`����<�m�0`�����Ԅ���92G����%H�9Hp�6a�\��ZSTq�#��m��R>�N��RF�·���.u� ���Ty��7 7J&��, �����Y���!֣�F�[���Y��pv'���=ꨃv'�\�}p#�M�((�9p� ��WnN�t������@ʷI���b r�7�6�H�8���-�5J]��X$&���r�B��ϭݴx�+�Q�������@I����T
��R�_AKH�)1a�{���w^lK���EHV���!?���+İ�az�Չ���)3��v;*��w�{�j��޸oO��"i�^�`�r^�Q�K�_vX]�kjc�k���/%pN��\P"��>DAqr�Eu�m\Da�4��f� �ɼO
B���yksNZ��{��fwt�j�+
�l�ٙ���B�DY�����'�:a�nUr�gS��0P.��t>l�w�/b�(Q�6�>d<8:(/Px:�	�L�+�U6�8�m�Z we�7ӅeA!?���4��,cͰ�de�;p�Y0�3#���T,7�z
I�Q����H�����w�`�x�W����Χ�?����O�I}~qʊ_���r��;Tx��U�#���jN+M9��oF^E(�3X�a���|���z!.�_ ���(��Ǐ�'�9�*�3�Q��1�p�F��$��j�f���3��(T\�&��s`����5٬���;Qu���%�DM��3�z�LѴ���P�1�ގ�6=���j3��FwjY����.��C�e��c"/�$�������u��2��%�l��)�2��qe��.�-hc�d3vrEk����"
�����C��5�eq��{<(^�P��ʋ�L���5����!��[bk�Ȳ��ِ1wv$���o��H�@�#�R�M�*͜C���ʎ�N��%229׳8�v���z��	�0z%Ф%<m��v�ٻ Y�6d� ��g�D� 6��V.3����:ѐ��\��K��J��ք���_��T��]�ŊC���fF���BJ�ҝ�r��.i<-��\
l�uI��R������ʺ��z�m��`�`��O-I|j�*���%l�1�J�L.	���țʝzV�)6�5K<}@Y�M��
��d�����֑���H`4xA����5g��U���ee���f�[��j�֐/K�*Dh8��j�i!���ʰ����O���t��cn����Z[��v55b�Y$���f�H34z[�����n|��Ԫ��/���3L���ST��}�UkR���O�!:i[$�Mg{Jm�bο�Ȼ�|jz�u�x阂���!���Bl��63��^��~����n�z���p!�c�Y<:ab�3�&˅�?M���CWBB.~���M��Q�
*�1�9hOd3�����Bн�̵�Z;l��Iq�%�	�H{fQ�o��/r����;5-�J���߻��!��3����O�]���}�Q��	�|����{������%����8fhγ�	�h��}#��#�f#tN
�dqG��t�-|�u�v��80!�e�U��ﴶx�,Oi�Aʖ�&��B���H��Y�=�X\�,��������~�®:�Kee����RK��-x���$�f�v�t��F�g����q��"�(���x�h�q$�펁�3�5 x\����#&D$���u�?N6A��`�{��G �T�ߕ�@��m��(|St2 �=J^���������$��Kc��̍xL�z�%���E�
�򼸻�&���ZR�<U��N���$\�3Z����!8��uS���[�f����[�y��0�O`�G[�L��<��iYP�+;�S�pea��e܃)}(>�@�'��U�,w}d�-�*�+v���c�x�B������.��Ͻ��zYtC ~A�]�\R�/Pb�S"����Ϝ���+��Aa�XX�$��Q32���·u���ˆ��+��|	�,\���Ax�2 9e�	�o��uk%��<�g�2����Z�ͷ���c�е'����lnmB�_,t���[���F�Y>������c���G�C�z+��N|J�� ݼM�y��A�|��i�R� �~�~�S$D�Vo�ą^��{�L��X;��I�]��JvZu�p+��.e��i 2�c���C���@(2���?�7h$�*|	J���r�E5�N[���pk4��Mk�&G7s�2�t����1�&nC�+�ǋsz��Z�1yG����"�c����_ӑ�N�"�j�q�A��J(|�\J�k�Yk�/
XH�lq �p!�2�ƀG��r/�xE��,:�^�X���kXP�XK�d[��Fu����b�ͼ%�y��\vq]�ASB�}�|S�[�V��R�C��#>d�H�2�#u��\����mM�_0�- ���r pR���R����eb2�>��~�ujæ^iΠ ����/��6J/;�a5�}����� �F���,�x�=׎늕���r�ʐ�MN��s����H�:�� ��ȡ2}���[���L�+N�c+��i�ݳ��.��Ԟr���b?E5�N~�CH��L	�2쭵@�EaL%�!���3���l,�;��i&�[ϰU#%�����r^��5Vj1���__/v`LeN�����X�����c����vݏ��9�|}H�n��*b��xF�S!&76{�9�J��A���0�Ϗ�L�Ǟ3�5�a����a�I���Q*��z��f���~(�*�Z8;~�� &����?o��Z�� ���蓝?:�fWG�{rJ�`�~�?荕�}�S�ii�zWg3u\�1O�� ʬ̂ﾎ��4{H9�0�\�[����#)�tiJ�J����:�֤��YEV�Fl�YdLV?Cv!O�:��:��(|�������L�8x����2gi�q?S8�4���9��W\)�\j�^��m��-����q\�Yk'f,[G�q�4�%&�q�W�nq���/�^�]F#�m{��;�k
�$Mu�Ǐ�M_��wvg���̀5�y�nm�:�w\ƓrWvI�����Z��:@�QD�Y�h=����4pCD�C[��<W�h�0:��`�g��oB��fV�dʓxȍ�¨É�y%� �G.�S[y�Ƌ���j[����ϙK*;;�SW^I(�{�f�:�99�:���A�@�oxjD>z�|�SxW|��&!��IO��u����9fb�.��S#<5�/8{�E3r/
x�t��Y)*�/��"�)��b5�w=�Й>5�uL���U:��0�)%K\�����"B�v��D��Ah��N�)��RՏw�
k�t!I:��ڬ��+����6�B\� _��$�ED�兛� s
���{Ĥ��H/�y\67�R�y�ȭ�Ύ5D����˂��c�;*S�^�Kf�޹2@c翐��0�bK���I�x��T�J��(�7������y
%BT$A��tK���K`�nO����<t\��j�dS����uV�����Ȑ~��Ao���L����{M51C�W/��P`8~�2ac��N�Re��k�KS��^,�y�Rm����5[������Gf�r�=�pS�ѵ[:p�M���o�:Tz���4wN�/%4���P�}v{G�s���)P�G�R�-T��ڸ��{�]��$�J���y(@+Na�+�_��&+m�N��x�<�}��:��n{�,�^�퐶Ց�c�&�FJj8���z�\!x���� Kd=)%���T.G���_r��P~�c�8̷��)�?:���S��A�R
;^:0|�x��[<�G�jح�}F2@M7Tw��v��ִw�gX�%����G�93:'ũ��.�2N�Z����Z}	R���P���޵zfC��EGhc���~T����ю����%-,$��%gf}@Ȓ��'I��v�r
�;�c�e$�������ڢ�Ż�|�V*���U�9�!��6�K���V��և]&�ob8XY8�ɴx[���(ifɌl�+�ߞ_;$�ݞ�m�,�mip���\(I?X���94ӱ���(�#�b�Cޙ��)dS�� H3����1����3cw��y"(�t��)�Sl]����o���a�� ooE�d��OK�P��6���V>	��f���麙9I5�[�D#2����Mb��T�ܘ7��hX���ε��u^#3_h,!��C^g���|�>�>���@�Q�<�N2.�8�rv(.�Hc�̢��N���3��c��L�%���D�l�@��m�� Wʹi�}0����x���=_Xi���`y毿��(�����"u��<�
@�Sbŧ}�Ly�:A�:p0?,��H�i�2�ct��)�-'}
I*aNIM8׌�2��`�s�T\/�6qxNh���UċZ}���_E����4&�%���)bp��O�P�g��\ě�8� >RIB���Tv�.2.�����2�	g�>�C�Ѕt�רd���:���	`ރl�V�6g�~_-Q���3��l#�_ޗu���=��a�f����ʋѳ�gw��n�'굢a���]�m���"�Q)�*�I���y�du����Zx�G��0���0b����?����tUa�R?��ߴ_ص�I��U����t�7q�Ob����*F����֙�Њ��PUG�uM�w�E�W$w�E!|¨a���������C�g��ťh��Sg/�̀ٱ��(Irt�tq�FE����ē��k|c�T��q��<!�k�G@)�r`���ED�5���6^��Q�x���aHz7�|TX��O��
f��^��aw:VT������q�Ԍ9*ŭ�z/��sC��va�IՕ6= bȖ�s/>�d�W�%f#K�ѳjG"��^��񄌑l�a����ȪF��-�¶Zj�8�9�D3>����$�><1���S1:l4&�Ԡ={���*��\�^�/����bo���lh�W��JX�`���_<�x���z�" �|��6�����N�/��� �Һ���N��Mu[:�	@'W�KC?W�:��	��'�e�˗��	&��MR]<��c'0���)�<_��c6YvO!��X4E8�u�LVD�#��h^���7�1�-E��#Rs���4�@��C2Პ�2��̒���������|�6�L��A��8�zn���,�Y9��z�7)�w �o>�=���;�� �0�T���+����e�4�[��,K��k�R���G��䏯��`>���n}�UF���W�1�4���ɽ[A	]��6l~���o�� �<�k�a�>���H�誾��]��v�X� {��6pZ}w�����Om	4"2:x�"3)K�(%������y:$��T@1���]F\���8���C}KB�P���<�$�Ic���X �d텓��^~K�S���U���svR��0P	7JKpI�hJnt��f�^�<��Yu@7���"7]o��м"�GM�3�c������l����W�"�Dt�&��x�r�A�V�Зx�(�*^��m�B�5�I��x��v���\ȥ*ж}1��A�#����KD[������L�݄��"\�Y�&�W�gY�iT�j��;e @�Ƴ+�������G�R���c�n)�s�}�����B1�tL?v�Jh�]X��M�1�G�4㈋�XU@@�6<�eÃ�[O)Q�X5���g��r��[�v{�nS�i&L��ԉ��c�q���T*ܷ�U[�K9p=�n@b&�s��[9���֗���؝Xp�B,��tp9��
��W��! �u"�?|�Za�~�;aӎR<�Pe�O�vI^�.�Dn"`��v���!N�����ۥ�UJ���5�e�}$}On�N�?R��Ю�t'�cj*5�%���.��v=�{D���uC���
2=�M��R}��h��ٙ6J����-:+ ���s�jT�;kUb�l�W����3�Hٷ��&e�X?m�'��.D���+k0��	e��h_�*�f��Vz��/��Z"#|���7̝�Q��!�CE
n��j�Wr��i`wuN��`��+Kb$�D!��$��ݩ�1��7�V�-O���0�������,5�ܽ�q����H�tp�Uw��lX��eF����>y��Gb"�P�N �G�$D�����X��H�H��p��x����zव��3B�2�AM�ڶu�H��`O�;_S_#`�* M���"x�ǣ-�RjʧPb&S8��D�֛!ݕ��q�J����漧u��c��[�t(i�{�c�(�����&}�죶zfT�����u��R�N�a�h�\��R�z=7b�Ls��^����<S��Rt�m��Jg^�����'|Yg/�a{�E�X�8�w��˳�T��ո���]���{�*�>��!#�l�y��k�.G�a��FLy	5WQK���\*܃@���q�I���,x���F[�׎5�NA�9L�=��u���!r��l�؜2e`ȫ�I"��!��@����)�����`��6�QAF _é�,�ù�!����,��/7�[����\��sn1��O=3�eʌ�L��Q~��G�E�M>�)|�%�s�I�`���^g���Fa�*�KQ�=�������܀��o�G�tʹ��*��]g���"������!����-���3GD�ŝ�p�N�Ա&�'5�,ֈ`a�|�%��b�L�#�'�����ҟR_a�g�?��$Ĩ���Y�%^ !�a�t���q�)��h��M���M'��۹D���@����3���.�ԍ�4|n�C��bc��?�6�9*�|�3���aq���~��Dw��<�\�L�\5L�ko��Y��tK�88Ij�J	wfɫ��˼hLЬ��Wۑ-�����
!��dF�@
-��l�)����{[7Zp*u�#�pj�;yiN�����뿗�p��Rឦ,Z�tn�6� {�v[z�����ѱ��q��o �[������0�(��節�a��΂֦�=Ee#�K���O�T����l�-vkD�F;������C;D��H����cg�����'4�-�ղMGA�� ��*g�6������oT�OM�>�_���E/�~ׅ 1��+��h-�|�>��'�iZd�FOI�\�9ܫ���c!��3�v�2W覱����YN$u���3�3�b�~��+�X�����?���}GTb5A���Kp�7Vy�61�8o��ǑKW��U��� (�^x���Ȗ|L��&�t�:p�w��ԌÔ[6��Wl�� Fc�!�\�_$*��\u��Ɂ�Ms��"Y�lt�S�K��z�[�L��Y5f�i�%V���(�k� \y����.�����4���w�ȅQ�Uc��mn��	�xP��O����&ݔ��\���XC�Q�l�-�ۆ"���t6���ų��*kQ��c0Rc\���v�z��{�7�[i�?8%�c
�{䢤&�
��BZ����~�ް� UKLgG;�oem}��t�2�(���Ku�b���Ld�[���fn��"/"�8�G'�Π?�2�R���Ӧ�`�h�`s&�f�B��u��0��0�n^���U�L F|�V��c��fa���G!�bF������x�b��@Q�J���2W{�D��6��������c��j'Ud�씄:n�MB'��/}�\���mL��spASS˿���% ��R��R�#����Bw!h_�hOߵs�B�����G��R��k��u	�'4�x`�x,
����@�<�]�g��`���^�%��M�Y	��������'��&�8d�2��/>�0���R����{���|��hR<R>CA���vʘ�p�r$����x0s�W�P\��Y�3�	���y+r��Gt�Yn�'U����q���T?u�Gxx�+�4C>}���yH�M;~W��e�TG� &֧���N�)��'s�T"�	��ͫ���1�,�%6��;�R��@���T���e����r�����V.*{��|S4/[����h��5^DHm5��=��%j�}{���!,�8�Y���Bbʭ������-���LU�%E[�mP��'���E��l��_{�[��+Ty��z�:�t�q��$�s��(���T�/�(��b��'CD�fФ�qؤLo��C��nu��/,�B����åCXR�p
yj�sQ!du�1�%|߄�F�:�/�;��#ጤ��\<�=,�Y���r�8����J#x���v��҅q)��B�6c����*�~�oG�a��`�.d�������^�ƤR 2�AH@��,�$g[`�]����3SO��¨�̷�k����U���� ���g�&	'׵@�lۂ�K�j&UH�H��!�7���]t�W��xԒ`+�]��^k�o�t4bߌL��'n��5�ȍH�l �
�5�\m	{*����ۡ=Ū�LN�kާ�IB)���v
N��6( �G<�ÙlP�2���d�Ί�*{F���$aӷ@�|t��>d��E���B	ag�j��l�e�M�����V�w�`R��hʗ[��^m.0�۹����'�}��d��c����t�uD�Yv�/��g�k01������ƲYb��Ŭ�:�gzЅ�\҉=�
���ٝ��Z4�E�����q�l3�S�/�UX�Ǖ�c,c�ZQY�]�����������e@��U+B�Y���{�:���m�W��2��4�J��E )4;q,WMnV{�|��Þ�xa��{U��9}9C�,�FsO88��H�8����kg�9��#1|��
�>cǍ��c N�+d1IP	Jdy�P���~�������mSJ-sI��<V~�@�{����!փ�]le�M!�id=/�քv�N����L��l��G˾���҄�����G:*�6.5����[*�<\��NvI��� ��\j3��h!�f��Ea�nǶ
*�+�+gk,��J|�Ǡ�Dl���4�B4$���h�dM{5Ķ����L&������j	C�����YZ��VnpUoh�q��a�cgK�Rq�c��������rt¨-��'�E�����C�%���!i��'"a���f���G�8�I�1(���h�)�<�q&��ZO�ʟ��ۦ�RA0��A��Q���Ho r�j���.�Ԙ{-bՙ��FB9��=OIO�J��	g���Ɲ������}g�*�{,H"<M{׶W��5 ��=hu�킷s�Z-���g�����&S�,��O�~�����켚oQ7����G��7��z0���a��D�
������-��G��|*˧��'��J���ݻ�r���b��܉+J�G�4h`ߕkk��+�+繙X�V޵˜���Ѧ���T��0���N���샿��x�ީ��Eg8�8���V4L ��OD�A�c�H=}ն�Z�?�Sž��@�j�}Gq�
5&*��ӇGX>��a�
?�Tn���$��ox0��Ծ�_-¬!�����k�<��nP/��uǂ�J���퉐�gq�u����h�6o���II���qp}p	���N�X����Hv�D���v�V���W����b��o��ˈ�
̻�
������
�z���[��bl��qy��)p+V ��d�
+
�kq�)��n�J�2�e�Mƽ�r���X�zX����֭�go��a���Xږ\��#����6Zx����nQꋿ#�&�D�п��?#-�^O��ގE���Dg4U�%��$�R�W�6&�傗����e�P�.�ʭ�,
s*W��ax_�O4
J�^��]�*>��zO�%�8[��>�������䀅ٔ��0;�?%�P���?�����1�\3�����8��x5*v��Q��9�r����(�#g���:����+|?)�`�z�^,���9�1>��i��m�_2�:L$K�;b#����AΚ[�"SW0_vq���Bf� �us1+�c~��
������w��<c���o������{�ĞV�X�}Ec^�P,�&#��ڼ�D���úA�շ�C�U��ߖ�����a����f��3�Ϋb<����
�P[EP�J�÷��U�c��א��N���:���y�vA9���f���	`�L�	K��� �#'�b���M&H�s��.̿=�=���A�L��V$��uWT�7�?Iu��K:�f����z�&@��.isz<� �A�"�OÃiJ��7Nh ��pV����
i^x�_16���e�͐�l��#'����gY]��&J�!E���P7{�����;sV'hܔQ]��7kw�B�$���a H㮋�O3�*",���Y�j�| �Mx��3�����
a5e�5&���N�)<=��_�[�h����{%�lm���v���?�[FG�/�<e+VnU� ۬�/\��
eӵL=��P�e��.���:|uI�W��5�-K�"�.��K���ֽ�hO2mz0�hPe�(���0Zr����&]6�`wd�w?w�0{xB"���8�~uضt�Yql1e�zH�1�@#�[���F~eXq٫I���e���@��m���<҆Ҏ�KP���fR�4KT%���xl,�5��J�N:������o8�Sx�ț<j��� ͅ�>%��d̦� 	W2���I������P��<���	�B�!A�>h��H$\G��U�C`�w͜���X�	E3l���7Ѵ`�F�xY����Y�����n(���e�[��8�΍"�k>.nyG/�i�n������0�K�&��b,-��\�Sa�eD�ؿ/<6�{�����N.��w�e�'�k[�f<��|���(ea|,���]��+v�$�ᄆ�D��B�y��u�`}K���H\����Q"��|E؟ܫ!����0��C�^�������Hm�W�J�ԾbǛ������{�:&^`v���ыk�?�;�7n;���>:��զy7!'�B��Q3�9�1D&P��O����nZ�J�$�.ֺ;q:�������A3���(43�ofT�V�8ުCW�k"�1��ۆ�4̙� �Ϲ�����]�}�IG�#C�9Y�2p�lY��6��@yߕ8Ԉ���Ѯ�mJ:!����}+C�B�|��ZKi!^h'�* d���z����2=hV Y��e��a�V���2K���I"��D���Kl%��H쟲��1�{�L��0f�~B���t.�hA�#��H�O[�쀣ˏ6�MX2"_Z�x鶑�V}��)��.,�$�/���g!�*�����b�내�k)�:��}^b�'��WEV��LɱA��5P��:�e#����d�?=޻k��b�����1�<���f�v����4G�f��>�y�FK�I֭�"�nX}�'��%�ǹ�ɥ���?�ޗX���dw���k��r�7�(����j� U�T�u� ~��FT�{�
��b!3�]��˵̜D���pW�����ի��l���I�K(`���s�ʙ���-
T7ףG��/��/?��;��Tn�`z0��3�>1 I�A�� ����ί@V�=G��Vc�'@���W�r��P��#>���Uu\k�2y�F�dV��tOR���9=��t��dw���-@�|�+D�;��<��ߦ<��(�]�_#�8Pæ��ك+����AV ����rhƷ�I�a��7�K_k�2�(���}���������.��RDOA�J���IÓ�8�Ӆ L+��h�����~��lv#���Ƶ?hg���bf��p=\Q�
�銣���9џùzn���2:ݟ�|��#�t��H}�����D9z�)��T����Q�v.w�]���0�;D�<�Ia���g~nP�qWAEo���Ӧ�Xu�5���SLi�F|�^�^ʪR�;v��D�/���8��ra�������)�~Ew'�]�V꼜� 2����n����o�;�7�����"��D���v8���7�|��s)�|����Ȋ݁?�lM�7P=�׮���r��#bIg��/�j�.;�� 띁I1|� ��@�j�dm�u$�鬤��}7�|�n������&�\wB�����r���T�Y����p�r�N&�9iQ���Me�����T�mt����s١(��J3!��@�s�?��
�[d)�[{.�@�ڤWg&㋺�	��c�5�rGo)�Td�p	�-~.h�OiyQwZ���꤈)�B��v�m=��Y%�x.�%�4�o�_Eh\u���v~sO�� �sZ���;�h�3�?L#A<H�rn_1��Z����)�-�����Q����잨�Q���ق��D��(�y�7�#���Q9�tK��,b�_ H��D�t�W��I�0�C�r��s�P*T<��nu�o���Z�*�t
R�"w�N��oP��.+�}���Y�c���Kn$�p�jp��[���p��<��;8�>��W�]��2�~��k�ȤA��e�.�>�x7�����Q�A��<��~�ڃ�0v�<�9�d	d��S&_F�vX�s�K��-T2��8'\���z}�V����`.M�n�=����5��z�խ_�6�v���]��&�uٵ}���ÔJs�#abY�$b)�f32���f�#�Be�Yl�Q�Ađ�r��$/2�C}O�?NMQE����1�mV��m�'j! �ir�ƠY��W$�ِ�p�M�_)�@�)�اO�[�T[�.\g���]πnX�O���:M���,��`2)�.��#�"�iDh����,��!'it���b�WUeT>Q�~����%�Cg-���T��jX��~�c�<�`k%CZԯ�q)K� �kɁ�b���mSG,{�2�Ci1�+���n��v1��d'*NV"7��R �Ȅ����WY��*M}/H�$ͨ��n}"��f�k�|���Ǻ'_���l�9�{�P�DK t��7�^!ZP[y��	zSHW�~8=�g�z -H!�Ʉ��XT-Sm��O-<)~j9��O��o������E�J$w&#�������*� ���9����@s���\F`�q�Z�#�D'v岖)�A�b���R��}�e��f}aQp9Z�V�7��B�F�G��R�[��ъe�^p��8�0`���)��]�x�,�(��>B2�r�3�w�;��нya~K�1��Lxz'u�B#���r�L�)�1ܔ)>��"jPA�)&��[P@)t�<+D���Ì���5�����ϒ��ʞe�(Sή�����tsI�U�������VcT��2%��4ŗ���G���=f_���N���c"tp�!B�
�<�TC��Γ�n��'h۳�e�)��X��ܿ U2�V^�W�Z40���M5��#��&�kq����r��FE��F�\� ��q�D��+���l��[��B��Y_�p��dq�F�6���_����ҋ�T�[w.��@�+'c����Fl�%�G;�]���^0��fs�e���Xq�;��}�U^�
��dr�m<��p����b��S���c3�!]th���@Ê�I�N������"{�̌g�l����8P�ϸߵ��Y�~	���>J��� �l�E$�M\��Z�D��\���344��ϔY+��k�����:KzRp��=lnvW�Ѩ_V3�X��f�Y��N!��ki�V�[��i�҆FQs��g �k���*��뗎�T%�9�M��O1���9�M$*#���H�#�e^���Ymq����k}��VF������/O7�*��^#�7�݅Y��q�����4:�ү��M��� 2,)%�)ZT�ofi@���fǙ�ZJ_Ѫ	��S�&׎��{�;��bD�2S��=�Wn�&�Cĸώ���rW�f���c!���>Y|�+ا�x؝g
�@?����
�W��wMiW�G�0�j��V-�O�-P}I<i�������IU8��j���L`��%��.�J��� q�$R����݆]'�4����\�'��s_�^êb�J�ʹ��
�ԓ+�;�Z?��.���|��Y=�)-�k����r���c��`�][v�]�I](5���=oA.`����_��n��$�h����d� aj.�h#o;:lCc�V_�0
%��[MB�����O������'�%�T�Jz�m3@�h��$�c�X�]��rB�{/CԶ�x�1���i�ò�&�����Ơ�(�?� ������d��0E�lM�q���Ƽ��9b�������Ͼ�C_Q`��C�,P���u�'��Y�+ R��!�	�4�%�C;C��~d���ʮ1L�d�Ӎxh� ���
$�B���Ae/;�,�>�P�Ưy$��w�M�5F�I�_�7�˖��X缐zp���л=�K-�MF� ������g�\�R���ds�!`TQ��E�Y��,I^��xV��i�B�ρ\&�\A�Țm6C�6�"=S�G����%�R�f�����n��[����p%�!kpB��w�%Jj�'$B����� �z�X�Р���ѓrW�-:ʣ��E�R��|�eso=�Y	�
n,;p����rAڸ�W�f&�������_��=�����Ɣ��+_�ݕK���䗩g7��t�`:��r�p��K��9,�1Vl1&HoR��-h� [�u��!�G�#ԭ��'j[�a©18f�R��������w�u�umn��0�;F�s�"�{�q�A�8�Y�Y,S�[q���Z�I�!�d�-�l<(r�0�?��-!��I&��s'y����"Q/��z2��69ظ�O��j�&Dʏ-]�B7p"ԋ?��-��٭W�c˩�����!���9��c���q�;a�?��}�xNߪ���X1�5Y�^���h*<&ۭ�h"y�
�܈��@t�g����}�k��L�
��&�a��I�!_D/�޳ �\zL-񹭜s�,�v�z��8�5�j�~��B�Lx�̰ymR<�+��[q��K�fyI��7�%T�`1�o��������T3Ɣz�*[��>O���L����ſ � �D�U����}�bJR��
^
K�ކ�S�U^	��dY.yj�꫙�D�_����N\���VT�G�Y�T����?�������z�	�������`��m���e�뼐Q�Q��:6���<5�7��d��"��v�#��F���PRf.3)o�C�`�3���p]�*K��nX��K{�����mcj�>8
�=�/e~���@��_wŝr�>�of��o���=O]R����-a�Z�w��5����7�[y͕f6)�WG_���l��ՇR��%{O�jx��!�#�h{��]3��b��{	�n�Y������(E90�����t����B]ǹ�?A��)>K�~�Co�(#�2��O92XD/�8:ܨ�}w��H�f��)3Q���oS?h�x����\������P���$���3��Z�N	b �0|-��<i(����4!�[Y�kq�DqG����W��%�#�@|���f
ZV&I#�=���r����I:��n� p�l�Ո��0�v�����	��Nt]�Rq���8���}�=�h�7��+K�G*?�@�%.���v�x�G�tW���!'�!���7��F�*�{`�%*8��*�#pY�:(�SO�
	A�U�S���莽Ű���}�ۅ0�1'�^y�]���,��V��v���(<��_w���y�:�mp�?m9����Ǆ�!RR�FB��J�(��hH�i8,�1���m�����s�Vz��l�L�u�r�����K��VyWgQ�'Z,�t�ѫ�bS��;���aߞ�KUu`�n�,t�c� j��bSH{���b$���h|}��_���Ѝ[����碉���(�.!_1g��Pe�u���봫.����R�]��>����^#�Ѐ��H��|RL�t3�:�[E.z���d��s������|_o�I�L�H�"���OB�q�g�:ݹ���"xsh��⟱~d�
�[aK5;�ꞂA��|�DZ�?cV�Rh�#��{Y!j�I�˵!ڗ�G<!�����Wl�d�{�g�7�N7�iRo� ���j�+-��ӵ��؅�Ԃ��_)\G�� u�!n�I�θn� ok7�a�Sҍ���=�K��z[F�d��|�.��[3�~:NԆn^��(;](�ض����1����Y0���ڢZJO�ȕe�Kۢ���چ���}m4A��a`�o���t`�6[D��鹄��GӼ��p��8fl �u�������������kT�'�{n/��!��&�y��D�#�m�a|�����Vઘռ�:�D6�T*���D�DKJ��a��`F��1q0�h���`��N%�C��cf� ���"�̢#�����5���3�H��2�M�� ���m�qs�6B}�G���?��Qg7 _�2�F��~���si���]s�)Z���Up��������	�*���l*�3s��.��h���sL�,C^7G�]�)8 �&�b:�-~ˋǣN��[1�9�d;�L62����;�q�i=�/��$�HK�D�������X�4\-l/�"�m6��'��WE���Hn�nR`���6��Y�JaΙh��*�Rj�㓈#��s�|C�V�;e�|����3l������G`�q��R/�(���,�q��x����Q��ư}u@�ɹw`G�&1��)�X3�_�����1�T-���E(ev��� vL�ᆨ��"�0R�ㄸ��&�Q��N��i�����.�0](���aJm��8��u�v˒���k�q�Z$�F�W����r�����Ο��xP/�������E��+�J����W��k�}"̐�%�d�����e�ִ�Uҥ�v�����B^w�9��Ɂ��C/j ���u-��]��g�����B5>M�GSXL["R��('2�\�6<u`^� xK���V�+���0\|Q�2��Y6b�� ��sy{1�&�\��l�A����D|��p.�1���m�#Ab-P�r�ڮҜ+rjA��.�p�
Q��{��W�@����G��*>�c ^�r��L8��c��m�b����'�B�����M9����`�x�L I�jF
HL1<�9�D�(����s���u2Z�vLTl�W�=���e���n�1.�(�)��;����,��Z%Jm/��NԑY���
j/�l����)�Uo�,F�8�&�]͏�?si��];B�iV	��$��dL�+
�(�����E���:�'�$TC��[��&7��w��9:�Ȕj��2%d5�s;s�'�4�ϬG�� �r1甊�0�'��j0ŉm�ǋzE�=�m�y��/dd�osVu8�#���lI���eTB!�%��/�x��y�1��A��yx��h:�7��L�<� ��rY�ō�E�j���{��e��cWf�sE�I����#�*ë;5��rAs���3��%�ڶ���Am��׸E<�,G�c͜"#ӣ}�ݸ���t��T3f���p��A�d)s�b��$�f*m���9��40�	}��ޤ]۳�w�zein��q�y�X�&�P��9E����D��y�4��{��GڶC�?JO�
u�h��\1U4c�J���of%�>�G�8��JӿGB�4~)�y��F��cVa2	D�(E֧y�p�ߠ��Y�a��#�z�%���/
U��̠��2�,�Wk�V��V��dGPӭH��.�?�Ԣ��`tG�tT�5����ϒ�\�1 �؈-�6'#-�Ðn]����ml~6)�#���}�����n���va[�ɪ�Ms��|�+��S,b��<�,]�H�u�8T)K
���D��ED�zs4�};�|�ePb4]I�kI��a����D�v���JJ��a��R���QЅ"�̗�
��Ӭw�g��}+w�2�&����Xy]��=�YW�Ol�y�,d%��+R��?���%i��;�����c|i�O�ŋ`SWn�s]��`Z��=��n�ݽԜ�km�}�����(�o�T���t�!2@$�(z��̺Ɩ ���8���#�N����0L�Kficj,e������]EjB���筟�h(C�'2��
߶����K�.���_Ʃ��O�l��~��!df��}�:˗ �^�������>e��@��c��X��2zt����Wc��f�֓��ؾ����|�[|M�I'��*�����R�����=�<��b����,{�*a����W�td�A-�jaW��ضc�N(�/����²���!�@9�X��<���
2����䑕�=����&W��*���$���	i��^���ǆ:c������I66�!Pi���"������Z6�_����F>�tq@�g�E{B�x�����dʂ	�|�ܷ�c�lHy���.v����-I�z�z��bw��;K�bUE����;�L��AE���	}1j:+L$8"�� GI�r&y�fu1�J3Q�i55*�Șrzn<�v��al2!M1.P�a�%�(9BV��x�O3z^r��{�-|�$�gnqq��zR� [Ixi��q˕���m>A��w��������ඛ��뻧��MһD��,/C���o�ʤ ���p��*��J��dt��L֣>:�IY���J�ج4�q���~�����@��Li�M���� ~"֘�������I����X���j�j,-�⾹�۾ۛ.�����yQ�l_�Q���.�e3���I��F+�|�;�ǐ1�AcQ=}L�ڌ��E ���V\�d�F�6�w)�FeF YO0ƯGn²5Yg���ľ ���$p´�����~ίgcxd���X��ƽ�=�l� $����U}"��1���$A/<e��J��R� >���G��-�\�l��}�v3lc<�i���U�<�0닪�f��C�m[w�I�"S����h��@��ƚL���Rĺ����om!�'/��Q�u�%���=T=����-����r��v�=St p:�ph�s� v��͑�{`J�L�&��vP��"��m�;Cn�9�z�ݢt��-Z���%=���!)�T��=ь/[��nC^�n��Ƭ����0��"ھځ`�	�N<B�����������;�^SRky�����;/��3	�M���٢jP��H�d���O��H��D\^����ihB�E#9�o��&��oI:ch�_D��w>7K�g�.*�Ě���u<C���h_.�G��%x�l
���f����$Ⅸl'��-NXn�>%�" �y���q�����״L�[Юv�#�=��u~|�"I;U�Tj�4���}'�Rຬ�	��<�L��mQ���W��+}Hc8 �#J��V~\��Z��բЪ�(v|�Y��~������*w�U�l�$$�+�{����I�<o�����M�Ί�U�+q&�UZ7�1��.r`f����;��~��a���]w���J�í�z��WE*i�U����<H�nY���bY�է"t�h�I�����?-E݇�Z5�W�x�����Ӂ�O.LnC�O^Φv��Ǫ'89N��{!r#ex"��A�S�}{uQ�n%���m�bn!��/��T[�v�3��s�d}A�
��⚸�pN99/���Ty�j� 9aD�6����</T�Bf(+��줿���xj)�,�I�ǝe�\���_-���8��D���a�
���-���r�����������|~e؛����f�3]���PM�'��@�D��~���#^�L5��v��_?^.��i���N��n�w(��iD�R�L��*�x6���_;��K��GaC�U��xn�Lm���T��s��tܔ~z�Bj�������w���.�Aɰ��r��p)�e����Pu��W��ׂ6�53x�6���T��f�Cl+����LK�0�^�������-֑�����}n�wȑI	N.`v.u��V&�}�#���h~�S��N��k߈�_Yo
�O��˳ �u��D���1u�q̇C�}Ӯu���?�ἅ#7ҡ����TA�B5��9��N��E�YV�G9�Wi��}H����԰��]�*����e�� �(�(aPf���y��x[y�)N�h1��I�����(B���>ަjR�p��9�C�H�$7|M݃�ͷsu���^q��`E%�����
���O�8� ��L��]�v�x�������	�:AB]?�s�)\�&���x#=��g�!��!i�i��q�S�3aS"�WV�x��D0�(�Ǜ�+�U��
��q��	ܜ�|^��,��t��jpӽ%NTOV@=1;SMVIw��O��T�g��2��C$ρ��Ҩt)'K{j��+[5<f�0��eTa��ВC�)��}��/�X�V��d	�;+;�)�lrx@:����� e9|z8Gq�K�X.^��3��I���	����|�6�����_���=n��H�aO�OJ#g<	���nt����F���^oIl>���dd§�Q1��$�pBeD�K�qav��mN]��$��^��²'_��E�;ڭ��@����]��b��p���1��R��ʰ���p�ӢtH��֖��!��
� X+�SQ�C�t'Li4�\j.��x�D�_�pdTV���0_e��ęS���}(f�j���&g�`�7�@�K�����
pT�#�p�Fn>e���& W��xWLġ@^<��-o�[x\��R<+�z+_q��Cc�?�:�m� �ʏ�?�jɏ.a��)������@��OCA�_Wx�S�/q!��C�I*�;gN}��{� ��4Զ��+�/n\�Θ��F���������|����Ɵj��|pi	�ݔNO��gG�HO���{�w�� �M��%X*D$��N4&j�u@'UkW�X]�݅�	��՛���qY�B��Nu9 czV��n�!)5�+�O'�.6X������`�v�;�������� �lDӶ�\f�3��Kڼ,vi�a.�0Jɿ�(Tl>kQ�uw\{'����l(!_����rX�\k����������	c� )��Q�b�I������.вGI#�<� >�i��4�ҤrR��>H�N��wW��z�W-+��'�Ē0�bQd��_XCzA����U_�W�I�q�5�UQ�]C��gD��^
d���dPD�� �{&����&L�M��3(��eskFx����!�S!/���,�4Չ;�C{r�2�7ibH��A�jvM*aRvс�w¦.X��ȱ#��W���\0lO���y�z�SD� w���@P�:�~V7@�d�-��p��B�}�+=6��)�B��M�}�!� .nɤC.�
Y�co\{�d��b���K�<��^�k���m�k�&u��ϩ�o|�<\�C��{�ϖ7�g-�Ύ2l��j`!pj]�m�s���T�`��Ard@t2���I�b--r�*K�i����2�f���d��v2�-�n���!]q�Z"C���������"9;���6��r�,
H[6ｾ�>�J�;_��x:�Mu�/p���
���o��n������ ������0L�K�9�@S��`�m���Kdj�S2
'B�s4���xßRZ1!N��;]u�<�ϖ>u���XY@�"x.�L[c	]�ֹ�E��+�y��*}�#��鷧�����}4U���ǽSK*&g��+
:P�8�B��[F����^J�w�!�/��	��D��.�%���!{�9�)$ȿ�v�V_Q��~�i�%"$�~�ݩ��
a��З�н'G�pb�Z�����j��.����¡�O+N��!��K�g�Qi@#+m�Y�\�d��H!&.����h������z�.��I>@�R} �����c˛�	��gt��ʾj�/_ۡc�f9�ԡ��O�M���D���0C�6����.=˯�@�n/W�1�G��oOњ�~*\-�V�M�`Pk��9N
3@���l����ϯ�P@�7���0�:�9z[��<!�B�����?�-���0h~���j$��ˠ��K���*�ٍ�h8G�h��!(�c��*Bo6Z��E��G�NM�)\�'2�&� Psk�;Cn��iB?�L��|1LKB@9�^	�0�Z�x�Ґ��>"3"®�<��ZRܙY5��Sd8��B;���W��1����6��i��x�<�CD�����]^�L{|{�3�R<�����+��^���yfH�T&K�#Kz�:
�W: JN%�����Rt�����gp��A �O��ċ������^m|�j���Ʈ��GP���%�������t#�רU�
-���E��t:`Rg�1�e��X]��*6�[� �W��M0Kp� )�K@��sk�l���%�*�%�-���^��<�b����	�J��T�`�#M<�xO��+ ��\{�T(I����VU����ő���h��4��jm3R�������<{�p�;$cOUwuZ����u��+�jZ}O'<%I
d$X�r{��z(��s�tJc���iCc��祠��";�����ՄNIb�9֛1�4X)�u�U,�S�,�ZH�Ēg=�jCځ�@qb�H��}�e%>:���X�Gو�#��1��@<~-�A��g5���z�o�1��Y�8|j}v�P6z�qG���tG�[�{���v�|IZ�/�N(�xHX]���9k���N�"�?[�,q�O�'������U6��\oE�<j6�`M�2�O����T�����>�t�8�,iha�t__{�Zs�'��	/����u��� ֯��۳@�i�q��n!�OBh���{)Kԉ�oR8@�y�����z�D7l���>��-<t����z��0��;D�⥮�L�UY=��Nӄ��P�Z�N��y�4ܼ��7H�Xμ%y���Ƕ|gO���<�<�k5�K���*jڦuvC��7���d��g6 ֎n�#�_�L��]��va��jU+����0���C��̦�G��.��*�R.%��6��kC��۾Q.�![r���<�� ���da$��X���P���6S��XrB�z!�xEq�G�iG�����{�˃y'�4�:���ąj��RXra=� A��	O) �K� w)�z�-��S���PH"��h�ɚ�Ƿ:fx�Õɴ�h�q��"�{o���D�%���߅���k@�x/�)�8�j}o�r�Z\����k��L2ϼ��Ŀ�Z9#u��e:� b
#�3oL��H�Y8�!e˼n«f��n�Rd ��dm`�D��v�iɄ����n,�39�4T^fd�6�5�Hֹ)E�$��Vi'{��̈J7��ma�]�u�B���g�ĳb@���+��ڴ��hQ �ZW�٢��y"�t�>��)1n���\ą���l�9	�Vb��w2��?�Yozp7kV?�D�_��Sb��L4;��E���@L�r3q���)�����ݐ\��P�4�ٟ�lªE/Ѥ+��2}�<�8lKk�h[���T�]�1v�ܵW`��������QmB��9 ͦ���~?��U�];����a�ƥ�ƏSg���|3k(�W�r���$Q���Lt`G���Հ�I�(�@�Y�ޙ%��O 6ǅd��&^qؚ51#�2m/�~�C�o��D �2��m6��n�� �f��b:��WE�wX�O�"K�[�>�q��:L
�JE��P��TK�Z2�N�	Ț�)�&@9�5�M�A�9��PRG)�ɋBD����g뾦$�_E<�K���u�u�-�X�b�2]��ƒl��i�ʂ[�{�8}� ��4G�s`��"my�a��4~BP8̡�W&~(��0��Ѹ�����wq&���ze,+E�aR��%����N��i!IS�>>]Ҏ3\���V^�~�y�D5AR��;F~��P9{}.���I��I|�O{�U�1s�U��o3}��<�K��J%]k���b�����8}�����t�/��iP0+}P�+s�q��~j�#y�唙���"B��#p�������(.Ԍ�j����{=f�z,�W�������|=r ��y%+�.�k��!rlw��A���ߕ�﹈�7Ӂ�v��p�I�vT�x9}l�=�l��$�&wY`�2.]��ᬕw��V�9�9����N���O�%s��&Z�}����G��9��_PFUs���	�ѽ�;G�6����j�=mhr[���Y�kF�KJ�W���-�Ь���J_ټw�|�9��N��ߵ�VE4��|9$�j�w3�(�fÌ" �T����_��� !�����Ř��{sf|���#��_ލ�2��vP5�M����D�/��a�T� rO E,�
����Z��q�k�	��me����T�@w�v�ӂ�{l-�ŉ�+�o��3�*��\��aѝH� �/�X��60��d�C��T��ϻ4i㽉 �R��2/��a�]��J��ġJ1�h�7~.��Xg������ږ�l������L�$^/�6�	�[<�mQ�6�@B{j�;1��o2J�����O�rpX��y�؈���!�C6}��A?W��h[��&�ǥK��ٽ���h(0���H�:gw5�~%ۅ0��12�x���ݥ���s3��.���wd���ݹ	
�jg7�i���q�jĂR�\��ρ�-����o�Av�pl8{�_/x��#������� �c���R��D>�$	}ʠn؛�~�2�*�}�u��X�e�b_�@�{��~��n7DH���qtX>�
�GޓX���Hҙ�[��E��%�}��I��3?��`RN-O�[��g�1.?��q�Y��lf�'G�L�PS�6-�m1�v��v�0���@��L�O�#*���)Z���%UX�&v�EÚYc�:��QCF��Q��8��B�.���J�K��N���=@F�,K"թ_X�J�ܻ$�R�#���#�~PN�����e�N��.���-�v������p<�L��u��޴y��y�W�$/��I|QF?�尔O��;�%��}\*O`-r������2WH#i)P�� �T�Vcz�浍~�K�9�9��dP^F4,"���a��Fd���gv���=z{.Ӟk�pKʧBNw%�l��ϧP��w�̔�J���)f*~�w��+��&�>JN��[��!���'��Cɳ��19lx�~�N�=7�::hӈ&�""��)f7��͸ߨ�o�b�<hR^��
!(9<�0T��,!h1���Bo_�aN�/?����\��Bo8�&��qF�d̽�uI��wQN���%�'��y���V�싕���"�HdP��,oV|�ղ�-���p�Z�L;�g*���13�JɎ�!�֓K���B��D�晈6��\�o$.�J�mVx�#e��Εr�g��t|!��<:p#���<P�T�%	�|��k�X�����@jp{0��:�0�#�h�@C)�K`���5wQX4��W\2��rtSa�6���t�b�M�l�r�u/Զ]1y������J������Z#3��K L�k0�� �1���Hm���������t�ڃ�BFd��s�_d(�B��|%<S��*r�Dy�-O�zBߔB���]��������[�Z�n�$=4D�Yq��_M�%t�ә����ڍ�N���b��l�XGJ��Ȟ��.A"��ES)���nW�٨���N~��/7�䶽T��l�y>n���?G;�!�- C�DC)�F\ s�U՞z`śy��r�ZO*-�j�Cx�9����,�WJ���eK<A�4AJ��1��h^`vZNG��n9���&f.�eY��Mh.I>�x��R�~�����mú˥q��Q`�k�{_s8E���_������:r�1ۄ#mg�i$���:�fÎ\.�wK�����*q��
�6���IB����̂�
8��ŝ0�����o���;��w�~¸
��P��Sܳ?��P�J��Q�u{�ۮ����۶�J�5���3p7�E�Py�o�� f���g�t��Q��L�1��t�MV��i3����u����zؤ,ej�ws (u�O�����阍�mn;8���f��)���h��J����`K؇������a�h(;j�q�P\Ü��q��L|xGP"LF�k�rD>�=��.?z%P?�o=I̕N@Ŋk��XKx�sgg�jE�_Wb.�Pp佮LY&������3�_>a�Q��c�A�o!K!�К�i�q��*1}H�jX�Z����[�;4�o���yݳ�
�(gMkds��ϑ"��]���u�P;�**�Ls�&4�O��$���',�B��2�U"x�	=a��?�EzL)
1M�]�
AT�/(���<\�1�;�r-=��+�d�\M\�l���VT%�Ɛ���*�b�l�~*�)#ih���K��g��������u�OAK/����C������9��  a��Ӛ�J!<l���n�4PޔkE�j H��>��F�N����=���o�c�]�e|ev���1U�$>��[�3Ŝ�ZWb���9(ҡ󰡿��s�Ǉt�˭W��E>&��)x�r�ŏOB����l�,I���4�`�>9]�$5?�)��^hu�x�a�%���Kl�}�<�D_? ���؉mDe�e뉎o���Ҕ��f�/�{��*C�q��	�9��	)��iS��E��y�B�7xZE�� `��_KwF��1dY2G��C
���n*�)Ē�V�m'��2�nx���#ge��f0���i@��t�J*�Z�?!��`m�9۾� �ܡtƧ�t�n��4���u�8���l��i7J�ԉv��
t�R��{n���$VW�c8N:��9��c&�F��ś��\���7�}�*�	��`���G\G�/iǓ���,xl��_j��� ՋF�Ee�M�4V�;��l�'�C���<���BhYSQ�߬�HBRzB�!EZ?t��tVDN���@��'���M"m����]�Sd��{V����n����6��`�����iR� ���>05F�n~���a����κ8a�*Z�UYt��vPa�b��2%R�C.wX��*��$�M1�0�f{pF3��<Uh�]t���C���2oXC���w���vT�Inx��L��1v���ѧ�����]����ύr�g۶4�]K�"���P�(iKd>(����,j��MqT9<$�� ���+��Dj����� �;s���/>r������,Cnc�QM����.�-N5Y�<���[u������`��L�8�*��:��_ɘ��Ct�e��\@�2�f�19&���U��-I���}�����6�l�\h���u���$w�(8/�	B-��S�,����G�/��w�����ɊЩ�p�͆��j��G�{ �ޝ������ͷ�u����MiƏ���H#��a@Q\a;1�j����߭s'=�$�qUVW���WC��"���i��w�� Y�!r�O@��$WSj23NÁ8��+W��l�n�H�C(!+��b0~�O;k+�Za�)��L��1�������&��s�nHVE$|n�'�& �?oh�vW�&�y�k�v�+�D=�j�9%c%�#p�>`T���`�Tir	�c�/�mxl�jl7גj�b���{�l�7�෸���_��☀���h[h�&�Y��+�V����^�J<���2bo�&]Eۘ��s��9�gdq��c�~��������#_��bg�\V:�*��޲��Y
$�rEZ��;z������!��U�LP)#��ȣFE��K��i�,q�N�YEt��ɲ#�&bì`l^}��Gx�-[B�2.~�ʭg{(���TCx��L�pֵ�t�?���C�����H�8�U6����dS��I�R�E(LsG��y�K�B�l1��a{��75=X���'�)�J��`\�ȍH�tM=�q습}q0��J��U�������ߧ�����KC9X�C�Jͤ�;P�P��Z������!�#��(y5[�/�3���W՛S|d;���
�����u�o��1�$a���`C���q��
�PRV1]Bnu<Tg�����J�� �C�ħ�ڤ1�%�p�Ɍ�lԾ����f�0o_0#�t�}?̍|B��Ә��	DA�����G��� ��x=�n<�b��26�O��7;)y���J�E�5n�Ě0�L-�^;3xc�U(Dv����4��� �
o��g8.l*��S���r�C�'b �/����:U��ǯ��L�>�fKJ�Q� py�CRg3�y@@	T��'�4��q���J]Ü(Y��.���pa���5v�m8�kT���#������򱗵Ž_?�� ����61�:��I�FM�i�{S�5o��q1����ㆨ���s�d�p����$�"fd��,�Y�yf��[����~��.V�]q�NT r=�
��V.�+
S��<L�KB]ȒM�xZ���c���µ��Wve�xʓ����N�Y����o�%Hχ���������h�_u�_1����^�'P�WG%<rh�@舙ҏ�+�reoQj�fX�so_�.X4*�a3!���"�&",���!�5h'�?��Ci�<�Np�W��n�7Or��!��tG��֤���|��
���@@�g5Ic�	u������6i�9�s9�w}`�DF��Me>9�9�Vx7�{���R�{��>���!o�(ı��m>� y�:oG��к����}� U�Gn���<��[>���e�0=��O�,Cζ�:��ǰB��U/�pd�$�Y%���-�R���B�лh��"�������^-QZ�ox�13�@�2D%�M�����+p͇Hy��h���Ԡ0��[��h�t ���$���{��#�RB�������ʹ|�E\s�G�Y�k�aA�E�˱�;ħ��ŏ g(�V���S�઻E���rS�#9���^E1lO�n����!V���Xt�ٔ>��֋���g�Kw"!���2�<1�J�����46ѥ�4�$��;Si�S��'��L��X��8vsn�f�}�Ѿ��(<#֝�w~ݧ{��ʅ��,39��j�)�:A�F*�Q����l ��!v�g��R����Ww����?@�Wk}�.tM�(9"��3�L�j��I�3G�U��z���%�)ܩW�Ж�|����}�-b�v��C4�_{X_�P3D�[e	���>����]��g�o���5L��sq�=�/]��$ރU����Ep~�B�kԋۅN��	l�AX\ˤs.�C'Ѝ~�?#�T�}���F�e��@cc*X�8��w"��3�TUI+-�>%:�fIٲ�Kj�o�e
֕^$m���9]��'�R��>l=�
�M͒��}�D3�p�>/ZZ ��U�o�Y��B�b��Zw_FD�M¥�(B��$���j"B}�oW��� ����Ht�)����r.aH��r��}Pkԯ)_Q�$M��P%�Al�4C�8U{��A���(������?\��V0��s���~V� z3Ǐ�����̐�у,̾�!L'��u���*�9Nx2�T~#�P��ۗƳ�*C� ��bӽ̇aw��J>,����T��*�?$#�O���L�3�Q~��25�ǉ	Y;vW9k:y:�������-D�Τ4dL�Al]{#���/��S|���֨J�0��D��9R��x.���:R�꣐>ƣR�噵�S��0���HTH��0?��5<r��`�����/�d�p<7�����|$ߺ�r�,t�.ٽ���M������1ˉi���\yMP��y��ח�E.ȶ�-!�q�H�o�0����
�`�D6��'�;C������z/�Iy��.��* k����-���+�e��R�j�*�$�lWr�MC�I;Q���XU:�V<���r�Y�OT�����������N$#gqS�@c3��ȓul�ᱫͷ�($�^�-5��o�����XuU������]�����Z�WzN �xH���Q��/C
cU���MlW��<)��%݌X�7Ԝ���Lsł��}��;U_�fn�62Z��K���G�qw(����;��6Q/U��z���z�q��i��S1����K�ɅE����g���#ve�l۔.+p�t���T{��������������E�HL�C�tF��^Z:��G��n��K��p��n�pqX�IbU8![�agۓ���׋QD{LN6'�����R.��NAKM!�qSF�83�}%#��%|q�)�q��e��Ț�`���6�p��F�Z��_j�uy�'�3�P�Y�L�9���k�wp)����ON�~��Êp�AEu"��L=�NB	�1T5�``�������Ng����K��K�#E��2��ձ7_�.�(q�
�Q�n�u����=a$q8Ұ߱�YA��]��%`6�3Z��@��Z��n�/��V&a|n���tm��b_�1o�pc_��u�5
*���)n ��J�oeB��TJ/11H�Z9��A����LZuā���$�v��]���FH��!�44�����+%�:q%i�hW�4������qo��`��K%ͬ�&�3���B�2�gn+�c��"G�D��.�X!��#�����;U�-�Q�W�؀�`�Y HZ �-m�A�g<�m4�ʽ3���N"�8߾��;�mz��A}�1���~��3�H�إ��/���-e�0,�$~_�agy�s[N�"f���2ӳn����1Q F���$������snU1�����S/T=�K,6�ئm��u�ș�mԝ��2=��t����-�����'#��Ajy�����^r��܈M�2[�(��t��(=�^��� f����>��}Ds�߭ʡ9\F�U�M���G6Db����ƚұ����^��1�Vw:	Q�vȔk@����9��)��84?�FJBՊi1���x�rT����F3����T%���Pj��L������{#r���:�R�r@^鰧 �vT�[�m�4�|��K���B܁���[���*�92E"�b$s7��P�#��J��K;n���؀"r�ʩ�g>'��a;ߵ�D��������FW��[3{�jղ7�[mǀ)�?�jd��Y���o����Q��{�,Z���l-�9��ˉ�:�^�K�����X�D���l�P��u�M.����s�r��K��$T�l�H�u<R�hp���J#��=s����ZV��O�2i<�C4�Z&(nM�K}�x���m���y���N����P��	�I�L��c$Lذ���¦6"~XPW��;p�$�^I[�#�PJ��k��XHހ�/3)#�ؗ0A��}�G�ح�(��s���ɫsw\'�A��!&}1a�;&54l����p��+A2;70�:4��O人�A����%,Gl��lXY����M����+0W~U{�!`�H@ט�ȕ׏޷��S���r��6gZE�ܚ�5v���R����זV+@$𒛤x"،��~��_<Gy�j��F��r�e��s+�c�g)�i�8��3.VЇIT0�QT����.i�Y���:H�5�zJ^֐�Oǉ�NivG[�ö�c�5A�Ս�c�.�-)D��ўSȜ1�9�S���$��u�9��7��
��u���'��`kT�q����;�Piy��-�_�6�����Q�o�i�p�MG��M����b�+�%�S�!|�qg��"F�Z6v���S_,3`�3��^��I߹��S���������½��?��H��� B�]Q�DnyNBG_1��������:]���@���Z�O"��c6��� M�Ӗ�@�0$5���@I�H����û�]���)�v�����F6�]o����~3�<:ۈ�({P7;JS��δ�W{%Jn�@��!vldyt�F�愭���9:��N]E�vO�غ1ґ�sc>sCK q���r�n�zq"x��t���y��`m�����.y�r���c̯��4'�S
6�vy_��3�U���Ӻt����D�F�l�~ܶI-F��Ć}�[����Z؍m�����
� �R�ޑm2��D!�_oJ���J-_���.�x��3 �\���n�{س`��f~��U���=GP�{e���|�&�%�����	.H �{���j�A�ا�Ě��<Y�P���+��IY"Z6k����Ա%gd�-��a���wt�s(`}��4?Wԇ<W���>ZMC�F}�QC( �O��顣֍*T:y�"f���u�O)�pSzL����EVf>�˶�}��_�
jCF��n��6B����^$l�Y��@⥋����? v�z�QukC��ܫ��u[4�SK�������{4?E���	$�#��%v��1�d�%S\�J�\��5=�Zм!��ru���ʉ
��=XK��m�1R��+X�ђ��I�M���s��1����&����ė��p���q�8�M~�;�ꡨ�t�`�T��0�����������MK�Xq	1�ݻ�Z[J!�� g]�xsdD��1-�NY���jq�~�ZC�.� ]e��~6/>��xO'�M�uqa&B�/V�d5{+G"�J_��Wr29��k�IO�t�_~��a��9_�L�
��}��j$��̯�u�Ii'?�3]v�bӗ���yE�=z���4�L�:�w�`Au6>0�l��v%�D)s��E�^O�R�@0�P�fc#KQ_�u�d1��g֚Ӯ8���s����:yjE��P�:��>}��⃑~aXጀ��̙$����k͇�_�qp<�nuV,2}B��W���F*��VC]����Z�Lw�i�Z�k���* �)ϙi'��l��C�U�(������X@�g�y�=w�QR��9X��	�ۏ���2+�e	M)�[�׈@�H����[����EV�рii�����c�$֒�vs������k�����5�Ptt������#	�S[u���U\5�~Fv3V}�Ba��Zd�1t�I�6u }�r�w�B�F}��e��	���.d��t
Z������HF����\�2U��
�*�XQ�I��ޅ����k	J���$A]Ӝ��G�ƳK�@P�� ed��#��9��B�s�`_�Edt#�%m�➓��W.�/A���=ݑ��܈LrI��wq��ȉz �?��-'��(�_�_ʒy����m�r��G$�ߴ��w����oqZ$��D;�{�y����~ �o����Ab�U�HI�C��@�/�oQ�3�֭���&�A��y�[V �D��
�7�o��$�����_�{�b~PWx���Z;j�²��M��C>��"C8	쑇�_�/)��C*c�{��Z��f"<��0[3�7����{(A�(�!�ѷi�%3;fz��K{U!�B��w�����1�A�L��9�0�T"$�/ˢ;�/\}�;�L���L
>?��~�s�dL;�� ��-ZG�[ݷM4JGS�=߻z^�\�����
A�]�Y� lT=#/����;�p�	�m'��[W�`�̉�-��zM^q� ��m�~�����n>rb�ږ����7!}�|Љ�&�>y��6�K��E��Y��(f��DLw���:"�`����c~��o�w֦rɃ�P`b��)3t������st�'n3�9�2g^f˖��fM�}�BD��g��M�Cx3��n�aE��@c�Ұ��Jt� ��8z�ALW'S���#��Χ�Ұ�~���'��.:gZ]�IZiW�g�ke[����MhAc9�3K�Aj��b�mc�����.h� ��x?_��f)�M��M1�݂u���%"�;*i�e��'�!h;�eB*��f�[��v~��ݯK��}�Ѯv�L��_��t��:�4��n;\��@�x"{��ut����Fo�c�]����t�%Ae�,���6Oɝ�|����*�f���J���;y NӐ�O�E�B���&�f�����D(�̙{l�8`OӼ�ΫN�S��.֢�n�T�7B��s7�L2qy@��S�5� %�*�05VN>��i�J%o[��N� ja��K�0�{�-��u�G�B�FP���a��i��m���lա����}�'G���%g���5d��b��奺���ٚ�z�|�����ڵ����N�9zfW|����$�4��;��F��˲�|Y!��q��S��N�w.��Q{�H��k�� y��';�5 �
��6�A%?ׇ�HQ�_��p���H��Ĥ<Y0���K�wa�vd�閻LM�>u��{�*���4�;��s6�0%���3�G8�F���� E�{��xCL-��i5�fi�8�gO�j��R<��-s�Ȗ	��R�`h��j������B�]x@
��hC2M�6�j*;�̓�v�~�́!2������S��P�;���zd��7YL� �i%�W5>�
l����+�w����_���#���!c��`�mK7�X;[�d�}JK�8"�8[�2@�6�f�^������/�Z�ݖ䶎�4��h"���Y^�M��e�A�ގ94v��#_X>Yv���R�*����e��SB�W҈I��J�����ү���U��8�#�" �>c�_�?
m���ZX����?`u���ݩ�-* ����wU���ݨ@���L6���1����:m�f����褆j�1l��S��t��5`�|�z�>�s�2+�j̷��&aT�C)��h��n]���B=�vǻ��V&H(O�}�9K:��$۪�5"�4jRd~
��ߥ�ElH)��W�%�q��H=� 4�pnsxA�8,}o';���<ff՗*�P�3��.�"=R�_k1p@]Ӿ��h�tc*p�9�@tޣ�շ��*q��!5��Nߣ�&a�Uݝ.`���]9�O|T��,��:烧�.�lvF~r��g�:��FIG<��1$'�:�+s���l��-I�w�u�f;��ӷ��nR������z@������>�C�?3Slɳ�uh��t˄��&�{�sXc�IfLkVm^v��=�<2��~
�̦��ۃP�������^���buw�I㹥�V�N��V@���E�ι���5��U�	 � ~Bv�3�L�Ѽ�ʁ��m+#t����ff��Y���M�2xG��Y.I1����U.�]b�F�Rj-�
�'���
�=:� M�h'A����ۑ���i�莾�w�k����-KdD���*C.����u�$-���$p�T�
�4��u�yp�˻|�b<�lD7ʚ^F:a� �U?�n:�sK�������oE"�`���Zs�7�;HN�?�_|0 {�U?t�^���ġ����./�����?���!����Ɓ�}:�~.|5����i�
�Ծ�K��_B�>.�7~U����t�@@�ZD���{�.v��A�$ds\鮻���v_�4݃v��]jy���d�g^��N7��j��o��5�����TOG��U'���L���E���ÏVb��3�ܞ]K��\������"%'���+"EdY����C><<1ć}Z?8���S��4\����oi�1vt����?~ˢ�EC�K��ao�?e�p�|њ���'L��l�d��L��M�m�Q[xܟ��#.`�
J�$ym~��fN �)�Έ������nC�bV+K��t8z�q�N�ƖJ�1�C&�XĜbގ!�݇���:�
�q7��0!I;S嚋'���$�6Śa�}Я�y"/�2�/��~˗�@D�lՐ��]��*�Yp?���N"}ſ�Ꞓ�F�D��wf��K�㤯�����I¦�4�3u	�$�B⌲�f��Ӄx�)��s�I�*.��)}&��p�w�Z�F6%]�v#��(��S�	R�h���IF!��]�W��./v���?���4Lz㱕%첐�]�a�)�[��&>h)Mu\\%�F:�����W��ɓ�ѝ���8�iV��	�͚F�~kI���C��@E���{�t���iNh��D�ru��[[0(,��`%y�Ɔ�����I��#�S���5��Vbz�5c��ڃ�ޏ�č�EX��E�Udi)��?�llTOz��l�9���`��ڢ3&$����vjFRL2�rr2�D��Ò��-|)^�h/��fH�N������F�zy���`�B��z˼d���6� 	\Q61�]ɝa�\��l���>�qO�5������H#��w&z�[��)��,x���k~�i�V���Α[,3k!�j7½��G�oGg$v*H�0IT6F鼽qH�bnýa�e�M�U�!��Mc6��d�fp�{I�64tG�C�*�S����;�w�6�WL8OP�_�6%:
�C]�4��b���Qdm��\	��b�U��r,V��qy��G�3�k\�GA�n:����?j!lm�����K{�B��nEx�I(�H�9�al|,��=��[���8���Ō�Hn#4m����?��D��Vg�T�d��{�dȗx{�.�vvn��  ��ӹ�]�ih�;g�oDLRı�F�E���Z_���A0���C؁.�~B�P�y%T�2��Sj�U�A{�ˏ������v$�#��ɾ��+�1z�C���lD�_;�J���g�v�*-ѝ;Q���eak����&o�4T"l��K���ږ;�kΰ���L�-_h5.�I8ޏU7�ŉ~��0_Y��1H��{���/t���x��zJܙ䊫��W�XQ6��r)�e
��)�#[h2�!�Z�:�x���>�{L{͇��Ň.���{*gz�[�YpO�6zA�i(Zb�z��CP0��W�uV߲<�V&�[*��ǹ+sa>l��
3+�%K��'�����i�f���$X\��-�fb5�ҩR����Z�Ja�������$~��jJ_oT@�I� zL��Z���-ݰ�=+�+���@\��?P|8�/��? �sj��I�2���3\��[�]��y�z$J�w�0�^��9���ͅ��A�
���(�͗��t��MM� �2�����#�{�;db��_b���l'��������YQu_% pd�22N��/��q�)Q	,���W|��M���[S��k3���[c'�!sg(=g�%�U��Y��(��<��`�?vNB"�aD�$�y>�F�>�����r�v�C��]3���6"��n�e�K�5�u6Vj[���7�)�T@�l�(�_�\e$�C�Ƚ��ޤ�7�[I��ڒ � 9���\����2r���l�%�F�ࣃ>�۔�N��x�B���IM͐7�+m��\��+mS�~\��A6�J\�#�{R�W���jLN��
�F�o+ue=eE�h	T)g��B�-3SH��I��j�W\=����ݧ.�_�����������
|�+�u?��oF����,c���=���U��?N�X~��P���"[ Pn� �9�}I���WBȼzG�"�|�/iN������ϒNC�Ѿw���>�~5@�]ܯQ33Y�jw�K����L����p�� �Up`����o�(�5n(�y��,��P.,��'����i�4!9N�m�5�u�}� ����R�(�~-MI�o%�B%c��]\��O��ڲu2�����7�<R�yu�TǑ�w��#����h��f�^�OF�f�dl+�<�:���%�0�nX����g7�:��M���*T��_��3�}���z׆�~:��R�����,{ʖ�ͪ.�����E�)�� �?�3_Nȇ��!"��[�}�6<��L\���63���k��~0���.�F� �iS=��ӯĘ�*~��4���f�uȸ'�|�o�pd�P耈|��ف}��;�z�]����6m�"�����;���hR���)Z³H�*Ũ��*���lڊ=DW(["�)D�)rp!ݱw�C�-���\8.t�b	�ftx�i�0l����f�����g
C�/i����b�/�}9��'�/:���[C8���Ҵ�H�0ś�ς1�0��=fD���Rvr0���lLݏe/#S��4����J��8��ėDl�� ^������06�3�����s�/�&��RuE![�ۇ��@l��w��	��1N��2�{s��e��i�4���t�{��&Hv/<�7�>���s�s���*^0�u������(#8h��d2�͝��M�w7��/��Y�B���<�;���0ս�I������S�q`�٭ʪ�֢,�����L�<YD�F�*�c�a 0��1� ���IO�ő� ���ӕ/���`����:�L�Ә�	6��u���� :EQ�1M+4�$��W��p���Be�< �x	�\��;��ۇ4�����#�Hz� ��~�c�9��Ay(�U`��-��Ka��&�Ζ�OP�R�G��~d^H���Vd�:�j�u �O򂡐J`n���zT,W�W.��a�ZUk�CY�C۽'ߐX�a�%�F��ke�;3�1�o@OA�/��\]4�1(�� J&�_gD��PE3L�o=P� �~H����V��:b-1~k~�8�c��P�����W%����(���+R��rg)�'Ii��p����O��:��5x����x���jO���~�A�Uˏx���WB����S�z��3,���lk�P=�Qx)'+��Գo�l��	��~�j"��P��TCxox%����NV�|=	���?�:F�u���#Wm��!�T�Ꚓ;ߟ�N�T���"9�'������x��e�4��%<20�l)���G)�x�6���.H]�v����m����Y�$3��Z�8m��O�۷��	���RE��"JA\���/iA�V;����T&�#Lh\-��B��u�e~���ɳK����K�Qܙz��?�D�d�[�V��6qs;�����0����<Qms��u	��W���f�������� ��"�f�N�{�X!����%J
#mxޯ"~�������Fֽ���[�3|� vY����6fAm��>5��R�#�N�C�3zP���3݉6�H|a(���41-p޿'h�2hh�*A� ��$�G�.3����d��`�%+$�&DA*&k�!>�!W~t{��4��*,)����6tz�Ɋ*�?�=�ly�]ӧ͌yZd(4���Q�3!��̨g��^�P�/�(a `$�^��'�0[�<�oF��n�`�E�R3��,aאx������3�`A]²o̖���	F��\�Ӕ��-��;n���(i�8a>��ܶ�P�d^ԁ?��nk�[�C����e8�� m0c���'
��{�u�r/��)A[�K��g�$�C4z��t��=m���4����̵�i4Й����(��<�f� ٗ��9����ܶ'4���`��=�hzd�v �1�w�+�1�x³��¨�.�0���p��ej؟��԰}�W��H�0Mr��_�N��F����7��"�ڡ���]K��A~�P͘�ݽ�u��������g�<J�)������wM|�2�B�L�uoF�p_	�q��J2��H���q2g;�ѻ���N�7^©�mRԐ��ѽF��73G���7�y3S�e�3�?vsN]���js9h��QV��8�?�Е���I���u��6���l0����zv�U�����%B�.��Xu���7��av�B��i��L��9���/Kx�qa�����XV�ƃ��sT��<GYm)"'dmh;tȭ�>_PnEv}d \��;�}'% P��2-@��~y�CCV�=hi�������G9X��/��UE��@��f�~����kNVN�m��,�^VJ){���`�=��E�V�n���	�z�V[�%� _f�B�)_k��$������_:�f�)�B#@�7X���4�j,E�4l���ֲ^r��p����|�3�#'�#�ӆ����q1�}��5I\�����Ucu���(5��:7����w��>%�8Ȟ����T��A�I=7Z���e}X��!�[�z#b�|"x����H��>q�mK�%�|�ȹ�RH+��5�57�b���;�lk��n=�
��L���\^�#�{@V{�=��!�Ȧ����R����nծ���4���'�8��t�,U)�\�n�����{ѭ+Z�gԭv�����Q�q1&w�G}����S�M,�L�n��š}
M���yʝ��
�m:�MI�a�Έ���0��z�?�Uϳ��h ����r�Vu�uߑ��ͯ��À.��t1s��yz2�G�w�fR��y[�N?)���� ���G������i�7Ȟ�9Qu�@��}��w��������Xt��U}AÈ��ݽ�ʶ�|mǻYbo;��M�p�
���d�u�� ��th�y;�B�{+�f�i����q���_��u%��o]�1iܰ.�{Dg�=����%um�S�0+t��A����.m����Ԗ~�ٖ�3B��	n�Y��pq4��94��&��c	�^�GK~R�W�Q0�&>B��rĔP����M
�~��)��\��Պɘ�KSh�:��y>�gݫ��3���5A���c��;o&�cs�n��V�=/���ǋJ��}7�>�^6)�B���[��Z��KI8���ڳE"W���N�ܝ����(��ag���o[����� ���QT�UO
:�w��[Hx��1o*|�aR{Z(w��H�#��Ȭ�k(�����gވ:�-S��=C 
�F���ͦ�Ȝ�Q4-�ҞÁ¼h�	
��eq�5��S�ׂ)�q?}���N8ZN�S�:�`܌���G�t���o���f[h���_��Y�֞�eg�O3��2�Z�|�T���Q7�f 9ϵ�*k�C�1, �b�0��Q��צ�u�mLJ~�ۂ�ܸf:�}v�I {���&X�̯J�%�81���3��6�[U�5\�no}���\�biw��1��Vq)<�"cT!r�k�Zb`�>�\��f��q�y�e�P�N!q���̼Z�Y ���fBܛ<�>h���j?��FP�ǖI��N�����I.�������N��T��<�ѡY$��Ԩ���8�2���� %���q�D��z{��p�A�B�����Q�	�	Zc->�;���[��W��?��,�N*��u|�]�h��q�q�QЍ�b%J�Z���
��y�v�#@wF������DV�ڡI��N��M��х���� 
�CV�*2��}���'��A$ر]�i,�-G�?�_
rK���!�CjR����%��*BTZt�y�|���k�i0Z�ײ��;�9I>@��1iB�>�Vg�jOf��(*�y�e*X��nyOZ����LU�/R%}�IgZ<���h;�,����;�TC#�#�#�o�����C�K�y���D?1�����-lr�E_����ץ����sx��U����{d�"tsv�"'����u�__��g*ll���fjqZ�Ex�F��+�$�v��M.�����N��xs��*�; v�s�8����_���RO�@t��ɩ����3wJ%n=���*�!gl�X���a��0�3⹗S��m��x��`!�_K�ŷ¢v4y�����yT���`qh�h\rY�S�G����,�uH�+�O��"uf���W�yk�_=���v�F�PUǅ1v	ͫ��~ؕ>�J�n��%	�A���$����ό�6
@����Ԉ�p�M<�IXTz���2p[�iq|l{��5�@E��4�ĕ�_T���{��� �8�,ZS���Z)�(�ƾH�Q횰�h�,���v�nU����j1����|������(���+!�Fϟ��ɗ���m!C3��n3pX�Kh���0@� n�&d��Ch"�v��Xl�6H5oͱCM�:}#:�`��Nё��6��~�]e0#�'Gz��?�a�(m[���l�1y�GA!�1����8ܺ�{�&yQdt� �#���7�,�s��k��}��:?�W�1aWH�$y�ƧQA$����W��i�"���D�*���E�Ȓ���Ŝ�����hwu�`�7�uA&���9���Y�f�^�D�[fc�h��fE�R]:8|P�m<��m|"^!u�/��U#Y>��,'�t�I`V����e�l���vw���.�~��c����������p�.�"*��\�	Yh�Y�W��hͲr�}H-t���C��ϛ[�Ï(A��W��4�b @@hzt�d��f%v$�[���iz�q�Z[w��{�G�B�����wS���:xG�{��+)"��:۴@/����#�m�36���<em����">H�����}سC�<k���藍d^�]�kÛKwl�/�\�p�v�7PsҺiݙ�@��(��9׌�>�����܆�h:%ӉY)��o)󺽶���:c�R}n���/OӪ''�@
��$|�!1N�l�]�
5���sj�ٌ�;��<�Tbcc�w��O�����h-ɉ�5�0��:e\�k�s��@:�H\hJlL�'��y�3��j��~�!:}S��,�4�J�u,�B6��!��v�2	/��^�D/i_a_kH����z6@��VT[F�AH��^�P�W`:��o%����������!2�BU���@3�i�����ז[طu��(�`]UO�$��1��V�5���D�ʅqWk5qZ/_�G�f[7$Fs�ƊGY�Dx��`��(��7%��2R%����x�H�SF�!�WP�:���yc��~�?ڡV�&l��WZ���7,���{��A��9��l�UE�7��_d���4,�������e�޲�Gd�9&)�8�1���C�؊2R�}�i�N@˗��`�N	5��⊵~�����9�4<�!d���d���ʏ�VL5I:\;{`�<�`����1F��B�b~��.��6��@�P�m��3A��� ���mf��)��y�LNJJ�ڱ�a��B<��v�埯�w��^�֦X�z��&�z����N���z�{�kF�NِM#�lo*#1mPP?#ڝl&�k��O^ѿ��l���;1o�Vb��^��U:�픔��5K��`|hx����@��C��gbbizv�D�8Ꚅ��a�{�+���� 2VFggajZ5��n��P��ݦ�:8��#�f���:���.Ϛ�a���`6o�1cKP�����6tM]�s3�&NE����>�� -9���{�(��2�m�LG�[zx���ɍ`i�ʀ�uid�������$�mK�K�����v���o�<m�g���y�a�@s	��vuer�b�O#t��n�� ���Pe��l���k���ۻ�3'�+���V�R�����g(����`OM�Mr3�����Y�g.��R$o^K��qwL�	f7ŭ�#K	��t*1=��3��.�K�^]�������Y ��ߏx�� 3�NF:�L�Eg~r&վ�6Y_�vM�-�{�����P�Z��f�ǰ���Y�hpx#����Umo7�eg$��O���4Y��D��5�����T,$�Lm������fbU����)/#x�Q.� �$ �\ To��S�o����������Dj�l��YZ5�#�V'�O�vR�ǆ�\肶(�o������Y_ٹ����� ��� k������[�ȒkfО�a���bxr��n�pg����%��㏬$�p���ח�N!�LhK��m/���?��d��=S4[�p�4M4)$����nh0z�/|GP��[(W]�j�X�MgW0칭-M�{��,��c�+��A� ���SD&��>i�h����5��bU�q��d���� Q�`���c]|�(7�,�l�����dPS��U��϶�Ʌ�Rي�lW(���]H��.<������fa���3"t�ޢ�k����9R��s�V���6]�n|��~��-��Va�S�;�(��[$r�� �ޗK�-|N�qc�f1F�^��;��f�t���;��>R/�cD��GzT���J`��5H9<�w��mmW�&Z�\J#��;�6��6X7[�l���FR񣼠�%��H.T���6��I����m�����ju� �.��;b`���P o�����\�B�V�"Ա���9��nf�ZL�ES�"Y&��eF��r�l�u����R����j�,��%��a7_�����t���V�D �	��0%������~F@!F���"�7�<,���v�a�zw��aMu�
��Ւ���񕵓r_c��ϷC���gI�Iy\H[���Ǔ�� 'Y��&D�>Q�������OnH菉���-��[����		�o����,�#��� r��`�:뺭$[)�B"b)�|�y8*��4t����Jj 7�ʧ�#����ǹ���*�<�d���fjͳb48�����*�i���ָ:�=듶�D��s"AڋkP��&h�'�M�f:��`��M6�����n�aW�:*Z�.�Q�#)[�!��c���F��1��/���ؑ\%VM���nQ(��g�_��-`��w+�r�����O�����>J_�ܞ�+|�G�[�|K��^2g��F�#��hj��S'K	n=�4�)"�<���l����_��p�՟{��ZR�O���]jo�8�NvA�\��ڥ샳F�l�զ���lNf%w{>V��髆�
���}�n�U)��Kr���|e��m�PL��<X]TO���ͪ��8�-����`�6N!gw�.(Ҹ�lO!z	�^���O�1{lDꦙq�R�]�@E��0�*i�e�ũ����"f�ۜ�,�HM%�$���e�jcz�g�xT`^��!�C�Ъ.�Bx�^��7�l`h4`&�4u��"^ C�t��*j+6E��gK2�F2�<�)JDO��#��b�<���47�Z�y%�����>lDbS��F�y<)��{_a�X�5~�I9�S��qo;4c{���尃2��+��p�:fɳ8k �����Y��Q��"�nBDo��7i�Z��w���ԣښ��N��Gq5"ds���ƥO2��bG�S��G�~ℓ8�&N��:힍]�>�'�4?����:hʸ�E�������:g<����-_��SgE/=�����I�7ު���_�AF�8�ҩ��m�۾�\N��~��w׼t!)���۠Dl[FU$C=7(��$�I��&����zX�`|?T%_<{�Z���$o{�J���H�&�!�="��*ꆷ_&�%����`4Ҏ94���㛙�[*(�\�\�ag(��H@X��r��C���:]�U�I�������=a�b���� ?��Ep��5PԅW�s�H~1�ʬ�6�d�aU�^��+,dE��=6�-S��b=n��X�tS`�Ϥ�{X=aΒ��g�q�H�,�2���к���SG�i�F��]��/���h��[k��˛�wj}gl��}�^���s�B.�_�=C�ua���cmM�x���P�'p�~q����X{�[O�Fs�'�  �d���3��d���o��*%�c\�
�������ɊiBĪ1x.h�!x���Pa�~��I�Ujfm�).=+V���� �ԙ&�˅������$3/X��n�4�%NZd��� I�Bހ�)��⤊@cbU@ϖ�Y��6�Z��K�K���̌���\cXM�i�V��k�;3̀�}�-�9�>x�7�V-�c����b{�nڧn��K5� �!ֺO^~R��e��T�M F�N��"2G��J��`\G����"ڻ�3?�Fy�{��W2@:�FUj�ʡ�E��V����z���|�S���8��5��en�0o�fuU��kN
z���9�\��J��n�>�<�$F�<���⬢c07�W�B�X}$�}ؚ���i��`���C�� ɒ��4�t�E7"�d�B�͠밬��X�4���� �ܫIp���">'���M���Z��p�����͎��L"?�Y�n���c��?+�3���ݚr\ӿ띚��Z���O����_��JpAHݸa[aޒ��y<%fn�_	���јרty��[�U$��tw5q{���{,� ��ySւj�4Ux|=��Z~�r��U�I�8J����c|��0�� �8˝|֍Tj+I!`sΖjK%W��l�a�Ս�M 3V_W�荕�`���",d�s��#7-�0����5C�'063�#�^\��K����k�"�)n�$�����WK��XB��~�1��Qc V4���	�PZ�"�T���F��@Ro�a�^Zt�S�xPҪ�Cx~(��^`���s!�^��%�ɾ�z�rR�As���T�oɝ2&`<6&�֟-(0������N�����z�c��Y���X�������Ĵ��1�6臶�%�F�̼�<~�����gv�*u������z�����A���8�����6=��mc�yO���f��Y\]Q�ub�A.*g�k����%;�̍���K�F�����q}�	|�S��g�S4��G����:Ӈ@x��qW)�~o���MN�A.�v�N:ؼ��3�ٗ�P�����}�nPS2�5&nJm"&Q��@���2���c�g�3�{�M�x��53ܗ{�Pu�-+>��Ͽ2H��4 �Qs x#"�E����?��Y������a
[טY,�\(��؏]I�2n���wH�O�����N���f�.�OXk�(���N�J�����I�mE��Q���f�ϖ\����0w�K1]��	���,G#D�!��[��ٍ߫�U����@J�E�� �U'��N�T�}J���tգ��&��3���l
�>��fc��|��Xw���#�i�5�G�� ��Q2�Fp�1$Fe���sQX� Vj���^��4�|�00��}��d���aAg3y��r����S�����Y�@��zK[�qT�V��ux_�����>��{�IB_��ՙ�/L���T2�
p�r����,3���Ų7��d1����q�)ב�E[�Cv�ʁ���ځۺ���)��q#���	)	�6���TƔ�L���8�o������Ƅ��}.�j' ��NiP>�
�����-��=�7	y[��2ѭ��pY��:�&�l_��sE&��2���җ��՜TT��$<nݭ�����<�!�L�G}�7C!������H���R�nteW��	���3�ay9�h1�F�����}s���۳���ߛ�?c9�3��_Y�e:�YfTرؙ���g8?�cg-Hl7��󣭂j�z#�;1r���p��Iٓ�C���M�5�[a��o�/����(qAe�ΆU�5af��  �v#1��*l�E\��L�쵭�f��y���8M+�+��廸d�9�Q��]���v�9r1{ ۤ����6Ð�l�W�[�`ˢ�~'�p����ZJ)�����q�:��� -0[w���3b��JԤ4*%�ZJ;�� W<��	��X�)|3_\`���eg��*���Q?-q]9�r��n�{�)��w���3}Ң�#JKS�m;U>�ș�$���������+{A���K��� ΃�������i.�a��}�Iڕaw���R[	�����K��,Mf�6&�S?�B�����\)ك�]��T�G������De?��N����VV��
@?x���{0�g9�	���/�8ob����^	���L�s���V����=[�'�دRC�t��V�rp�{)�x�h=��-�cd���ù�f-K��#"�{�������T�v��ȃ�i+&��Myˊ�h�>�t�H{�'�p��q��'~�V^doJݦـD^�'��[U?�����kRj.#ص fx��?�a�Jf����� r^K���X�v�Y���� 8��|�{��E$?��wP���4Uls�K�i[q�OU�� �D�z��2�7�x`�d;��w[A�N�U�3��b�,h��y��P�~����������ه�Aۧ(��~v�a����)%^�,�݆�Z�/|��5�\�|��X��s��V;�(%7]FYz� �A� �_a�?��е�7��|�	�vؾ�m��e��E.&�*zV*��h"ZnIB�9����c�c���	(}+�g���~�g������}�F0��bq��B����Ύ�?h�o���S8��~�{�\�r���9����v��嶀�E4�P��:h��x҂B�6�=����Mq�R9��@�	�>l(�8�8�S���zP�<>S��^�e�8��Q���I�a^v�@b��>Ul_�.���/���F���5�c����D#��TM/rp��Թ.>l`ϊ^\f4c��{`��ͮz&���HM�݆�[�c�TP�����#�X�##)Trw�C�*�/ς��O�3,`o�~g� �G��[ɳ"ρ�v��On�L�8'ȴ_���� Ŷ&%�r�h���^~������<�ԣji,7GN}56)���lp��J�1W��,h�o1:CI��/�����{��,��*��z�V�2֔��\�?鑉M�e��^Y�闿|d��]}z��Y[�[��d</��^�!Z��-�&C��c�&|�"l��j(�ї
יeA�?|���wl�0%�4��Ҩ%�-yrLG*��]�.�W�i��B_�Xǎ2R�,L�#��}�ѩ]%�B��_1a]ڄ����̧�d��l�v�{
�`L��a���"�o�8 ��j��I��t<��[�^��A� /K��o�T$�&��E���ڞ�3Ѓx���VX���G��
'��k,�6��F�QU.��;8�����n(��X�u8�o�<(a�ŤR�R��70M>0.�R����*�a�5;@7��v4zj
���?H�=OȚV�`]-����_�kuU�7j2�c2q��#=�P��`�֐z����?{d�������@�h�m�Գ9�&-Z����y�yP��t_��{�o�)Qz�΄��ߝY����V��Ӊ�F��Q�T�m1w��#�XE��'��P]$����lճ�H�+�z�_��0�˦��-dRv6��`E]2���8Z}��F��D��ܱp�I�Cr�|��_�����S��̔��|�/�K�f�L�E\ۑ�N]������/m�2D�̣�a���"g�kec|�'ot���Hp�R5P/�.�l���LA�K��r$� ���"�ef�5j���/��/��׫)2.K��P�):Z����K�^&�X�]~z�]�pk�T��.�c����'�w�Y���LC�ڦ����f�>U��#!5˒N��M,���y���A:eKkp��<\�'^��������� ��D��>&\Ԅ���1� �+l���O���QS�G;jSA6!e�^-���� ���&���R���(�K���<f��4�-D���ط��/�_�ԝ�n���P/���u$oZ���yM��#�L-��2�T����f��Mz$hc�P��C1-5�}���a�ό�ءOt:]fD��\��c��9�>�%�e_��Y�!/=�����u���XS����'bnXy��JVu�xl�����E���i�씔/��$���	<$>�=UG��T��?^1#���8��$���ՃIu{.��.=��4�/0�������z���?��Άm��|Zҗ"�垾�佺�2E�e|�0JNmi0}a�'�+Yr`[oJ�B�~X̓uֽ)r!e�������2OUn�[e]aY�U&���8��l_��X�I o��n+�,�T��pL�����%��y��;_���n�o�'�l=���)����>��<Mf�TD��e�5��d(b��}��"���p)�+W��a��i�Eq�N���G�+�́�0�n�M���N���a��]C� B �N�*�D#.���	�}��Χ��*Q��H�bำ����I�+E��3��w���Mf�u �M���],ʕ�CL�g&YC���m]7׈���3Y�\�[\nKrq��5Rit�\_�,��_�҅�,;A��V�l\�w�ߔ����B��>��]=����%F�%�5�yv]�����d�A��$�@������#�]M3<}��,a��#�	�Q�j�q���*a���.ެ��]��:���ԠC�2� ����)�p"+�Xŵ�q��H��}����R��*��wQb������z~.k6��]\u�t�K�[8�>�4)Bi��Vꒉ��M)�
���QZ�*y)6u(�0\�XWn�L@})��ǳ�4ʇ����E�a�I�m��*��[g�ͣPCq��-�k;���N�|C�I���8��R:�|_ J��q\5l�",F�W��˅wZi�]��VK��(Y��"�R�<8�m K�v��3�qб��
�����(*��t������Ll�.b���|ߴ����}@��)PT_܍c?t�]�x� }��9LU��� ��W�+�#��ծ	�n�UvjW��-�!�o[���D_��zlۅ���Qh	��GTRw��mD��e˕b�{«krC`@(��5]�m4��aR�0 �Q�U�1;h=�u"�ĸT�^n�)g�f�������u�F�s&k2���"�aB��2=:����c�;��,O�7윞p�Ф���B_��y��<�Ƿ��;L�Q�c?)�vAIZ5��+/F�̪�"'k���|c�oqT�
 ��ɉ`�׹5��~u]ec��ji�����J,��H���4W/f#?�6��2p)�D'%�t_Ƶ�cϭ��	���-g�W��՜-��F�̂�����E�K�aI�jFN�\�Fӑ6�E���ëb�)}�G�R�a{䥬�^��y��q1h��-5@_/ԯ��>3V�;T��\�n?�I3�2�S��ˀDA���~��t�#��_�bc-P}Y鎴%�d��@0���N!���Vƌ*�+�	�e5NE�	=��ؚ-L7�����pf<	�B!�]�H%b�d*R�gK�`��.ri�~�i݃2��0~5�l�D��\AV���&N���r���:��K~`�����������f����6)�i����s-~�əәM��Dm}��Y	MZN�N�+�ۇ`T�j45��� �P�r�`��}��8����J�1�_�5Ü/p�S������T����D��j��><��g&U��L�@�.�ʸ��~��!@��د@�,�v��M�C��m�\�� 1��F�kD��9�Js�o|��8���Lѽ]�>���vF8�*��`=�^�?N%���+UBxji[�։�x�ބm���x�<����8o^���3��p�,D��jPa�R�UL�uG�Zr=/�'�ϦT���2 ��}A�!��&��t?��;����J�������əziq���ڄ�;D�d)��ᄞ�V��~O|�J���D�����A}JQ󈥫ʇ��4s6{���ǐ���(���-�4��xC	<��<;�S%�F��L��B��+���)��.ʷV�=E��t�q�l-�3[��J��|3=����5dsгd,@qʸN��s��Ʒi{l��y6���P�R�rQ�8������(b;���׵�c �q�P^���H�t���J�+Z�o* O �ݨ�o���A\2�ˡ�Y�*S��;�O�6�������E��I��$���j�Z{�
����ֆ8v^�a�^	"�@�BxI!Kn��4Z�-3��J�����6���z�ŀ˟�N5x�N� ��ϑ��~�1�0b*~[��2JM5Tqf�z���X��@�������dZ尰�A�����%��kb}�Pyg�&���;��ppDTő��|ϡā1�L��B���m`�2n���*P���6L+�S\�T�*���eg�
�0#ϴ��B�8ﶘ��_�hq�.�z!G�/�n,l�����Q�:�ȅ;���P'~0h��ã�� >#)�6f��n���W!,�7&�b㧋�Tk!�_-�o�TC4���*�g�4�Q�9��'�f�:�k[R7�%�ısE�P��KaW��]��J<ဲ?�l�r�"�߼��m���[��"��ت�s�@O��M.l�t���#_	�4��a$Փ��>�]�&�Ζ*�X,�?���w������:�7@=3C��<u�Z��N�H`j��[�B��}`H�i���ů/,Q:�X��t���'7ax���C��e�Y
K'cGW���X�؍Q`P�=�^�}a�T1{	��mq%��6��\2���6�[~�b	V|�3�N�]�aG	E	�^-��,i�>��ReT����o'�Ǝ��]�.�(qR�kvs�ӻD��0�d@s��K]��g�{}$d
�$Hrw�aK(\�ګl���mż�9�i�w�
��55O���}���`�`�Q�a'�ӣͮ�"p��o��Cz��E��\!��]V�F�, (��zoON�_��y�|D�އ'^��S6�=����V�t'5.��E�V�8�z!^�`��A�>ؓB������8��z9��\'h�!c}��5��j�Qu�l���Y��j�9����Mn�VI8n&W˥'�k3����>+���IT�����P]�z��ۖϚ����H��"��:٭k+�5.""��_��Oa�h�1E|:į(pkLZ�
�s0q�'�j�"�����y_<���<;��D얯��K����D�-(+TN�o����!�L*�k��!�-qN`ƕV?`i"�,6dJ��~L��&0 ާ����3��5e]`�S���\=��2{�|e�9�
G����9�y�ĭJ`��DVUc��>��%ؒ۱�̸O�<��F�9`�0��IJDM�ߥ��U��41�U��!�0��v �c��~SH�ǝ(�I�dW��0�� 8I���N_��Cqw��R�Z��u�,hO�W���k"ȕ�2G��K.��v_�qM�di�	B�x�����?`AЬ�:���S"������#�*0N�C
��wĊ�Λ�@�:�������qb��� �ZޜO@}���%�)����|��7>ùN�qV��[�x�d7�*��Ŋ�pņ~;:|Ia�	�O޲6ķ��Nk�������1�w�i��n7g~��<��"��c_�|�K6�B{��8-|�Z�K$>��H�	��NQ:G{m4��%tC�Ը�B�:�CZ�/���Ǎ'�3������o]��� �a���"�8��G�Teo�͡�ߑ!V͓P?	���V1OoB�����mTp��[R@��b�dlY��r��2�Д�����2���U/r�R�
[���e��f���1<�L��59��Un�\��
����Lr�����H& '���Gv���,D�Y+5w��4�-��ӂ �d��ڏ-��13yzl�w�"ػ��V���r����b�1>Q<��Xk�Z����#�>�:1�'+Ġr]k0���gͻ
�@#\���#����*<m�p�{p��?9�
·5>ȚԽG7%��4uG٥�w��'?�v�<��Д�L��1�J��"��O%�Q�u7���D8T�%g�3Y�b҅H�����o���a\<dS˲1�dm����Y�/Mv'��\X�l"�{�����!��Uo��I1'�[�p#&z�G��b��æ���.�j.	�D��U�Ɠ�S��z�]`�>C�ۤ  %�E���3YO�߳��F��y.i��$�W��%~����M
$Ķ� Ɵ|>mM)(��r!��W�_����1ʠ a]1}8���a1��I.��ꟑl���V���_�s������FF	�{WU�1,=9�z��4�)W&_�J��Ama������{�8?#�����_���	��L�l��9r�y�,���;vs��-_�}Q��pd6�]����#ፆ�K�ӊ<���@��e���T����,��>������FI>a?���3U��2����Uܵ���>^�B�&�����&��^��"\�D��wO�ut��^����+�sf�����Q�+P��e�`�.@���b��9FfUPZ��/#�q�3<�ʲɏf}�}y~j��
��z�YG���-D=qbqo���1;�X�&X�UJ9ꚗ���A_w��f���
�-�[�k�@I8a,�c�=n���Ԛ�L��#�L�� ˵I��A����$vj@͞�n��Es��l�n{�2+?�Nt;���q}>�����#���ԥCѧ��}7H�}�┑<[Q�
��\��{z�,�Iw�w��|�B��y�s��������2P����c��8�\����{��0���]�*��߹G&�,5�aSv7����@!���fFv��̚�k�(��YȎ����Ź�F�2�u��d&}@�[��	��zQ���m�^}��)5����2)�_X���D�d�����M��$���@7� V�vLw�����إj���] ��)Lj�qm5եw���K6�R�e7��r5I-{�?n>��31�Z�%�*���(]���/�x~��Nx�/J5�xXD@�����%�^��2���_�~�y���?���m=��%�ؒ�"0)�4��"�����ԥ`�"V�щ�ND�����qr eNߕ��Ds�R�9��.����r�|���_pC'���c|�s���^�%���}Y�i	�������G����qM���b�ŵ��%W1�Fքh���|�{w���J�]$�҄��V��u��i%�]��B�r��R*�vOa�_�wr���X�|�\�N7����?Ջ���'%u_��ӄŮ��
��R��u-p����!�-�W�����G ��
Y�*���O���wF�dW�u�� ��
���9�"j��LB���>(L���q�d/I��Rs ��h�%�*��A�lXr�A���e��:� ��H���~�*Cge	rXD	���:��*	*sJ-��u8E[b�J���!�^W�a��� �>��wʅ$�S��\gS��3�c�@F}E�`]��ɓ�3$s�r�����?�$.5J��Jt�F�4����)v��t	�F0�чo�wa�ȧ׳c���:w^2��A<Yވ�G�&2	k�&���&��z�@�v�I�v�d������1�:����ρ��k|ZM�Z�<��6��>3S(�q�շ�~Q�K�) �K@���[�n���g��JZ_ �5��S�݂��v�כ&E�Y�	�ûz.�/&s���+�Lr�T�`�7	��؀�V�%�ͪ�LU5�q
K�\������8+���s��T�� 5�؟���,[�6x�i�KA���)v�^D�����;³�
�tVb8����w6���A�������E,/�S�׋���]�D�z���0e`Խ�c
z�|�5\�ff�ť�Hߥnq��ޤ�nk!���ZoJ�.�����`[8O�N	!���GOp��B�v0����zzN⎤��-U\��T�OƔ����{��D���	�p����٤�\�����. � HoҮ%���4�o��� ��?��$��0+���^O"U�6��@:��l�p���D����+���=Zk��Sg(�Þ� E��Ӱ��φ�8(�C��]�V�o"_5���������o�i��ث�J1�ݎNB����o�@��C$"�^K���-8�9�s�Gj�K̑)a��E��x�ԮN�t<�X�)�3��@�gr���
1�/�k�i�^�C�tB@�T����9Ymw�=B���K�ώ:���3�F~�z�6
�F��f�wZdy �=�wAְ͎̞���ԜX��#�^w'V��`��@���AQ�Rר�ȍ�&l]��s�R~���H�F�	�eU�/�ζ����_n�9�DKwQ�@�����e�C`M�Ǉ�������.DX\�*�޿R �% 1�G�o�K����@�F�ݼu��:���S����`����!��؛J���㬽]����A�7ğ�{9*p��(��>v* ٰ~(s`��l�%bi����M�% ��:���C��Ѓ����eE�L˵��[���V>x�z��>����Lz-07\rf����P�zµ�v��|��Ӂ(+mGL� Gd����T��=D�C[<t�����Xc�YĬ���W~�Zk$�4/��ζ�I*�:��s~�ƙ��P5NR��<��~;�n&��H�H��5��-�s�C���F%`�:bρ����[����e:�w�@ޘD�1V�}�:�5 *���0����}_�
��㐦��Zi�^�r=��M�� ���h���B<j!�I��	����l��fQe��60Xv��i~�A%�V���q�,S;[��iR~�ʹ՛��W�ߛޣ�IUSAS�.#~gRƦ]V^��e]�?h���b�j[�P�-[ݬ���Q{�m��Hk�ںq��.��+�Dl��Ƶ�/��˹����	P���.�m`&k�q�ΔtW��fCLi+7E��*�u�ѣ6?������:Zֿi�d��?�)��;s"�)ʺ3���$b�2����%����!��̯C�)�T��M5z��Jm��9ژr�C��g}�$�O�?^���]����jí�.=�d�%��L5t�`���8�H���[*��J�nr2���2�x0Ʋd�K5�a���gGy���ۗVJiY��J��֘P�I7��H���R�漋xȔZi� |:dcW�ȍbJ/�V��TI^+aU�w)�5�F�B9���\�L5�}9��t�W�_�w�uj�TJ�DŃ��t�x����gL�򢯶�:W���Fs����,�E���P99�p�#Ԗ���h�BCR�H�]L�mb�2kn�|�p!�T$���Ū°�g�[1�ت��a"1'���EZ�WxԮ��L� ��M5�k���x0�-:6����t�1(����V	���-1�y���[@���U�b�~9Ig�s>��HH*�~��-�*>�x0p=lCP�/����`'��m����S��F�0�U�ۉd�҂�Ϯ�k������>�-E���8:�G��� �w�NG[jȧ�٢K��gڐ�Ց�>^�!-�����s��_��˩ف%�=h4i���e�/��Z�}p�V��8�o["�7A�fb��Ȃ'��S�y���ja�q��46�����FڙZ2Gz���􀷃�'�	~��݆?z������흸w+o��/㕩�^]�1��DkW��[���T�`�o.~gI��0�"��g�K'I��B�fj������l˥��Yd-K���y� �����ȃ�:Ƈ*����B�Y�;� ��q������� s�j������*����*���A�>FH>���&��q콊��|v�����3�4�p5��w�»�:+��B���Kw�=i>�FV�j�2�CgC����W�d;�-\�&��u�).�m@z@����1���������`�ޤq�^��9���¼����Wf��'���8���$��r@�Ւ�Ƌ�� YT�xC�����{]�[�o���K��>�"O&Sw���Z�`��:�Q�n?9aj���u�u�c	)�������&���c�R5r�\l\�H���\�d��p�ϺK�%1���� ["ù�]���OWogU�^t ����U�k�Q���{-�yg�'����WB n��g趥�{�/ h�7�d���]�KsU��'f�'5+�!Zߨ�s��Bf;ȡ�b���M5���4���ǙDf&��o� � C��Q�vL��-?��!g�/�R)���/Wmo=�SJ�
�4��Pz�{qj��ǥ6PX87p�2�����3*�whiB�s��pEB2��\zNp'WM�߸�;�_��C�{U�]N��l��~���-?GشR�	��7N!����2p�2�_�7��l���P¥ۙ,ƣ�Ʊ�r�~� B�Jhy�~:2�[u������n�P��R'i�ɽ��PF��nV0ƴK!���|5%�9T�@��.jd�m.y����Re�,�K�h�|=P3;ߪx~�ίaޣl���b÷�z�rUc�@�\�i�j+
�6���e��ok��r�)R�6���o;@:;�Mq!vܳ�LAp<�Q�ߧ5,3����������j�8L�&��B������hs�<\^��c(�-�dS6$i{v-��p�J��U�A=c��fIM֎�M+�OX{c�0x�9ͷ˯s"���5>l���>�u�"��P���`)0��Px��P��x^�����rm�JK��~��HW���M�� �9��T�'�]�1�S�d�Ҷ7X����K!��}R���z�`0T��_����)￀kA{���bV`ui� o1�:�vr��"�,ݿ�*4�?�8F��/��D@Gh�����0��$�!��'�j�	�N�&�0g�m�+�g�="΍>I,{C-�S��&Y�V���&��
�:Ub�~#g'7�fj�\�@����n参z�w�´�=�mP������l�<�I
*��x�V����*Z<�O��� �ar���@Y�TP�?U�}iԹ���Ą����a�ё�_ql�K��;M�$Te+D,��A6�~��`e}S�`�������g��
DX��sҢ�i�SAv?��	�N�a�m]
m��W_�,}>�ϕ�5�Vg0q�y	]fq�5 R�`9�`�OF�n�d�"s�]�n��i���U��b6I����z4�Ry�i/����u'.ض�/AXw���������[���IRRZ���Pw��)��{S�i�\�4!#V>aO&4#)��_������pG��(�'Ӎ�^Z+ER˖�Ş���d_ͬG��F8;��֋�>�Lc�%��:�Vم��|�|������&8Ķs͏��w�,_%1�\Uw�=D��%�<������q�H6��[e��oiЩla,�7 5���/S�������M�]R��?5a�J�
�m�D\P}n ��+*�Nd�ojg�dmY6�����oL_N1P���{-K��$�H�_&�����-��'�~q0��P����nA#�w�Z��i�b@A����M.wz3j<��o�94��R��~�@�eCb��R�����$Bڿ{��޿�A�NL��E�Zm�"���+���ɗ�o���4��;�O6����8�&v��U}��PL��@����ش2�-�FC����&����;�=��7s�e,��YA+�7��1�@m���ߎ���8���6(h��[�!D�!���36j�"lk����p'��̎>"���}�1�|d��Lbا����_c5h�1��=�ߛ��g.�-�-
X7e'B�q�%[�Dz 	��ٍ�	�xWQ�4�}טh�^1ｆ3�W�R�G.H&�x�T2g���	��~���z���S'Y8l�M}�[�=�Q��+[�C	���tS���T�fw��rŽ��A��ac�J�j�y�6��(�Nyϊ|Y�����Y$��.���۟��;ĠGBn`Im"!�1@E;k%_��b���gӠ�j���4�n� �5|�h��s[��fڞPڥ���m-��dwd[����2	vX�� �9c���r���Kst3�cC�����63�?z��uO���<���%�w�b���u�q�9НM�	�H�dc;��%���!�X�*�ޖ7�$v�I�_��o�ٴ;��5"k�������.���U�>�e��d�Ѵ��%j�o�:��7�+���7 ��i���¥��4`>#�M�?d����h�c�')���+��y��0ʱj2i3!hl7�ԛ�K��ʰe�L@6�S�9Zl/o�D�d��e���6����k��49��Hw��K�_���
th���|���E�7Vd��:��2���R=���5yR��N` �ɗT!�L�vVp�v�mrߎJb���]�̇��+�k���V���,�)3�Bނx�{lB y*�k�-�����,�=C�t�_�J���P!|��a0��_�T]� �d����w�o+.E�e�4�E��g�rN�ɿi�����*䲺��\��@k�N��;�����qR�2�=Z����Pqt�s�o3�h��>;Be].ӵ�qo��49H�\ESl��T���+合p�q�����vh�[
�n��/	�|Ñ2D%�ۚ���W��л��8�q�}�����Dq!t|�w�U��e�\v���}������J��e+B�{��������~�&�����}����!�k��J�:�hRd֞.f��oZ��H�����H�0�'��2�:�|�
�o֡��r�O�#�<@���M�>{�W\D�+���8.�!R	�}��g��v|<�ϑ�K@�5P��=l�8>L1Ҙ/���m+�p����;�*sô��ӹ!x������*��֨��"�A��4��v$ m"�!�j ���;n��#i�i�Ԩ�pZ����|��A0 �h�MaGy�s�_��	�0���j�vBS��� �{�)�	�����u��H�Δ2b>��� ep/��'����D� w��Ir��&�\�Acs'/ ���|��'�C��5���˫,�d%ϸm\ǻ��i��.�oKw7�CH}���5���P�t@S���16uK��`�Q�P˳C�&$�c<�f�TF��N�(�p�]�[n���b��0yI��+V�����`ڶo���[I��2����P�2���	*���a���_��i�e�)=��{����&Vԥ�f�NF�{��V0�^=�m��Ͼ�����U��71V����ΘϷx�|�u����%��wB��5�l�P��|�&�J�'�L�`�u�ؼ����&��h��i�Y�S���b�p���BZ���Y}dz�F�N6@�(����J� L�F���2��z���w�;�����lz��X�"6��]粈��۰�!ĝB����.��$mh���x��I����R���@n��g-�R��(��!�D�v+��Pҽ��.Ũ^�\Q�m�%U�̹�Q<�*�j|�1�\(�Ѫ�;m�1N��$��C�v8|k�<�?���G�aF��ֲ>�����C�@>/.)�[B>iW=�w�3���)x��]!ւg��H�Τ"��;+R�5���.�PX��|R����6Tׄ��q]��R�@nt7\��S6��ԕ��N��t5��@Q�~�Ȯw����X��T�l�($M�ɞ!��T�Rb�>�B?�i�����	|�����4~R�=�g��H��;� T�}5�x�[)C;����(�@�QtI�XO�R����� $>#�b�����1�S��gW�es�������:3����W%�b�%vS=Г��c��ҕ�ȶ�Tz�%�T�\El�V��"��܃�X
��VG>��I��a!5��;>)����?���*�����n�zu�[��|*5]SZ�����J���e�>[�w��9���ŝF%.����O	�Φ�C�#�A(���*.����]fcu�гb�b"m_~�r؝'�Yj��ױ(V^�a	2NI�<��%�`S`-Rg�f�_�&��w�E8�	)�2�+��G����fg�c�q-��)��֡=���:��8<��e�}/梍��O��˷U�[������^M��|�׻9����t�֓47�2�}�U������Њ%^��s�
������7��~u��֌Ǩc'~;�u����{����(��p�}z?���G��kf�_�eZ��\BrE!�zf6��/��O�֐QǪL:���@F@�.�nBI�z6���L&��G��]Xz��{ѳjv��rS��ۨBy���7��%�-��eD�cVٌs C��{E�%����.����N������e��|�ՠ�Mɚ��-��ǈͥd�'��TbL�!��F�L�o���F��RM2�qZ���iL�ch��H�`�p!K��R�KR��֭��:�ݙ��4]���F����=�6�n8+����Á&�IM�;�P&��
wQ�m�|ݔ�5(�;�����u� J+�LNR()2���85U�o�'�zw����Y'A�q˭' ������Z�����
��H��J�ڟ�WPI�5����R1���Y &_I��#��xޢ��Y�C��&D�==$fxM�\������s�f�A��$�Yכ�O��T�1.ȉq-�/~@L�f�ay|`a�~�dPԜ��&j�-����T��2(ذ�E��M��Ĵk��|��P#��<�? ~�����_5&!sT%-����zk_e��%��4�oէ�#O+T��:� T�Hw����Y��v>X��YM� w�:,T�g�Ʋ�WX,d�qH���Gvs�i.?|�ؚ%��~ë[i��/�]�h��Q�).ngW��RG���G�\��F�G�:'kx���us)g�s*s�/z���+u��t%L��Ͻ^�����y-�9�	L��i��Chs������k�}ܬM-Ka3e�+:W�q�����.j���K�O�>������B�#��|V�AJ�ؖd0�w����`Z�т��u!˳�+�I�\�~�� ��������'���P=>6��_�Ə�{~�uZ���I�=���M�Q�zXU_|YO�B'k:Q;hH�Б) 'Y��y��99�2�ȉ#�vW��j���Z�,O1�6l鑊)3��f^��r8S��X$����-��JG������{���Td}�υ��H�*9�W�u���F=��+`C6A���u#������Vs���@�RT[�jD�ű�a�J���B*�<�4ps}�q7�l;Q�)�.���j�$�U,���1�T^�®��c���J:Pl�/�`l��_��=3�G��x����Se���$
.�_!�I�fw��,T�|���驁�U�e����$.T~n)����t�I�6���^Fe~�o������}+dE��a]�ԏ:z+m��J��:]��LW)�4��V������t�2�I�O�nv���Z:���sd�A~�[Y�r�LMւ`��;6�P�����B�eyq+U�aJ:a�Tc��WV�6き�ޜ�l	�������z���A���@�r�H�)3{��+%�ͧ�`%-�\�����P~��J�H���ICw1�������g��la�/�����2<��"������K��6�)E��?w�4�)C@���8�
	BE�yd^ �09�͐��|B�]�,�7 �,2[�m,vT{��z��)��J7����	��a~w�����$_��Mc��oY�f��r�M��X��&ө:+:y��Y�O(P�d�ҍ�l�,/�{�3`���QS�S�v=(ϑ�C/%Z�H��6�M;Α�ϓw8�|���彜���)̿�U����Tt}��j'0=�i�h�݂A{M�}Cֳ��Ҝmp�gg�=F����c���`{I�^���:}#K.QWj4����^�II��i�Kկ��V>�:[��G^i�uB:�A�W������8$��X@��6�Ł#WXl����̙M�s�x�w*qx��)�s�6�O�W���=`�pX�����ρ@�$�+�cJIؕ���\��L����r|�p<�������A�.�2������E��s�9�r���eWË��B�q��pw �����@P�/�~�Ct��C���4;q|C��&�E�S��L)B�u�s=��{0lS��r����x>���r���q��ّ	��,�s�:!��Sj �Z�\��]2�t�'*1Yo�C�IwƗ��e��W��T֢�B�e�"�]oT��x}{�����8k��]�Ԝ�a%�ʸ��9B��c>���.�����H9�^q�����M=ο�A &���]a����\{f]	�{�Bu��!A�#��#
�B���!N��yz� ���M�U��n%)\�ŕ�9Zд�N7##(��!K���g�Pw��)%5s�#��hQm�l����b�x�F��ڔ!����	�&�ed�L<�1��ސll�'��[���m {�fb� ��Nڴ��r�_T�+�_�2k�@�N�J��:��l)ՒѬE��r�5���ظޢ�G|�Z�OVPg�Hc*���	O,1QF �����{�6 Hb�*4+^��a��*�&4
E?b2&?�=d��OC��c������2J0QA�u݌qCוB1꾶 �(X�����
j��wI�S��ɮs&$�kׅLr+��陛Ӧ�	<	�������;��F���l��/gqH䆎�L���d�ҍ������f��1+�f�$�󡱚� \tcKW3��F��~���;p�yc!����5�@UZk�{��G�g�0��0,��gS��������J����ch�FsT�Y��s�^��GX��X�'��u,}��\rap�Y�&�Y8�0!�q�D����X:;�[��=<2��	~�]9��混B6�:w�M��7�f��q��|�j-�fiIW	c��߻�6�����(��"�sv��y��[K�=.�c y���21�'�nM"`�����ds^ݱ�]g,S1�ͼ}-?Ț���v��t7�����c#����9e� 2��X'=��yF٘��0�v��QfM����+)�T~n"����dtb�I:��dk���~Z�T���̧,�"���|ft�p�C��U}Io�`�]���(;0dst�Љ ���e�$9u�jY$�VgM�0����]�ŧ�z��kjѭ\p�L��'U���_L�G�(�4�&�h˗&n&��G6�_Z�6�f� y f����L���� ~]y����Bd�o��0�B�fQ��))JVJ?M*<PF���'X=��_@��F<���c����>ƚ1荞��Q\br"�#��T��;��@�O2����z�T�yT��se!����7�F���{AU��H�56I�]�C���ײ���`���(2x���t���ˆ*H���y�|�,sJ�v���p��zqv��[C����T������3m���*�� :}�yEeqv%�wx]��[�O�D�t��7���h3���/���L�q����5Zs��~�����nMW0� S�ںꐞD�Ydz��ګ�[0�.#�ȋ���*O/����s��V߶T+q	T���Ԍ'�OφTc�l�>�;��6�u���暙D�͟�A��8�<� �x��Qk� ���=j���j#L^��)o�,BT��<'������r.���<P:$�sF�����ܳ��uP��|��J�Ge�g����)�ނ�l���q���nu<	�1/nN6�:�Y
��eZftv+sugl� 2�P|l�:)	κ���0�'+ƭ�5��@��6����d�I��F�Y.�#&�zH
Q�뮡�yu��Бm����ŦY�9z�/E#����r�=������حH��z�ӮS�B�1�j��tH��f�jh��B}	_���L���o��^3's���CA_�Ë|�}�y-cB)g�l
�t	y�~�Ƣ*M�t�n���q�����: b�y��Ѯ'�IM��wx���#��/K��3ޝ�[�H�JP��/5�e�p���+����.��ӵfl����
�C㣓!�S��Z�4+İq��j�����l�UH���¯�
�֖��K��:�*9v.<+~D�����D6<L��Gy	CmX�X�-
. e�����%�%�K���*��ܥ�����!e-9O�a7T8�?�nIB^�)(� �p���[��N
'��"k!��Y�ѻ���Ƚ�yZ�x�g�Z��n�j(%:ږ�tV{�K� ܏:\�T�"��� :��gz� ���O�~��N#�O�_5��䙴�_��5kn��rAM��oi$��Q\�K�h:j.F�μl��[^�OSJ¸ѾoB��b��ɶY��p.y��Օ)P�
iCx���c��dv����BOo�RϠ�Q��?e��C]bݎT����F��v:��j�i���ŃSAA��
7ax5�0/��hP��Pz,��$�_���Y�~t�3L�8E�F��w�M���aTק�!�|u��!�XPCӹ��j��d[{��e8b^��H�bw�8K���I�I\��e��:�i�6M-��g�Y��3V#b~D�ڝg�c&�1;��������Kg�w�Ӆ-�,��b��<	��W����`n��N�*|c�6�j�M>�>n�u���
N	Ҹ�Aߘ���dnu��c]u�%W�)V1�I��U����P�~����J��C36;���n.�fo	�Q�@8H�PlA���g��-�J�Fܛ0/d��Y�#��lD�',9djM�H��_g/_$W�n}��y̜�Xe!�5��L�����xǏ��\����\�@�嗴��:�v�z�%��o#�U,�^�t�9�]��@���n����el�!U3�K���+Μ~��gmt�a�_�5\�C�v906 .�KIhτ����NDE��+�Y��|a�td�a�g�n��O��M���[���Xca�} O�5#Bڬw��t���Z�:�z��$~w{Ks�����ŋ��્���沷��i��~�^�[ab�U�XMtXp&F,A�k��&2�����!���G�T�	�|Մ�7���c���l��P��.:tq?g�'|s��+��k��=�-��_y�����p&m��4��
yoY'�A��Ղ��1<����u�	c2��9n2����Uƿ��v��ޣ������2��ȋj��v�� �4�[�--��ٹ� ��ypYk�2r����Em���Q���H��xBJj�7��ΜE���L��GN�
l}�i���]d�s�X&��́��E�,���9�K�oFx'�0EeI
?`]����D�iğ�a�[�jS���ᲃ-�U������D�Nj�SǍjIӅ���F�%lЎ�]g�+һ�`%��{�P�WL �bd{̾�����P���rd�x�'ve��''�� (���'��Q�/vl�)Wnϐ-�q�+��d�-���6��T��L������|���@��`H�a����������#��FV�[j����&��C�xX��.Jb57����>��0�=8N�i
^�ۂ��.��, �}������ʛ�Px�W�uŰlr�J��R;��16�S"Oz;g���EXH�W�'-b&�!�T�h
Z�D�!Lq��d�:�/@Խ����I�<2@�H�L�B
!r����耣�&���!�<�����[w��p[�7W"Mmut_��5�:�*I%�9��b���63�5�&/t�Ӭ_�j�A����{��*HI!uC��:�T`\�M���#�ܜ��s��}����ܪ���G��6����>�9m�'���p��v��*]��\y���s� /�X'9�&*��-`S��*ɹq�ڛ� �)�����Tp��S��?����׋Y��:$����s�X��U��|݄�1Y��L#����Dh���j����iޯ�3.uw�r�����{��;_$7_t�Ѫ�1sD!Yr�&x������{�K���1���ܵ]X�G�g�b$qJ�
��8��\sen�6J{0cfĽI�z_���)?����,<e�WAC*�"8tj���@����<@и���b���O�xP�/�T���9c@�s`�� ��9�{�<�4j����Y�/L[yD�i�z�F�#�2�Ӻ]/��W���${h_��-$+Q��C�;�k_��*���ع��W?(D$B�>FR�tz43��f~�a��9����%�U�Pϩ��M17�~�|����+[�H�	`(�'9���f��}t�;'3�g����?;��e|8�1e,:�t@�+~cr�~&h�2��7�ub����^�q:�^�b�zQ��:�Ҿ��@��$z��#v>��i��,L��y�o��:ҋ���tg���s��@t��̓�H9���,�z����ü��UQHv� P`��2���$���N�U,�92����<B�4Q'�)���������L?yo��c�c�k�c�F#��@�J��m"�e7ܛ%���Q�q��|���ʰv�ќ��nĳ�s��G���Z��i��,��ע�\��3�
�|JE�ac�}ŗ��9g�����1�}_9�@f��s�.$�b�$���@���m{K���&Ś�@Q'D��spD��"�XY�a��A�G�����E���+MN��%(��ʘ@>2��r�n��K�fo�����f�p'�����Wg8 P8�q������6�~�심�%�����̨�"��g��}Dd���_5��a»PK���@]Ʀ�tT�n�k��,D1x�g�i��H`Ù�����?�Vc�ql�x���#]D� '���$���w�����lcLV�oL�A*������<��HdU]��� z�j�U8�� @0�"R�PplEc��:���el���1OP{�Q�P�>����=M���}>�G1�r���/��d@��زq0��_Gh��/���qB5����6]�E�=��2�6�e%\�IM�)�DM
Y�KO�&l� �Pq��na�@oi�����������U��*�wo�r�S��I�]�z�Ѧw�����!4�I�<��/�`��$b��U�<�m5t�\���cd�u�-]1T	y�'��s��$�]�L��h�8�GD�>|,�c�[�r��p�
�*L����Rw��m���<MI��><�{��R�	�ՖJ�9��Fc��9����y]~%����u8?\��<Z@
��R�yW�W�j�MЗ -=>���$B��d�G�*� ���uc���:Bm�@���]g��.�Aj1o$>���
�Ph������CQ[Y'�nQ� �2�(4�~cCΐ㑌�A� �T$�L�Ψ��Q:p�2�H�z\����_�����4T���Z�x��D �(��Z�&{�?F�V��L���4����>d8�������.>��&���0���޻�Eۖ>9�������o��I��h�<�Of1���f�կ��[�5���ſA�� �6w�����N��eF�u������]M����6��E ���Z|Uߨߔ����	�^�k.��G�s�C4�C�C+6`S���~�HSW��xt4G!zi{Ra�&N.Tj+Ts�Β��G�-���������F�{(V]쪛b���YzBD����6��6q�,�`�t���N�7����պ���scmd�lM;[��M���=���8�rz���w�Ye�$c��P������^�!�ִ�\h2�
?~(���ٙ�>�9��?��}�0N�@k��RI�_�L�h>��&2�Lj��f�5d%�whѬ�ѰpOc��I/)�b�Z��$@��� A԰6��t�����p{�B2�]�&�9�v)M����^�����[(e�hW(�M�K"ތ�pIG��M�F'��{����f��o7ׯX[�������/�ګҴxQ���BmU+Ʉ3l�
�g4H_t8)��V�a�Yg�{��L���}��X��D� �
��vX*�#%�,��fy�du>M�յ�\�HQ��
��?g�"D�=�W�
���M�m0�#�*�o���APyQ3կO����F�MN�06,QcGMמ��3�#���p#U��g�Qa�v�|���
���^���y�þ�F��(�L���+�m��9�%������RUE��;�����T�3����������YqluO�a����<��N�NY/2�0={��߾;)T�ʹ�C���	碡oc�6!H�ު���� �u�(���6�@�{?]��`�ΰ��S�������;�G��̑a4IQ�!�>^��r8R��AK�)LK�ZGO�hK��Un 7���?$��nk�J4�!�ǁA�JG+V�q�ҮDS!��5�Xb��KWa��� +q� �`\)� A%��{a7ò��ۍ�(1R�g�Ji?�N�J��w�Z7"U$��_�s2��仚+�������@lN)^v���}	yW��
G����&����u�}ur����%��ʴ`�s���~���s�H��i�$�b�/	F@{}��=H�'�
�z[_�W,o�;q��2ΨЀ�Kw��`)L->��l}��*��S-ˆ�TAD;�*��H�G&<�׳��,!�sF,�G��
4���3��Djl���)���(���������?[` �ӈ�;�;���/	J�������������h@�ۡ�5
{��} F�fq^P	����.}���(�Q �� ��~�r�D�{���[U��H`2J,?t�Ix��g;��5$ѵ7��b�����7cN |��r�;@���[*4��mW���棲���mQ��O��+���nѤ~4��Zk$���#��0$M�Z<�#5y~:ւ�hs�(c'WTXv	`���<zk��pW��=0��"6�U����̝���}�]���5���v29q76-s{Ѝ�VA9:�|͆,4����Z���!���VOU���z��r���h�U�@�y�OT&��쐢/[�<��2u�2(���ȬĲ�����O�`I ��QEH魳B��4��o�R�`������y���c&�xG������ܜ��g5����/�,�������k� _��0�3(�/�~Qdx����U��Ie�����6◨�ӬT'�K��g�\H>��*8K��� 6I!��D�d}TH�kbG�T�Qt�U���9������XSY)�oM�q�e:P�b#q�{�7�?�0���E	�n�{<y�qQ8/�����?�%5j#q��s"4�}�-�XO�XMT��?���q�`Q'w*�nSަ�%4/c�~���`�� F�z>�}��V@���{tM;������*q��j���0)+^f|�r���a�D����_"��=hΡ#��DfJ/C"��P���]o�|'�r.o�C�XM/y@]d�G�9dytb��o���/���^#+E{��jV�&v����#Y����^��[�`�몱|`h�b9�N`?2d�t�uLI.��]n��lD�g��ٜ�áw�2{���T@dIy)=� �T�f���'�o�Qki@�s�]|�Z�t���ǉ.�|=XW]���҅ͺ��Ti�I��tQ�|�#���W^:��7E�i�4����u������̒�R��n�M�\�Lt����W�/��ԍ�2�ix?��=_9i|H>�L�ܙl]���GA�:j�u������J�^m��.%����_���1����ؖsΎ���ہT�R��[˭n(�6d�{�([a�+��p��A ����1�R,��{��(�$�N�p׮��GP5VgRE>C��v�{���GR	'� �Wct�^W����[P.�+2YƤ;�@���������l�=V�~�hR�۸I��紉��������8qY�Yz��i����(m��a4���7�Y1V���\�҈��7�E���RJ�*Z�΍#�`����9��}D�.:Bw?��+�Yp�N�R}=�,��C�D�������Oz�q�8}\���8����fn+�!�CT ?����]������m�폻]-3$^W$���B�G?��=>1��?l�����9��Sq��k~U�P�x!��9M�Q��u+)�ziQ,������XX6"�"[LG���\���b��V5ld�����",__�^���]i��۳[۫ƃ�B�����#��pw:��s�1��?G.�'�$�7�Q#=�e���~�n��#^�#)/ ��qA�_� d��]Ӱ:ߜgoyN!�>m.�J)|u�b�6���L0�(��%<�v�d������8�)T
^P����c3A�@=��3�{��x���Ҥ�������~��Z���Wj ��7Y��#@��n�R.&��O��N�_�C�O�A�B�#I.>��U��B;�D��!�����V>K��R����W,;�V�Ʀlむ'��sc�w�l���K�_jC��m��U~�Ԯ8��s��a��|�Y�R��nhׇ�._��h�1�
 ���6v*�I����?��Ym���
�����Q#��(�C�7��P�f�_��&X�Qb�l]��SyW���6�;�iA�4<̽���YE���b%�j�!�D��[uV��:Z`�M��[3�`SŷE��a�2:T��.^x1��n4J�g*���ғ���}.���Z�����8��j��L>\����Y��v'�t��,`���j݉�RD�s'6��*��/6�*xM�9VaQ\���x��ۅ��Ղq��qW��'	j�?$���$|�R�~�����+{,�j6rHh�j_W,���T�#����U�>���:��zh�fO�>�r'���5�!����m�Y�6g�<�%�?-Q��;Ϫ����	������!$��T֞���ںv�K�Qr{i��FC���*Y�,�Pa�I�|r���h�$� 2I��X:���W�}����
�кQlt�� kĺ&=���C+ �J7����p�B��v�:(̀TEfI/�t�gN8{�ʌ�q�9���h\ލ˟x�^��3������}�X�S0���[��]�K63s�눕�UWk�;�PX��x5��&]OH�~
ԯҗ�I��!*�xt���9n�����<��PY�}v�\?�ū!��;+]�����67����<�C�����G�� �	�d���>&xf=����VW[j��/���:@�,f�9��2LIv������!�����R0vap�eyr�:,D�E5t�m-�u�l��(��h�E�*����')Q@��J!z�;r?�1� �,̦�In�	�(x~�+�>�����.�xo� O;�E^ |�N:~B�-�,��>����\g�ngD�����WW�P �А@�yU�6a �mޘ�`W5�~+�n4��i$�È�0�钶�mo S�ȴu[pD
�7���k�8 \���p�!�� �<x1.	Lm�G
5X�![�f�]QcT�!�w���Y�/�a�틪�4����Wȥ��ǷC����ctA|}&ABK�WF���=MiH���Ͷ1�����S�(��Ԡ�a&�|���8m�Q䀬:z�N&��o�f���?��_/y;��	'�v4�4̞���I�&���h�Sx���Q������ܥ��j׍��\�7ʮ�BL�vO�8e�`�e����h����wT�@ �C����_�"�?f� �Y�Á��S|��ukɣ�E0m#�]���k-ځ��kZ�:��|ۻt*آ6��g�Sy=+�oD����v�HVķbI��WCjQ�v�־qa�Ihiaȁ-:�|�qaG�+-�<)���15�?�@�JV;t`m�L�k�m��# \�[o*�勤��q�^d�:r]C��j��S抟t�k2Q�O?�y�or��re_�@]~,�dɚ���)�)�>��.x?�.�}M\����%Ri}��Y�w����sn�x����|R�G�-5kQA��1Sϴ.��SHK���J�Ѝ�� �DBi�诃�|���V�{�M��Z'"��1-�3o�]����	��U����i���c��4�m�kvw��ׅ��z)w�\�3"3�2i�[�ba&�վ��zXrT6?�8B1�(���3c|�`��b\�kӅcN�Ҵ�Z�~��M(�Z3�Yb��	���r�}N�����p�%Gaz�]ò�PR� E��<��:���N����I��E���n s[� d7]Z~ �\m�e�ȝx^>t�V�C|�d�E��8)f��"OՉ�v�=?�&��\,���y�,Lv��l�w?�b�O��Λ���/���&1�!�7&�7�[���*�2'>G�+�(%N�ל#��7�D�aAÖ��Q�3X*�%+��M���.�����.��p��
R쑰�ăL�p��I�>�&�+�Gu2J-�mԱB���b7�8.<h��1q�v��,��&��A!� KA����Q�*l�� B�n�Kha�V�/�0���;�\�Q�n�u9o^�����HW~]��:9��f�z@�7ɉ�P�F���^���!����,�N��~ľ���盭�(D�0c�P�)@orެ��Y� ����5�^���y
�`A;-�A@x��F�М��r�y��L��e���-�RՈ2~�g�r� }�p�p�����8�����{��,w�1���U*�q۫8[�`����E��u�\R���6'���OV�<�-����.�Eo9�k �u����ő�n=�&�M�K��je��mJ�+q�tdy�SL�=��#�_z�q�>\B���P9���t��ӥ�CA1�%�m���_�q�n��I� �s��JA�3����m�$E�5.R5m�R�V�K�����N�۲2�O?܅	��e�&%F�н�k!+!��5.��Z��&wciW��,�f+�X�造fS�j�(f:�:�ۑ0F CP�cy⥸	����MC^?�����$i�r*GE��Z�$Y���a�E��/��t[n�zV-T&�rǈp���fn�V~դ5/� �V����H���[i�J_Iꌆ���摙-�]b�H :B�I�x���?��r�R]�9<כn�*H����������=���Sq̔!��UȈ�t��O9B�N�V���	�b��p;���9�x���h�_K��]v�7�2��/R7�L9|�`��`䓸0���P�.Ky�R�Vz����Ŷ�B�M]�.����1d�2��kL�d�z$o_��䀻l8�JG'��[agIVGp�C�B��/�l�^�F�:��� �J[�ln
��a��#����W�{J]-0͇�_]��e-w�ҙ5�=&�2���BHH'-�X�"~�j�EjV�����8��~fҦ�������
�9#���Ƚ����o�j��ƅ%{�9{ߣ`ܰѹ�r:.�j� �����q�g�!�����`�����rF�����P֙��BU���񌺭8>h�"�jG�<��bҚ��&�V����D�L � �I�SYlʱ�����x�)���۪+ߎE��4��a�lv���9��X�i/a�R��!"=�,��]D��9l�ށy�YT���~v�sQ1��߯s!�0�E������h5o���>��m@���&�Ǚ-�^F�9�e�<{�fjB�ӌ���[� A!Or%F�ba�4iq�(E�O\p�|dQ���d�Ra�r�pO�'�;���@<��en<<�`�E�8mS��֧�vp0���F�M���|u͌D]�S(�K{k�s�l�����c�X���>؟;c>� �Ύ;Ĝ.Ƀ�uo����=�֘2��p�����Zx�<��2z���A�5�M4pr�'�5���ϧ��qeu�-����G�����b�n���Lkպ���r{L��	\_>��R{�t+�R7�@;va�@N{�c�ʞ�R��2\��h1EfSJ�?^T\���	G۾��x�J��O�'��Y�c�}��5�L�����[���7��H���'�������8Pk.M����;�t^�ʯ��jڔ��J������X��)���s��~V��D-v��A1�w��i���V�7jN� +M�J�բ��Rw`�m�vA��Z�
gl�I�4q��֒t��M&�~�Vh�V�r�K�]� ?�3-T}����`�D���	���>B��п�1�����#��(����AQ/���c�������+k?�:�]}�X��s��γ�8�����D
&�#��z�) �P��� X%��ˈ��j`{���%���ًx��+��&��}�k쯊�&1��m-z��{/�}����i]�`�H��.kJz�-�<F�'1�Tv�I@e����Lm'9�+yS43H��$
��z�Dr���?X��5 >yzX�AӇ�|a����� I��洟���tN��K�d�aob���ހ��?y���A��t����#��_/�X	�Մ���ag�����B�&ڽ^v/���{̮u؛�Tu��Q�L>5�? � �����-�ʜ��T7�m�5��ǿT��	VX����J){Q#�
�t��P�y�RsQ0�,U�6�0���޵&_���}"����Tuh�⦭��|�"��ԕ��X��(�#���\�^�R�sI�m�^��-@R�(p6J6Y����K�e��&pA�X3u0=����4�.�h�Q��j�+&�������Mb
��t�ԥ`]C%m�vW�)t��.���G4C�Y��xf����:�MU�
���6���C��=6q^}DW@�,�4�l���x�Hc��8:T�]n�I�8Ϳ��	ñ8~5P�!z�S&��Fq-�]霴)B�=���M�G������B��t�Z����^A˓м�:���[o�ڨ��`�KQ���	aS��������6Uj�����6u%yS�}��>蓢F�94�xFc bI�
��[>s��t��n�Mc��"�S��Tά�%�⌋�u�1�qZ���`ͫ0Q��7�E��S��@C�/�L�h�Ќ�\w����7���3���T������.$����>l��bnQe�R!Yg�9K��/KFsT��Q�0M�0w4Pj���W�����@�g�縐m�jթU�}oE�$q~�`Cs�,�W���'�;�?`�>7t�S��V���u��r�-9��Ur�ˏ;�
�ހ&�.��#��9���	��ɀ���O��PG-Ϳ�	�5�'3�K"#A��8�(�t�.����Ҫv,ը�D�|�С��x�;]���B}"���%a�H�ek�c���^x�6Yo�$U�g��s|�*
|F+�kD�k�;��OOe�-�>3��zV������n-Jg�Ln-��{�$�k��{v��W��s�>�>��x�P�g�3o�]e5��G'P�F�����s� VT���~����Y1�>O�=L�ۯ���c�gs��ag���H�3���\� jyF���<��I���i$5'��"ʼ��ꪯ{��lz9�;'�:�BpC�w������C���F��]t��N�j�y879���O�S]Z�=3�NS�蕩�ɏ�Ҫ"�@�f󨄹������;#g��~i�(Ss��b����vט��]�W�6�e��q�X7�S-���8��Ȼ��(�7EG������w���Z���" ;��k������h-�] �z�h�6ѽ��ád��`鷺�߽�ݏ�y�B1p�A�[��*�9�D֠�Ȳ���hݐg��:��Ϧ���x�۳Y���J�>ݘ;\��q������� ����P���[Ϛ�g74�^ԛ�&L�w�)Ә���TR��T�`}��_T^�|���4Hj����fA��誢ռ����G��6�<�����3�l/R��/
�P��9'�4�,��I!�d�:JЂ����~�mJW���iwvh���=�,�X�7уUO�c�H�fj��|@����Z���9t�W:CO�����ui���7ɸ���}��|��d�Qz�?\�j�h�?��YDVu)e�g
�9�u*�b"��&�Y�N}r�f웝�^e���sd��n87̂/��W�Ϩ6.��vt��2�A�z�෇�t��6�'�:qd`��[Ʌ�#/�0��C��@�4n[��b��8�(���+�F��B ����ZB����<� ��\@�^�~Wry���ڰX.-���h]�%C��9�v�1� 
PP�A�[���V�cx�gY7b�n��?����JB@����J4��&+R��zLܿ'c��V�~����N��{�]W���,x9:�ʿ�⣼$	�r�WԢI�8"�#�]u��;�[�!;���Ӛ0�=>��yZ7��t��9�}�Ҿ٘���$ŧY�k -o�u�EX[�L�\��y๣��I��������/�R�=Ȱ2��Z�� oh���\���8M6#�|�z���h��_�}d{�ޚfq��RW�G7�V��PuG-b��Ah��ɴ����G������06����f���.�3n���-"�N!6J�%s� ��^�&�&έϞ�ƪ�hǐo�X�tlTc?�
ײ i%a�ګ�$8'��Fo�4��y���y����p�be��V���#����z�*@WZ�(ŎU ���̆��f���o�_��?���s���|���t��鼑@���G7��5��E~sO��q˂J�K����^��YYb���ʋ�
��)
}ӣtP)J#if��Fʍ7Ca�u�`H��	��N����x�M���	���F�2�oy�+v@ �24�?��[�E�r%$d�E��`Aj0�_�[��E���΋�{]G��)}MU��a#���q�)������2��� �E_���j�F)V���(��ρe{*�O*�:@����w6�}h�[�
 ���V�:.�.��`h 򕊽L�i�5�")k�b��f��t���Z�Z)�K��AH���J�tմ�'�dW+;=U�dr�r@��,Dd��������c�������''N[I� e9�/Մ�.���
2& *o`G��BLɄ���C`�&���=!�lbAL�o���s�IȲ7�DH��*��;��j�,�B'(5��}O/��t0���C!a
9�y�����i/����n�n`P��inj���F{���tE�]@վ�⻇�+4�F�]�;�cbW�A��_	�%r5������5jN�`5��}�[�ɭ^�	���A��c��3v��h%��n�vJȚ��;q�hQ����'H���a�ٓ�ض���iD�5��$ �H�l��K�J����Bu���Y�S�a�����,����s]�(@��/n��Ѿa��{�\�"�C�d^��"-k��y���F觕*` huQ ��z�wB�&����>��ЁC�B`��iO�P*�z�Ei91q�{�/J�sVh�$�J�J�M��-�rf� �x��L��j��+�iۋ? &��Q
�u�<53�f��RX�3�ꤋ5R;��4V��ʉF�+���K����/�)Ь�xwQ��o~�Km A�Aņ-^)T�C�R���7��s:!�>���G���N7�{�>AVHa�(��tREA��?x�/�6���ͣ"::_��'̤��ݱ��a������5S��Gs�}d��h��ץ������N${�j%�IlJr!�����q�iC�aҜ�m��Zkn��kM<�k�J�L>7��q�ʀ�m�$�)n9��d*'���>Α!aƶ�
�T̩�r��]�L�9�:�b��QN�����[�~V���(�u�H���-�����d��[��~Np� gް�& �������ϖ\$X�3�AC��<3 �jg�w�:xw<&��>���$}o���<�t֙8�jŅA��̄zW~Q��5�(�-�. ���Pֹ.�>4�P�P0[o~�NfTԶY3n^� �:5p�~2��y��l[�-�@�#y����fIۯ�@.�6oX��?��3�~�d�Mncɬ��(�+�D���D�����mѤ�-�A"������Ę�Wm�7��~��XX�%���.���R�1.�ӡ���dv:� �9�~ $W�XW�r�M�2R"1U�t<�����9��|��?�<��Ȑ�1�h��m==S.{�4��V��`ս�c�I���ٯ�����D��j���oL�׎у"+#�_<��!��ʟ��7�vo�[��jg^J�����u�N�@�A�穁�HB��m��$:���B�I�6�Yu��DM�Rs=02��@7�̽[�	�"��M&�������v.����h<i��I�a��]�
0z�@g[�˼�����T9�Sxs�	"O�Y�r$�H����w㪧�����K�{<jzq����"��R�1
�IpNn���3����@L�N3�׾� �Rus`ᣲ2���k�U+.Ύr�*!��|���+�t@�7��9l�gݤ�ESņ�{2�۟�y|�v����{�� �$�ؕL,�*S��E������ҡ;y�k����0��Z����!��=]�ڳM�J�Z�"��'O��C�[O��m�pfVF��cSv�M�-�QG׼RgWoW��F��:�/�ߩ�����`��[��]q�R=�-]��I�^�ّ�]\��n����4����^#X#���jlG�^��䃠��0 HV����-HBw.DGFm�K���v�۫7|���_$���!W�Z�/N��N	���H�"�&��@����.�!%i��������5&��I(ߓў��KwP����GO˱Ē�+i���c�GfȄ�����K��Ln�"�ڦ(�j�.5,�H�M�9���P�C9�?D/+Su�د�Ƌc���t�8�7?T�1�q�#�kt����#?Q��t����օ!IT���읷��J�ZX�E�D�,�S�� 6K����3FUtJX�Ǖ/�?{x�N�ug��sx;4*c�伵3`>�i���E�!lJ�_���0��a�p�9dǝ:q�bk:�[.��^�&�;߲=���?�?�*��n
/s�8��
��dN�;�d�]H,jj.����}���X�&�+fĳ�P�B}���S��2L�f������ �r1/i��ɖ�{\2�Q/ �y���Y]}�PsIL����o�R�?��R�t��.J�3g�@C��lx��0��Y�:�g�]����]�U���G��Zq�v���� ަA��hQ	�^A۸q�8�k�!fE�������plB���t��0Hcs��h�]J�M�*(u�c�2d�<����͢!XIhR؆��O+1յ��h����"X6X�sV"�J�I(����e��:O���B���1?���cxz ���Ep,�K�>��]����s�W�r�:��
���ɞ\Y��e )a#^�\m�P8���_G텚�����)�־c�K�p�j�
��޹;�e9�T�����:"�[uh���o4��p�iJ%�?=�΋���z碶|�'⊋�/Ai��յ��&8"Ɗp�6�N����c؎]�D��&�#�ü��	�aΞ$❫���7F~����Qr�W. �Z֑�~�q��k����FȫxFE$J�����m����aK�^��������<��`*2�E���"ug�܄O.Éi;���D@�<�2_��c��a��#���D�P��Zۄ���$�s_YD44g�gt�ֳGF���|�@�[|>nȦ��'�%l�Z�\Y�c�w���#,.�1n�m���̭7��3�3��{S&���Z]�1V���J�鹻,8ӵ���J�J2cJa���dc?��*hI�rY�+ROҚ�����:|}Q�ô�mK)͋M$Ġ����l0(���hgI7Q�dGeWL�W�l�T�{��V4�
�Ha��s�'���A�iUqZ�
���S��r�;�e"|�<4Sd����,`n�W_�GF�YaK���1J�&���Gk���p����� ����p��,B�! 
gBֆ���(o,u���?{qO.�\��'��rG���6��2"�D&��ȵ�b�b��TA��O`H�0�U�ƿ~z�Q�fUV=M�#j�fl$�"|9y�Tw�5D��'�/�P՞�:/t���t)��o�P�OSЁ��Z��~�����c��g�󰞦��U���p�B@��R�-�6�:c>ȍ\��[(�Y�y�P�S�2�vm����QB&���P��UG`���:����ȼfZ7����Y��!�mȊ���?Q���j���'P�m�%��GD"(�'���9S����>�H�o�^5ݕ��O����<ۿ�ÀyJ��g�������ʽ�g���6 �Gm�D��W#d�ұ�bՈ�C0�D&l�nh������	.��6+Q�M��5|M�nua˟��N�r��e�ˇrJn#_�W��!&�ZN���F	�潾���������5{T��|rʻ
�c=zP���o�QWI?��t�3�L�����̯R��L!�o���6�2N�ip�����Vx}��V��HY�����o�*#sr����tv;���\n|ㅏ!m�iibn[)z�>�+R4>@_����9S��i߫��nB`s�x�OQ��Sw�w��1��|O3����� :'7�2�g�2h������`�et�u$=y����� ��5�?*��r�;��o����^�� ҇M0���ٝb���~�΃ݗsK�Sh�cז	�� Bm��:B�sJ�fGq�����ez�҇���7��J�?���'��4r���L<=����ϷF���D>aw��^���9�/�خ�V6�/�՛V-�K�d���t�������j}�`jA�=]d�O�s���*+dKc�u�(�<��"�Y9R�l���E����nY_�c����5o�R�Oס\W�> 6�Ą��wm۝�g�>O2�E�-�˧�G����{���H�͍B
e�0�Mٗ��� $ź$�#'����!��.*�~��BfԲ�n%�����e�f��)�^F�KN�P2���s���\�����L/:l�����Y{km-	7�V��I��}�H��W�#�Wֽ�eF0�����H�K����q���D2��9��Z �/�Z����������T�F)8����2cm�.�K)*��&��e�%#��I7�z��� T5�N��k�g�q��qa�e�@+~	���U�.,	rӹ`zο�Fy׺���5V���c.�X�����n" �3��K������!���1$�����ѕ&�t���o_Y�Į4��[8ـ:�TQ!�L0��-�W��.x�H5��ߜ��G�J��"Ь����%���f�X�FB��#5��j��*�5m/�2
<�x���>�y���Ufa�'Dg�r*�Ĩ����Xz��x^S`���D�K��"=��sƪdJS`�r�pXB����K�G���6���+%F�to*5qf�t�/��P8�$��^�3B6f��c�6$�f�Ӳ�����M���M �������V�1�G]GC��?N?Ցf(j���y��vaF���!R�+F���)��N�n����^~�Ƥ̖�#�7t���f�K|-76	��0��0#<��\����<>�]?4ȍ)e<�p�0\u�����]��d���S"fe�����o,�?t�� Dur��p�+*� �-�2�t���zb<�`%�S-\�z\�^>�"���ųi,W�-������mS;���H0�;q �Zg��TA��AŁ9�A��鶻����ão���ŰP��t�����P�L0�!�R� �����Ĥ�q�'��Q�q�7�� fČ^?��&�0t������?%�(�F	�ˀ����^�B`t����7�}&1��*=��]/��� ���'q ����]�`j"P~%�x�?qO�YK��t)y-V����es�-���O���n��>�P�B�p|��%V�^��A�������Kj�g�$���&�g��q�86>�KZ�@�ɥ�Ìy��,
��Q�е�0M��Ɲx��L��t�W��w��Q<�JC���]���I� z�í^�rK��R<��X����靖a��}�\m�xHAb�&h�,�P����6���Ry�}��'-C F��k�e���^���D�3'��ݔ�c�CK����LP��֑��8�[��x]���W��NpS/��AǗf2̓3�{<�z�X?�߃E2n�xG���{�qب��taP���̞��&���Zb��	k�M����t�=*��5TB� �֫D���Mm��Ԍ�/;|�����{
(3�)@��p��;W���j ��U�iVk�u���2��0�ڹ�R�7#$��2������d�}���ȳ;�6��1��� �j����"VXڽ�_��G y�R��ۣ2����?Z<;��c[4�*�ga����[9������#a�5�P�+N���:$�c�]fur���k���p���=4ƶ����1�V1̛Li�:N��c�n���
�uEH|^�!󿶄���x�ٺ�n7^ׄLͫY3�g��S�V�q�a��h��fG�2�T�	��>�������χ��V S͐��������V���mE�i+������F_��
��������|��o�i�h5����0��g��r1R:<j��WZ�@+�o�T�{�Iq�~��f4�#���Fc��YY�v�
*%�3"_8��TU�e��q�:��w�� ���A������u�{��x�Us���PR�/G��g�t���[�4Y��v3�� �@�'�~;FMC ��`�`�j+`�]�N��M�0O�&݂��И���W�.���(��ʁ/I ����_��6�c^���	��1.I�\-��J���R�����i�-ԂQRI۬-Fzh�B���1��R��{>��'���S�����5]���S^�ㄦ��7��=�0�e��ѵ�����ZH�����(d�gI��K`�R'�GE�?�>���>0!6�ay�	���A�w ��Our�T'��me� �1-2���������������KAA�al�a`>r�{L������������"l8KmI�y�6�'ډh�gc�L�`c(���őߤ��t�gpa������o���X�}�*E�<�W7^���ǰ�[o�X�:��&9!oDB��1�