��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n������E�u��#F�R{��:�b;xj���k�8������Ԟ��6���@�T9N_m��K�K֔��~4�YV,3��芦��v� ��?̚��}[C:f��$r_�^����M������كN�ڷ޸S�s�Fߵ�<õ�����s9��]#��o��Y���]�+f%5�n�n��Y�C~8ƍ���|���g&��sD2�r� R*-J���O?A��n#��\�[��T�lv���eA�.���~����f�ٖB��_�����.���I}F�C��Jٷ=��VC"?�Bo]���*��;��������dPG��On�f�
ER�Rn	��LÝ���ݬ�&)咽Y~ˍ���1AZ��ܚ��&�'�Ɲ��%�x�3�"J�z�)�[H��������Nx����:ZO�K8�]G*�o ��<Λ0���َ5���[#�=���kΨ��mJ��iN���	8j ����:��r��dV���Q������sf���%�\NxO:��ri�aY�����<��Cu���@�f�v&�F��Yd�y�m�s�rɔ�yYl�͛�{�C����n:'�[�wŧ�)4p�K�Q��O8p�r_�;��ˉ���V�do����G2�+�g��TS˞�+�l�O�d�&�y'��!xpU� t��E&��y��|=Zg����� ��1�Z�2��R���*6��4��t�v]��蠝�돹�g�{C�I�$��;Bp����	G!i�QX
o�|�LZM�8��N)7�����l�f�/pI'D�V�p��aI-���g��z���<3Oj�'B��N"ߵ|o�[�t���O�m�*tD��.�Jz��~y)��&CLM#U��6d�#@�����i��n�FU=aN�va�h\�v���q���/T�^t����a!ݪ��Q����4� ���2K/ln�A�T�E|�hW�y���Bhy ���`!<���q�s.�T�� �X�؞1P����k����.Olx�+�w�Nܢ�PYH�
�[���n��=8�z��y�V_�$0��o_Ç�"p8'�m���bi����w�Ƕ�m�s&3��V�u$���xF�癤�g���g Na%�Q(h}ob�V,ђ���^�-�ݐ��Q#��0��m��n�?9�׉0��ECL�͔m��n��V�W����c���a��B���
��T,�ڍ�z�J����E��]�M���3���mS�ɻ���.��ܷ���,����n�$f�]�q�I�3�5
&R��M�%]�Qx;ٔD����l��$�^��Nm�&FΖ��֌$P��2Pӌ[��mb�Y�bD׭h�Kh�^0�C�*$�0��d������������f8�"��/��b���Ü��8��4����EWk��@�;���J�z��ŝ�_�siw](�^���l���n�y2
�w9�Vwg^��ίf�����,��`(�������i�݆C6�:=C��D�:��?H?mr������,� �(��AJ��FG�.�����Nٝ�4����RZ�:H&�ش���&x/��:�k	ϢS�PI���e�q�X_zY�ٌ8(��}8�Tόg�[��t�%49+�¶HD��ʶ?RCb��?�TI�U��vlt�_t�b�Ǒș�9@Z��r�^yʫ��{e<[���u���uX>���*�Z���V���S�S�=8�x�_�>M_.�:A�E.�	٧�c��?�p���5��p�+">�Y�eA�\s��c�Y��4���敾�X0$��h.�"�쬀�kAJm��9���54h��#�A$I{Kf�ݹa��kQ^euV��?E:',a!:�V���r3xsȳ�>U��|��l�"(T�J�wy#�wj��_nR�[�Z�?]��C���k�v5����@�)��5�:7e�n�?��똀0���J�� �.+�"���.�_��Ka��-��`�`��c�m�Z)DK�9���E�\'�L�2��/�t�j�	���A��Q�2���LHXWx�P�f�_#B�O�T,|n�>BN!�gk��e0��R��'HKP�xz �j��˛��ؖ|��%6����/2l;���~��J`F�f,5�z���Y	��&1���Z�W�/Vo��۰�D���D��V��ɽ^_��m�ן� �
i��4�$�1�f+�׾��j�.o�N�S٢nQқo���N�5a���䠹h�ʝ�"���6�V3��pxJ��Q�u�rT;�.RX�}�Y�j�P�ڔL[��A:nNx�p8��o���0��Q���!���bH�܇R�ݑH�\�@�Q���LB���H�m���8�����������2G�3h�3�*�Z�if`��b3{�����yF������h�_�<ʔIC��`�-,���;�Q+��RJef>@�
�Dk����^D-��и�A�h�ثI���g��b���ʀbe�e�!HR��k������sn�%��`�����o�n��K�sz9 �a&)��f�=����&���fYH�{�Kb
e��SH��){�A {�<9���Ӡ���a�2bS�"x��b����Y�7]E��7��4��Z�Y� U>+ʠ����oZ;����Ĉ�hA4yD��X} +2�;�͔d��+��(���|j�p@�OI�^?_�2!��i`���|��Q�Z5�P���w��F�.L�9e���n��#�ˍu8����]������l9~�����f���c�޹88�o7A�I|2��U65���H�g�*��R��D�_�2 � �!�XR�t�>e��p�񛟚��?��b�s�v�/v���x��W���ƥ�ɦ�M�i�L����J[�h�9j_a����ni�e�9.;���2�������h���o��LL�<� ��D�/a�W ���)�N`�a�Y9/YH�yŉ�mI�?#��i���;�z�]?�|���P]/�
r�D�%��#����V�����ێ��n�W)��V�H&�h�U��^4'�9;�=y�B��?�߿'Ip4�cC�dm���]p��$�y�3��0�}� �܄�����o+�W�1	�W6U:7l7���n�l:�U��K�lAD�t������퀔�M�Q� Z��(���,�(u_V��Cd�WX��BsR^�B)�'���gG����� ��X�JN��AܠRM�W���q1��AP�.n6��byf�P�r�K��og� 0W55�-�Hsw��bR�7�e>�������SR����?�S����e!����E=BJ� �ND5|kB(}u�	�PNsYL�g���&�|�jS�ߞy&ʫ1I���N�a��%�[��tiC5p������-�����s�����E�C�e���^����X��IƝ�(����]_���?�H`�L�H�9	~�2�A�jw�7�]�k��)��){���Xs��{�x.0�Y ���<��
�.U�Ǚ����e8o6�/�l�C��[m��G	��|?�`��O�p�P�66*�2B���g������2l��sꕷ�"�N��Q�ʊ����o�%�aF����24*��2_)G��8ty��=���0��1aG<��/2j� �!ѩ�!���LoZ7iawKo�"��D��*�E&�x�%R0	^0��=Nڪ+(�����k��2������b�h��q��Y��>,`ŀ��;{�buA
�u��@��J��y�a!��f���XF�Y�\? �M�sa��w%~�ܴaU�-%O��|gwv4<*�:��q5u_�n�VZus_�?0,��? qXc�.�M{AXy'�L�@L�y�^յ@)O(�0�I�D��Y��2�$�iD���k��T SG�I`�̂���hΌK�!�V����p�Q�Ki���o2�������F���7��J4:F�]���H���Ӌ^oj��s�F�?u��9���dY���c��'��W)B?=K�L��ByďH�n,~�Km~E<��*�1�����4R�{T�/7
p���� ��S~���g�����9s���ҽ��fg�ҟ��Ť��&0��Ѳ6֒�9Ӌ��6�S��$a�}H��eȗ�gř���>�[�QV�q�R �g��	Șz�Y�ᥗq����/��A��m�Ր� �֮f�����>��#��.tm�}�r��i�\��e�a��"1<�3������"�K~F