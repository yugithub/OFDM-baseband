��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#�����~H�����pl�Um�v:��L��Q����;�~��?U�b����1�w���`� �2����:S���Bq��6w*��v����m��<�,E�H����,�b�M��1>k�^��&�SV%�n��b77� ��������m?��8��O�07�����v����-��Z�h�-"�f����v�Lk��em.������~A+@$���V�����z�K�Ex�;Q�2���Ij0�P~�ZR[�J�>��As6�a�!9�D0��c7�w�䔋G���ITwߦ�8k��i\˧�Ǚ��3|�İ^?��g!��
&�GCW��'W=+4=i�;(Eq��;�1!�jE�O�UX:k�9�M���L�Y sƑ�~%�{ݽz�}�Cz'ט���i�6�W���H�O��/�ӧR��k|����a�rT3�Gqc�T�T�Kq�bG��E*]�)���-R�����TR�z�a�Ћk�qum	�"v��<�E+w�L7i_��vB���=H�L�(�Yk�j����>`�g��ݖsJ����"Q���m&���P))!@8O�h���Q��(x]��u�=�� ;L}��9��3h �v�6	�?��B9y�?�x׍��Db�n�x٫FY>Sz�8��:6&�~�k6y.���Uָg�$��7C_V0O��"��l��{Ez�q��dB�H9��k��.5�^Θ���3t��BP�|�:b;eN$��/q��T`K�,fm��Tl�^�� �ו{���;N2�|=��w��ͷ��yA��!gs�*��V��I&u7.]�y�ꢢ�"{���'*���#�_3�����^Y�E'H�i">&h=s�� P#'N1@C�������7���k�d��c��Û�i+Jr3s�j����l  �DmW� ��X_(M��o<�4p�j�����e��Q��]�lG̵:ۯ��3d�Lcf��3���EC��*�Xo��}�C��2��\/�f=Z��wHۑt�b!>3ukeSDe;e��0+�|������F��y�-^9�o�h>i�0{� �����W�,�L�&�_�о��{���+�}.z]-�����9���kg��
O����8ì���%iG~��U����5��K��$�<*��XR����'�L8�h�����s��՗�J�W�-��5�����
�Ee��*���+b�ڑU�܊�@�躬���m'#B �R7�pr�P�a��^X�Z'�Ci����'5�~(k�f��5�wl��6�(6�{=�al�U�e��y V�-]�x��������i��t��%�o�P�Zw�pes��q($`QM:-���ƽch[��r��/�Ѓ�aT�`K�`~з�VD�ءJ��*Qu��A�(a��0	{g3�W��7�˸��b�,.|#X�ԝl߹1R��yR�Z�g�'���H�+g�*��1j�|A@�CR�Q$H���<���|�$� �	緋�6-�_�_�k_�۱[�v򈄈pP("q�P�րJ��c
�9�(��̦fU'�y�N����1��芹ġ\'e�k����GE� �XI���폟�B5yWHXF��HCY�r�?��/ل�c���߃�B���X��R����.T"%�FIk8���W���tC��S�B��ܣD������x��䁘F����rS^j׍ ���f�����د߂��;
�+y�KзV��$WPK@�b�,?o�p�1tcŚ��*\6��Sr^^�=����ew�?b�r�.����Y{Si�?fV���˨�@�H��ZAh:KF����e�Gvo^{��$"��8����Y��@�ᠵ����Nh��-��Ϟ!L�$�9����
d�����Ⱦ1��O�PY/[�~H��"j��g�d����'(��]p��sj�`F�ŷ�5�jY����;�#h
��]~�`]�zH-��a����g��\�%FW��C3[������|���I�Z�	�W�z�.�͔ȁ�(�-^�TBѧ���#�6�����8��N���)Ւ*�wbRt+�y�8����{[�"'�� ��#�����
";ߧކw�l�|��.�/����kH���"��n�)��DZ74K����qixi�΢_S�@P�pܢO=�ϭ��o��Mx�41CK��2��h-�7�~��М������� v�\΂$H'^{���p&5�]ȟ�<�|�~�ʴ{4����5G�^u3��#�#��c'���Ј1����~-m�֧�KTy~��{�o1��l�� Λ��	��͑ϱ���v?�6C�ғ��IS�cV����U��'�aR�����l��X(G
��c��x�Kĝ �R
{q�x� aڊ�hȏ\���^]�� ���&�+�v��������ͱ3��C�k���ￛ��4���i��*/ Tڕ��Ot�o���ԁ�-�eH�q��a�[j��F�æ�ڝ��i~�jʲN�weJ!���,�W8�%I�+X�mJTV]�nZ��\^��ZZ5�x�{��`�rtdRN���� Ț*AV��ő�j�bѸ�0�Z:�:+!�:۳v�Q�IĬ;����~�f�H�����tP�Z�Cr��L�'%"���^2�|��h��8�愘v$⼴�X�6+�a)!E� ��Sj�+�=��F~.k^�体�:�zF����]�e%x�g^ܼx�9�
�ZX�B�V9w�r��]-G|Ŏ\��:i�~�Uڢ���REk����nf�T���a-~+\Gt�Z���6\U�j�";�XV�DX4z�i�U&>,�G+ⵆڄz�Er-�� 0�e
���`RL�j�
�M��7%�F&��T��`%�6�oU�ɽ9��g�x�q��؉'��N�Q�65Mm�8g�y��w�?Ȁ=Ƌw���7A52��(�)�qdk=z9��,��c4�3�g�˄uH?�������I0!�����c7�Ki�l�����)n��2��F��z�̎G'�琼�m��7��-�v�7��4�\�T�M��?���>�4Q��z�gb��=ܽ}WG�_HI'�LD�)"����C���{ӊ�W�B�����a�p7���Q���s�h�b�+s�up��'^��6���
�w��8��-�Au̬~8�H�T\E�]}MO�4�~��	�P��&��a������22"?��E%�Y�V^â��.�xT�A�`�0U�GOj١�w��i(Q�'�	d��/��Y���P�+P0&�	���oe=�MQd�۸ޯp���:��$`狯���}x�S�F}�21g!�i2��N.�� ���*�^��$X֌=��a����b�)�,�z��8~T�W8$�5o6�2q%�<���=b��-	�.�����Ŕ�zO�	���7u��V�KbL��`���u1�Ð�8���Yg��B(�=em�ή둶���D�r8[��cb�7l��Ö����Ǡ	����Nl�x�&�-66Z�J7��*�A�3e����9��Q��:QJ�]��	��c��Y��/����%i��ˠF�7S�����v��_ʱ������\�B�]rJb��x�ݢ݁��f���^�~rfk�rD��ڏ֎�Ɔ��N��.{��睺�b?��Y�ݪAe.�Wd�jђ����n��H�[�;nFd���ތ:).��&��l���vp�B�pW.#�Mף~��rCI"�Q�G@�M��`�\"E�l�����m��H%��@��T���{Jn��ޕ`� ��9��nsH֚U
e��.Q�I�F�e�n�徖��M�ܓ��QY`,Mw��K#�:s'X��s%=DB����r�͑�Gx�a��Ҽ'������A�:�Pt�O;�uH�&���$HQ�f�r��ǉl���]z���h,j�����5�P㝽111�Pq����˚��嫺�hz�k�}�`x]���b(�ILjЦ1�ߑh�������+��d ���8���jt@�@�UP��^(uG���Lv-ءf�+X$]t�`��jD�r8��D垺�{-3�}��p�P1�"�~��:���]¢��̇�v�ܳ�	���,����~�r���
�_�皝���[We�T�ј5-�)���y��W��1�:��NF
sё���3�"��//[�Oqf��%d�r�^'C��0�g��rɎ�e�P�2�?T`	��c�j��L�N�ݾ���-�RP�~�i~#M�B���&�}c\�z:7�lv������sDJ���x���T)���q?�P��EJC����������1oD$��|o�߂��J=h0�?T�,\%-�6\�Ɠ�^ّ*� �T��D*F�ћ�)H�X�۔��KX�C�7�"P�0�_�"��bM�'nj4X�G!��i(<���ۘ��ʇ ��(�8+����@7w�t��LJ�HEl�f����4�Ժ����4ɦdzp2;9�FT�Jt�����6TȨ�s�s�Z��8*`����sc�̬;j9Ǐ,lXr}4䍜�-�����%����[l����Y���6��a�{��q�E�ӉjWR)^Y��x�p�4D�dvd׍��"��%��y���n�ג!u��1V𙸿�A|�	T�Ow���Ә.M�6b����@��������<��]�￱l�X,v(�0�d��Ak�	m�b���n��Da��M���Xkn���^�T;3�E�6��Q��Uo�, ��O�'5I���p� ̷�cF��)0=�z���lm��?<���pbU��.���h�r�d��L����A/lg�/�;d�'@y��:Z�����0�p!�b?Ԭ�Co�cΰYᄖ��:ku2��'�N �������c�����J��w=���q�l��I�<���P=<��x1_�v��F4��XLo] ��*�B�n`�ˤ�9�38�� E>`B�����$2v�jk�Bk
ܥ�Z�h��klU�������m��RR���!���:H����gL-U ��������j�)�w�dɨ���Ĵ�{CB��y�����{<��k�]�6"3�z�D�<0Hu�羼�R��-�c��nOq,�KĊ�|F�9�I�m���әue�M�r����\�V|;8�7�s6A�o�7s���hf�����i��=���{gZW�6������e��n��y���x���� ��?�͓Q�R�V�����by|vz�,��z�s�q���Ftr�.���l6�=��*�0Q�p+�s�]v.���e�[�c�*}��03�0.<�o۷�}����:����#�A{�\�x�k|k>��>8}�s�p�P'�y���5E�9_��2o����~��w�ϧ�-ѺýK�`�w5/{)$�Ѱ�_J憖B�.����]r�aauG�T��΋O�M�-M�W׊}o�kŔ�}��R��ni��6nҪ`��u�����_r�L�g������~�r<�jޜ��.�i1ʼFä�O=�N��s�Et����/� ���;
�R��}A�-l�з�
����}rg7�F��Ҿ
��65��g�^�х�=����y��'�o��DK��� ��2mS�[2����Q��]�][����>i�u��H��Nb�����Z�"6��������ܦ��ж�g8���9��b��-.�DM�,��N4����v8�+�q<�U~o��s���Qp��`����qpQ?�O�[}�j!�5��\,Z��tD�cC����K�����������!�f�7I�@�'\IPX+��B*Q#	��u(#�Jj�laP�<i�2�w$���U
���&��
fb���5������X�d[��i���*���.F������V�k�}Y�b�����[b��:7�t�ԧj�y����Ho�<��%R ���)1�8п*�M���IGF�b�F��}�K�_���E^>�����;/,)9��Z�1+�o��4�Hh����,���(JSZ�oL��vQ5��G�����r�"�}I�'b�$�����g&��� �MJv��#n�ゔyA/��+�]�*�e��#>Hl��̞�S�\)��%~��/V�K����ݖ�	=(#�y���]�7�eǎGNоR�ǭ��v 7S{��~�)�nF��i��huuD����Zk�.)�D�AV{P7�U�a���]p����M�6]:6�Sm�uv	�K���:�qݫ�,�K�uKS�m�hGW, 2��7�r�0�)�?B�E���ZddXz�%�Nz�B��4���VC6����9$P+�8N�3M�,E~����p�	#��o}�y�����fѱ��p�U�� �a��+���~���olq�!~�E^$�0�',��' ��m2ar�	v�	�ퟆ&�8>X:��g#�8���;�H�ty��f{��ʉ��FC)���3*
�#Í�"��� �va�g&+��p�h�_}?	`+��("S4��H�fɱ�.p&LM�c{t��/(�A*�5�06��3�@�§�ٯ"Ն@�yk?�{L�ƴ��@){��WZh���eo�T�W��_���.��Q�E}ܴ/����\��M_h�GBa;PR�ci����~���.}�GL�5����G�4ؖ�5�m��5����*}�`)K�O@��o��#��k�3��7G?���`r����?�S� ?�,'��%��2��CV�����(����do�Ƿ#�l|��ķ/d'9�a*����/�P'؀�Ź��O�.2$sQ���t��BQZ	Q���O4Tqb��[��r��UU�c �����Ñ���YM鍭@l�����	Ŵ�6 Q-�@E#�ث��Ľ�t��/�����h��HD�K�-Rq�dhb0�>�U��uTBnܱ��9.�a��V�>L����:����Q*^���/�^E�bT� ^0��I�r�2u9'����'B!OB��M����C�*��ى�Ŧm���?8�r�ۉ���W��Z�v8�O'�r��dg�S�<�C$��̡〘������:861�@�
��L�ݓr&Ц���!�ʈ砟]��GG�J�H�q4���j�f��4y3b����d~�Ɖ��=���6����q��1��m�qi�2}3��(p3�w_$e��9�;�����Iw�ZM��5�<��K�!��o�EeNC�.`{�*�5>���ĸ����x����/�Tt�(�b=�lH	�� )8k��	wd�p��F|��׹�Eh��`ߌd�%F��.Oɋ�Ke��x�����g:zkO ��_+���X����Dr����y͊f����k��Q�F�14�s$;�?��6�A������n��`�@5>u�ҩ˅�j��}����)��z	G	�V��S�5�~�Q�(b<vo�Fi-���3��b���B�x+�@Т����ؖ�nGca���2�*(�@r���i0�=B�&�aEe���|#�Qϝ��a�}��9]:z��HӨ��U����0��W(�G���!�  DZ,3_m�V�Lk��}�R$QJ��r<I�����u��0�d�Y�.���Ө\1سQ����9E�I ���*���5�U?�o���<�ԝ1]z8���uAV]BA{�_��wz��&�L}�X��S�}�Hg֎k|ܻR�5'c������0{��͌���/~����Q)	���FT����D��R��?4-Bs�!!�Q�cGy������w�E���>��A��%	C�:x��ڏ�mv��"�%�[��{Q0m!W��|���I0|��2n�h�� N��k#Mlr�A��_ERT���5 ��f�BqP�B��/�ۛ��4�Ċ��XNX�a?�1(�W�$,-��!9a�4�W�:3�E�	���X���:�uY�f�%�H��1$q5��jy��,u��zb5@=�*<v�\ҍc?����h9}z��������A�3Qx��bK �c�vb�	�������xb���Q�[�R
�:���V3���Ɩ��`H�Q��$���m�+")%�BCh8�!V��6\;�si]X����������gͰM=X'�I�?u�s��.�V>��S��4���&3k�S /Ě!`�"��Ӹȕ���(8�rO�K b9N�pQ֠�p�2(J{�/�O�!;��j �;��$��y�i`�᡻6�q�x����F���7{����G�5��s��@eâr!���:w�P<�#�ch�;!��wg��$�T��$"
_�
�.�;E��i�|����O?h��Fi5������|��-���t@�W^\�0���s�,�H��2��u�I0��I6�eW�2���W�2N��׈o�e�Bڼ{"-n4 �'�6%BD�C��ϖ�z�Ĵ��|!�z�"��ͦ:ǿ����+���Q������XPS�6\�[Ml�wI���P���!���z󰺟R��\�|X�����3#=����=�,�!sO��w����ΰv�V�nt�$�82��N?u��ʕZ�?�H�k�NA	M���ݾ�� ��!��@G�p�#��
�ȳ(FԹ � ��B��B�|��l̗kl�]<'i53����!3栗6�k��݀ϓfW"ͮ�O���Lh9tE}�A�`c�k6�6�륒��ř�e������!��*$������3)����ꦇ4(�R?�c(W/��N�f	�hKl�� )f�#
fK/�֞L**w�Z�3�P��s��&�8d;]�SO��D�-Q ��ؐ\��[�z�'�<���*���R��_V	��	i	�$�"gq-���*��9�����S�Wd+_��u���>w��$>�8 a�%�0Ǝƍ��FFw�\]�XN۝�b㚽��eU`��>k"����=G�D�d�Hw�Ʌ>"dɂ$��ݠ�D����^vğc�w��v���{�� ��ڴ�&O��ڥ@�#���@Û��@��o��eJ�:�L��Q+�]�:������F9ln ���-g&z&�#�ഉ�I��|�u��|G�ѓ=���w�(yc�0�>�~M'�:� 3I	���)M��H})��~��S�&���1�
6#��o{� ܼ5��l�%0!�k|C�a[W|�>�I-a�G�h'���V�M��%9�s�u�7���=n	����늌�����y�l���FWS��h��Τ�>U�LC�,:��8���a�(���,do,�:R~~�(�� p��¼����丆X�	I7�^^u	��<����t����O	�p�!v<7��eEܲ0�􆢔d�MZC���x����Hj��w����vj=����J 9x#� ׿�����?3���/PӢ�l�FM1[�tlm{�U��8K��`Y)w���NSe�?�o
�N���E��#xZ6� ��0?ʪY�Ӓ�j|�.��@ԛ|�aA��U �ř��*�(s��'F��7��l�o�R]?*�g+�ۦl�ۛ�������#�'"��Ϫ�l:��9���{�b:����P��W��JR���HoM�C��]��i<>����oS,��R`w�n�J�CET��]{�/���A�����-��:��^������3ld����l�H�e�ge�%sp�ժNhƑ"a����!eK\^������ɟo�{|���9M(�CR�oO�##\�U�>d���&->�%�!9����,*c�Tq�n�#Xv�����B��L�	h��n�K�Xv�McC��~d%�U�'*��ey;���ќ.��#�T{���7P�Md��Lo��!Q](��R!&T�c�c���#l���A�w?z��c����>�X�}?��3A�.��X�a>舤_���ہ�H�Q:Z3_@#�W2l�@�����X>��Fh8�s)4�`�c|e!�I���9��|�'}�Qt�v:2t~�t�z��B���P�m��)#��7�`���U6��.�r���d6o��c��/x}�♑�� �UX��b��6���[��ՄI|ɵFK��.�������s�����m٢wJ�?t���ܔ��ܞ�y���㑜�NW��*? y���H��H�0���Č}Ng�ϴ�i;o���X(�ol�I��a�0���"EDEs���h*o�W������s�-k/!r�;FY��qA��2;�����O��i�S�¢�Y���w��`�~�[�R��0dYAj��mݮ����fJdk3�r��i��4���^17OFZ&���מ�R6�稚Lj������Q���e�p�+�}���ߎK���<ٞ �P�� Ĉ���y[��0�a�gh���ؿ��8�M���͖���\t"8H�Z/�ӣ*?_�)���k3:��>2���Ʌ��GFCM� F&}��>������ղl��E�d4|ح�?�B��8o��@�]��){�NP�XK+��DTכ���-,_�t�R��a���Ֆ�4ma&���u_���C��h"�!����Y&s&�U0]W���a�m}V����d��n�}#=���'�P��%7r"v�UWF3�%�9\�Xa��pb�^�"7f=�l�mm��PZj�m$Z���9�'�C�����+}�{F�}���Q�BXW8&Йb̹��	E�?��1�[�����=߄�(������$-�NU�����a�hPD�=�+�v���J��G�	�x�rS���L��{���͓�X��C���5�h�ְ$'OM׾wL`�W8���U=�ؕb�]����p֬�����l/Yx�}��Ji��Y�"N�#e8h%U��9�>�|��;�M1ڄ����_�m���4��D�A��.�N|3���_�;��nA��^ާ�mЭ(�j'o�m2������0O�����a�T��_���Z����^��K���N�&�l�5Z�v�2S@k�_�����'^ڈۨ��p�
���lmm��;	9��L���o�[�D�7��G���a1�R�[;������Gd]�^R�>����gB�y�� S�/�G��8��j�7>!�.�����^\��m�^,{�1�.לu8d���ۗ��a"�"��r]U*NᲮ�[q�^�,���d���'=��23����Ut�P	m���v5�!��廯� ���(��WAK���O@��6��JJ�$�KQt}���U�[q�b/�{�~ŏD�y�6�G�����,�6��o�x`J>�,�F 2/�H��:��2uu��V��h˃ ��Y
�,�Q,�ߴ������b	���8]N��^l�D,J>ޮFx��w'|�M�i@���'�-MAm�5_�ƬH�`�5���.��$��/�6���$�S��8(��RF��+���6h��Ĳ��]T/rx0��Lǖ4��ɳ�$��!2�sMU��0��(P^hgX>􇕯�(����3=��q����}ۑ�VX%],�S�%�w�1-�P�Z-�*�@	��cΟ_�����&���:�1��Bw]P��kfѵjV��$[�pV�=��B���=h���2,�s�Ħ���^Z�,�Ƚ� 9͏��5=��y��gx�~��'$�&G�X���	ףg�"[���_H^?��]@��J�o�d
IҵM��l����i��O>yQ�q\~�ze����)��=��Bx�ʽ�[�6�ܸ�!`�3-؋���l�����Ѫ0���Uœ��Mvw�脢{�uL|�:�[^U�I^��UU}Y�p�OE[��(���
!u̸U�����V6���܍�;bQ���CeϰT$ �6
��S�d[;�8�:3k{�O	��$ǀ�5T+4��]����$4O��c8|�����ylҁNζՇ�$ۖ �*�Г�.��%���������7:"-�MX.A�<˷�,B��Cԝ[Ưԗ���c�в���2y���vl֘��4y8��V�΄�h���L���ݝER�>�[��΋˳v�MEu�0�#%��7�?2�4���V��m-�w���=N�k�٬\̙����X'f�֜1�������m��m�-��v�g����c&��4␔[U�Y>��)U�$/A�dr(�:h>ߐ�O�
t��ʿ���B��N�.?��M�;m���M7,� `?w/������V�}����U��]���<���^-�X[.�k}��28�
�s�g��>	�B���a��vH�I���ݐ�1	]g�(d���0p,tQe[�0�
ʽI�cH�j���^���;2��;&���ky�_���&aX2�^r+�Tp�6�\�y���=_��,fe:�t�f%���2���DR��{a5�'a �jmB��q��H�������1Ӎ�ņAD"�l�@�B�����-KbI*j2�tn=�l}�(/4Z��ľ1�NÕ�E�* d��&��;Rj�ݡC�=�00�dq݇�Q�����*�8��G�ĒI�ba}�qZv�P�5��yHѡ]* T�z�>�G�Z��|?�s8� �dGv�y5���گb�QМ�����^,IC@�ui!�@M�����ԅ���/�*U*�2��s���3-�����T�q~�&�O�\Cْ�y:v��(��Z�4X���Gg�[��b+���s#K`n��C@�{=&���=���!	���$�QP��{�7��+Z]eFY�ե���)��-�O�	�6K���tQ��%��|��ק iSص�I[8>�f�s����>��/�
��u���mT��a��F-�T�F܇�s%m��"��c|��3P�"�œX�xR�7��<^%��ϸ�]��]P0Ԉ!���������m ���?=a4܎J��<��@fto�Է#��F85�y���";J��0G�y�~�M[:���}�tL�V�V�s�F�ۆ���~3>��s��uI������M�WF��T����s�ʕ��up��ݬ�,���1;W�9��b1ZܙGK'��eΜ�9��4��-�X��Z#������%:Ռ�c���J�vl�S�vr���fA0�jp��z����*�>�U/�T�#Q�3�����J��4�TI|�N�>D,�Ӄ씁��Ê�o ��}B_UR�>����=�_��D�HW#y]1O'1H��k�R����Eى�m!2���J5�6�� �~����R!>�B�9�e���̿3lï?���)�v��(; �6y9�"�{���G9�v�|���/`�����H�ҕ!K��o	&�)�-�
r�ɑ�����A�~�M^����y��|C�U���K.n|��6�������"G�T��5����S0�P�%�5�cV�Ɓf�AWC����GvGl"Rȏ&���a�����@��T�+��ܯғ�F"��`�k7��ǆ%��/�GO��$g����Lx�y��b���R&�(m�3���Mx�`��t��c(���.�6Ht�!�_܍
�0���� ����GaD��<n�:�O��aa'z*{d�]/��Vz4�@2;�9:��L�֗ZӇŜ�_�;�����'C�U���r�1e���"�L���"gV{~տ��̰��u��^|�<�0 �oRt�k��ֈ�{�Vt���=����@��o)�wA�η�M��	u���6�����\/`����a  �ƽ���E�mB'$��cF�ߧ+7a1L/�ԕ��pL7�Y*z�a�Ӊ��h!OKN�}��Kȅ9�Mu��:t8[�ZR�fǉ0���� ^��o�P��<h�l����\X��$� �t����80����2�Gqo�o�JJ�Z#I��R�M���R��#ǻ��AG�ă�(�KF�o��@�Nf2��Y�&D��� @9��2]�D��vBZ'��Ǡ��4H�d�c�u��_��0��Tn<:Y���f<Xd��?�뀲��W�܅G����b��kY�찗%�ő{�%���U�}�I|�+4�g�P����^]���H'���y>���d�E%.E���{�`�� ���#��� p��/�^��ב��`F��7٬����T���!g��^k�mt��&�i�z��u�����-Rx˫�8댣Z�`�>���\���3�4���Lē�+N���?+1-w�� 	igZ
γ� ٞ���.2���l��ж�i�$�����5=���r���"="<�Z��Bf��Ş���u��x�ǔ���[W-���7o
u����̰���\��,3��}A!s����-��XI���zu��wxf��SCMQͺ�"�G˘�����	���=$6
��U��&����ՎG���x���pou�^�Ͳ�ҰBM��V�i�f�������l�4]�"SG�	��)^�x�#��t�8� B)�];�|�'*V)-�2MN�o..��u\�M2�xI]x�Xx���3g�E��2���I�4?��6�&r��ƈ��#�t�0�k�>�Gv{W�-�/X��d�޽AAv6������XO�'<�h{@L�؃�*(���=f��H3�� Ty>���+{:Zkoaq��N��>�XP5d>������c;���
��_���_W�;ê�m��[ڛGgb��
/�[�H��8��箿��":�Ez����n���T�xH�>N^m |CR.@�`��:v�m}^�Y]��f[ݥ��=u]�/ײq�Fz1�5M�у�4�ӑ��f1��V䉗W�k�����}����͊9"n��N��r��n+�SH>����c�7�����KӵH�ca���
�gLQ����_��Ӑ�[��Z�����{6�V���R����-�wݟj�,�)���mغ�`SJ�?|b�>������Ԉ����X�-������ �8�(����7�O����v���vQ����
����_'B�J��3P�)c��q�K2��1E��hDī�r	���E�ʅBMlG�.�n�����"��5T��^,rY� �j.�Y|��}"~A�%�\gD+N��5���2�1U��3Y;���e������tL���U�
a$&
m��Q��YD��KS�Gr�*��Ap� r�7m���������m#afrO�����ڦ^��j��I���5�7���L�d�M 6��`��S�q.1�׳ P~ѓv����&��W�%`	X��.FgF-��x�[r%C����ѵSȌt����P$_˱WS��S�ܽ��s/D�Hp8n�� �6��!Új�V�|�����*јPQD�X��p�3�٣k����a��
6f����
������l�,����U��;e�2I���n_�B�R�Vʷ1��y�l�Ь�(��J"�v܈�������O�����~���� 0���S�t�_	����'��䗲*]:��ຟ%�~�-_�i��N�H��0BsT�'�,ud��N��-�#��,jp�����6�x���	��/�w#o��,[ůR3ʠ�^�:Z��̶\��;�y�ႁ�
5
�r�2e(�	e�@$ޒ���ʦ�nɃ��%�Q�psE��"u��	#4�����	L�#���c�}��e�����s�N�k
k�����E#j %uvz�Zn(���u��*¡�]��X�3ډ�p�5�Rh"�qI6n{�]^B3;�"�:��y��<�O�y
��B���l	�h0��}�U�m�jk?��,x�9�X��U�Im�8���.�>�}Ѫ��z+�W/*���U6�	���� �Q��Y-�3}�&�O��ת�^?}%��π��ۻ��A��,ƫZ�������|����h�9�"��ws��p�Z����&~�z.��]�u�b"�P}js�M��Xdnu�{$��R:�<��m7�sn>���HqNQf� X>�P鈥�mcU�ݜ��ϜãFğ7�ϕx���䜌�	rU��MD���K�� k&��K����J���F�]
�l!S���Du��9^����א
��������NW�L���	#��e�@aj�#:"���E�T�Y�YԹߤ_�~���ia��*l_ȚΨ+�A�c%��6C>�0���E�w$�!�LP��M��/ƽ]1�eƈ��1<�nb���nd!�v������U��<$]���P�C�pv��k��W'���cN�"��(�=,B5�S��9��Ux��(����s'�q�z�0iA��:����gp	?������ƫ*��E�"d�F��r�:����oQh�g�μ�#4t96�:���h������{^���k[!��*�����P��.�2۠�Lh��(�(��R\&*�t��R%��Y5o�}�c��$�a��A,���X��:�G��F�N�����\���P�rh�4�7�ߴ/<`�1_L-���e���7ÑO2���V�E���e���b��]%��@���c��5�/UW�wi�^�h�F��>}g��ӎ}�7��
#�J2��,8�nq�U�A+�����O~#l��4��C}*S����c��w�Ήl�o�
���E���:���Ge25<���B��}|&*��0d}o]W�
ORb�=�J�Y��w����;�l��F�@��k��F�k��I};PkX%�u0��)����ع���5�)����f� %�"��wY6ǝ�u�����m|'ܳ�'zk!�Dqu Ƅ~�J=�[���7��H��f�TŮj���o	)jg��y�G���e��)��|���}��~��Z-��>#S����
7P<OA>bu����`��VWL��%�	��W�����r��Q��'�Ħ�����ZY�"�#3d�I�)�I��g}3^�oL^�Ղ<�zap;Zx%D�Dx�TdG�l��"[�rã�ƳI�{*I��I�ͫB���o�O��Q��E<gLٺ&�j��s��˾��8X9�K�B,���v�x��J�r�Zc<� :�{��WH��2I#�����!¦&�[�["�FM���|'�| V���|���8���6���;b3(�.!�Wg+��y���?���Kd�R���
����Ζ�x �}R�ȝ�s*�χ��~��i� }v�& Uu!�amh)�+{���#F�vI���D�!/;C��e�p51���O]߲���c��*�eP8��T�����=�fVz���t�h��X�ɳ?{���3du��Q�سlQ�? I� �|�"�sԈ���Q_��~߻�:-���m��P$���D.ªꧣ!�}r�����mߵ���#=�Zj�$�=�^=��^���jC�.���OFI�&�Y�Ќ��uƾݮ}���+��}$B���[��ׂd�}�8þn�F�UhH��TM��	��:g<n�:tiw͚�'3��6�Wt��D�MQ0,e/��Ћ�/ؚ;����C	S�ɩ�r�)���y8H�xx}m��Tv��@�"�?a�e5�
䐁9�w�o�j`S!��9d����bD�W���ʀ��7ţY9��+a��Nz=��RG���w�b��QpQ�*�����x�Q��%��rK�G)��q�<mw�Y�&��|]v�j��r�'r��[�=�*z��e�R���Xc*-y�YR�N���u5�\�4\��5	�����H=�j6-�����6��0"1@<���W�4��kt&��Z��+������w������*�����c�h˾��X���V����}�~�j6������r_��n䠌':���jGڷ
�
y(���*�_��D�IF�|7�X�.{լ��7��� �	�"��Fv�	T���a��FO69��>9r?hw~���B�ȓ{G��<��|}y��E�������R����}a��(��B� 9����;�.N���E�UB�z�C����i���!��X[Ա(�#q;^ؔQq��k�,cO���俱��qs��عV�?4	;ޟ�'��T���L��*K��n�G��&׺��<�8<-��r�e�x
g2m��ul����Q!���?r���ΩMY5�_P-�]>��lthcs��C�0x��?t�7�1��<<��F��7�	����!Ɏ�,s(1�[���D�uU�����U���!_�8M�s	��7���s�L�-�|=	]����%D��2n�8�ͦ0\��G��lM���z��"K�n��Pta@����l��vArǫ8h՗�����5��¹_�+��o-��B�����͟9��2�����14g$�N����g�k�x9� "�<:^p��lpsg����89��U��~����"���R�j���ɊA��5��i�����Z�����y�0��pyه�}��gg[B$}�0�IowF������:�߿*��b2h�Ƅ8�Q���F�3����4nӼt����ݍ��okjE���K]��^��\W�O��.���</��ba| �Ƈ��F�9F�?�_�{��0�z�dr��ik�j��Q��\���`@fNO
��w;
�P��s����Gt(*��!����X�]���P�B��;)��Z�f8g@�E�&k!}O]IA��8�o��l(x��ʴ�'`uB����d��`�x�2�jM��Z��2�6bI4{U�]�K��5��r�6t����秎L�'g s�KN491�z�0�����ײ��F��*B�c\{U�G{����=��Up�ͽ��&�=n_��ok{�i~��m��:P���0�<��}g���S6.1{�Y�����K�|�3��JU���L�k�����������7P�Z|����ߖ.���v�G�PEa�E�Uע�Y��|G���eb��02;!818en�nu����\~���#�C���%?�)b,׵�0����,7S�-�X�Q+�M�^ᩤ=o'YV����^r�KG�����<�S�^��n�[�(!���=DԬ��tۺ5�/���%���F6��F��=�g 墳�2��a�<��妩����c1*.�w���\f��}�,�m�,"*埳���l���
�-���Q���p͹[�&^KP�,�͆��[���u�&85���9�K�0��n�rj��~z�+��5nĥ�>ۻt��~�c�Q�ƺ�P�U�A2"+<�RE�L�z���)�z�ZL�ٞ<�G���A�l�rۺ��Z8���<y��'b�M}�f�r�̷�_��Z�/�e�%���ˁcps{])���0�'5���5O֍�y%�א]�����{A�F�C���w�{���gت�5�ع��1�]�YTLh���[������qg�?��'�/l<���D�|*�"R_{��*n�6z����C5J����8g�U�<f�t2�"��Z�-zn�d����	ǧ���iU��,�/��y��9[L������Y]iB�T�yS/v���g��i�4�KJ�����[ד}�4�1YcXo�[�I��q������-'�G%;����v��d�g}���5S�-�����tf�Έ����&{����B��e�e��,��@�Rq�ᒁ����ԽM}ֆR;��|�z�#�Mu
�̒��p<R����v0��j4� r.i��x��V�/^��Ŷ���"�O���"3�sҨ��L�mK�|�a��}SI��z�؟΃[���@��g6q�_~��@�-�����|.��6c����_[�:9�o*�����䟈�% �������c{:=E�U�6RA1(t{���`f>�#����͞y)&���64��ZG;��y�f~V�( ���m�6�6�)8[�1�2R w��D=��b��8���$�/���g����E��x�c+;>�3���qɢf�ǩVn{�ؗ�LZzg2�o��$Zr���p�����90��:���T�~5��ܰ��&U�&�N����=W�Z7����������0ː_ɪBbW�wۏ�-q)�M��Js%�V#��OS�T^���aޡ\������˗Ѱ��|R~�>�e'9h�T=�j�3�X���4xcۜTjzt2���Oݴ�a�U��ޮ�Ul�8�/��36��S�&��#�,��ۉw���%�k������*i(|vc�8���n�"`7��Z����4������CR@u���N��e����Wԥ
��k:ض'ޝ	M��{����1�xZ5�"�\}�'�Gt�@�M�R��ķ���j� �^Ũl�#G;%�ú]��`K��kjZx�<eV�I^����gP��}FQ�P�n
��~�*'5b��j��BF�*��QM�QN����f��a�U~�.B���rQ a�Zy}�b���ˁ�d��ԑ{/����֯97]@Ɇ܈$W��7%K(�O�4���E`1�"o�u�u�}(���KY�����w]��������
#��
w��t�O��D��d$+1��\;3�'���rlc2p�	��H�n�("J�n�c�E��p�{�V ������Ct�s�G��>}Q����ә��銟��QV�}�Qt�X��P6��7҇��-�E�&�a^��S}����?m=tܚ`+N�i89�apx����U%#��'Mu'.�(�Zi�jD��><k1�] �( ������qIS�Nݼ3'���+��ҥo42xf���UZ��Ca����'���Dj��b�Qt6�$5�^�s�����R:W�E�P���@'\��JoAT�U����[��?\���H4 ��&I�F�yQn�:F��ٕ��h�����I>�j����QK�[�[��:sf�N>��!��FxI�QD������p��+�a� �d�C���E�.r�Z�GZ��n@���Cp��WNٖח�UÄ�����<�ņO$�[�����������bn�zB�������%�c,cFX.��\��ĺ�85��tᨄʐ�'y_�y�]����y����}�+��N<��4�ȸXT�UC��C�x h2c������.)�>�S�A��5�����$�6U"ݘ�*�2���t>�e�XR������_�W�f��\?�w�S����w�r�&�$Ώ�j������N.��yt9������R�����R�j��6]Ot��?���16J/Gc�!����o_Ɋ��t�[�9f������^%��IG���>a;�0�íll��V�Ab{����2��ͤ
�vi���R�5j,�P�0�ZNz���[a�o�@�䳜��>�ȅ�"D�
��ǀ$���H;�B]�ڜy�ó+"�G��	KG���50��������{}���o�ho�aOmJ�T�s!<5;��R]��t��ʸwx&nm{��A@��p4$��D�7x�����~\ ΂��L�+����U�������	ٖz�v�qH
v\?c� ����oJ����{��?eL;���fjغy�Q9(����R�%!�5�P��l�D�,r�� �f����09R����𵿾�L�*q3#�����b��(�k��V}���\bWY�C�Sk.;�8��=�-	à�-q681&O�Q3X0�r�XA�evNʛ%U��;�OG1��[TG�e��g��b"�<��4a�%w)�2A-zi�wՃ�D@'�Dj����ж�LzmL�E�k����ُu����YV�5m���K�EK�Fy2�2#'���ܿ��7�7]�lHkj�H��&hN�n���o�Msӓ���I��|bQT��솁#�G�P�� �y��e��nZ����A�&~��;�N̢�0�\��8����Sd�	U+��|]�]3�x|�s�=Hc�F��Ul�kC���\4�)8��"��|Jޝt�ְ�d�����ߪ�T��{�.u�G@�KO	�G6�`�O��kpɺa2��7��y�l�	��Y��!P��+a���:ŸUyy"k��h�9*PAg߃Tj�l�9�1) E�yx���X	_.=�mPd��럤1� �lQ�{M���Q&/�W\wQ/*��l;Ur�_v�y�&(��"��w���fB�"������~�|�?������J2��	b�]z4�k�bn�;x$�Ň�W���㤳v2f�W矕�S��q�M��fWNDHێCr�٩��f���PlP:�X"Y�i�=�3F�Ǥ��^�|qF=�i�w\��BWB>����99b�T�L���s�7f}���|��(��T� xftش�G���W�=�U���r��k{�V;q��Ȓ��^�P=�A�V��t΁S�(TRSn�*��|�W7y^~R�T�6B��a?2��r.�䟥շ�(YW(�u��?��.��EY���6§K�_p��3�kC�v�S�I��Hj~�F_���d��14RWz�6�0�;�V����|�s���i���n#1Hu�c��˻��VI��so�fpߘ�)9}�(��R�3���6�˱Ɛ|��Q�
����m��~���=��/�&P?�d��\j2q:�YN1���1��{Bz�H�G@ǧ:�}*��_��������#P�}�f�j�cI���$>b�ؒͺ� nO���4n�"Y� ��E#��i�z����á�H�^C��$�]��U�C$]�g�<�����Yo��r��w���a�1G��H6d�s~@�9��a%�f��E� ��/z��M��Z��������������W�@��f��ܣJ!"\�wNK���G�=%6��j�6�_����}��#���� ����p��O�Q����}��[�$ !�vM����̧���vR`��׿�(�����$)LD�r����͎.�	�i5(kr����J��|U� l��\�D�=A���*W��U����%��MϏ`�gL��zR�|3����l�a,VR��PE��[���B�.�z3�x�s�~#�IV�
j���}��%��t�]S�`��Y�@��v�0��p��ò[����n4�5I��e�TZ̅`�~��� r9xgJz"�u���^�2�!�5u��5� T(��.���'nZ�����K�P��p�h�� �n��ր���x��W�^���K�,��e��'7�рP��Z�3��J�g�U�j$�[���<�ܷŰ�Ӫ�$0pI��E1��GTO�Q_ܓ��TY��X�Bq���g�NKR�i3]�'�1���;�^H.�� _J m��ݓ�+a*����V�Fd���B�-��_���tW�n4��t�Ax��q
�J���3��rͣ�����u!d�;͡w@��h�?�UP���en�����W��r��������؅�ꑧ�T��	�c��3��t�������	���s�	/�Ѳ�r����ޣ��~������FӞn�uxwaޏ$A�<��U��K��Œ��Ѷe�sK�u��p����gx�7��Iȕ��d�g�cr�X���ĥ��K诈f��Q�ҭ_���U��'$�`��7+��i鵗�t��&$:��7�����1�=r5�n(�ǲgfMIf�����*���ߩ��Q�CM�Ϊ�O���,�-�WUg��RP1�H��kj2�����p�����;c)l�B�2�Ns�U�wE���!�Kb+p�N�4��)��>��n���#�[�H ��GF"="x�Ϊ��٧��>t^}&��8��U�D?�$8�J*�޿�Ư�-B��{�����p�@8�\�Vl�41E���e!�/�L�e��c��%�@̼
ٟƭwz m����sk�g:�c4r��k*	ʱ4u��@���4���zw>,�%$qk��QK��%�5[�E��Q�`��|�6z�;c���37�ed�Df,�3�Z�
������yA�
JE!M�5�5v��.��ל�����vQ�$� ��-ކ���U,@���{���ʎ������nw�����(�Z-����3�SK;?umkm�\��(:�.1�%�2^Kx�3�<�n�^ʚ��׽i�C�EC��I�z�B���6���� �ؼ�}���������6L癰&XV�tW��)����Z'z���vp5�?�T�S�qh�nPҁ4_��a2&zA~F���������x擆N
��ķݭ@Ǌ_�D��C��U�2E' ��4�м�
�K�7���wq��CuidA�)5` W�J#���+�����V�� Q�<k�m�3I{ҩ�?F���0*�)���մDS�<��v���Z�ˤ������eraUHR�@�LJ��'zZ]�G�+L#u��lly���j�M���ZEe�[�:)���ʞ�]�8� r$j���~̖X�\h`����@�/�	�Р���F�UH���,�[
�-yؔ��=ϒ0%�6�NL��� �(�\���*��+*l��kHv�`S-���PT��
5����K��A�8a�VCV8m���
�+�X���c\�r�T�zr?P���\ؐ�z�b$ሓp
�:p^4��������P,��b���6�����y#]7u����L���;<<.r[:Z��Zr������F���!)�I̦��`��s����Ǩڎ���a��E���6?DN�o�~j<kԆ�r�|C�k���");>�˿�R�h2�*=�:i֐}F 1}�V��,a	�ڏL	:K{�K-�Pp߈�L�N(IA�3�$�|��йs�s�O�L��m0g��B_?e���L�L�&�_�d�ѧ�sSe[�K&)l��u�|I�{m���~ƅ�U9�D��OD�{�m�p�U���#�)]�Q��������,\+3�^��֒�"�zq��r?�I^�:�ϏvQ�U��7NJ?������H~����}�"� l�j[{�0�$]���� 屢��0s�X���σ
�tu#	��{���	h�̹�,�>zᘤU�D@�ј|�C#������cr�s�aC��x�Rt)\�No{�Bk��4�@��].�=��6��*J�<�>�oԳ!c���`c�U�����wgf�A?��bT{�u�������|�甐d�ƈ����;��#��tʻ�����T�5�'L����?r0lgC�sHBk�)���J���'NQ�]�
���w�o
�؍mTH�������P�K|�>��h�F�cH�ȅ��'��W*D������<���:�.���B��*�t3��^����*�nǵ�+8N��ykm�뼱W����\Ԙ�q�R��v���R00�d7מ�O��D��]h%�;&3����=YA�pS7M�.~Zz!��c?,�n�~�j">�Bt�^)��T� ���ȝT�������ԁ����ֱ��,���2ߣ���/��ܚ*%���m�������&��!r\v�P+��<��!��~��@"΄��^�Q������yL+�J��A+�M�V���2��pg����V<�C�ֶ$9���ɶ|�:?@�}�פ�.
��k�g�yX2j��}�]�DxRϐ;�xYR�YJ�'�(c�?�V.�I���� ��"}�)vj��߫vvW���ǈ�?AؠS�����Ǽ90t5��"�i��;-��u��_��>0��ӫ���Ӎ\��V��n�Č��35	���H��5h�� 1"OJu�2�����`/�����<��V�i��^D�	{�eW��rq������0�*��1�ț��@rOǾ.�K*]��r^O_�*d���[�W�p��@h�g�������R��d�nOyd/��Z��]$ޏ��T�@�B_v݆��M���s��!�4�#%NUH�1�E)��k'c�q���'L�5f�)gN@��"�I\#�?jQ�v��<�k�͸��r?�#e���^qoC��/����M&Bɶ�s�V5�wŕ�����@�^�	C۹���D��Uc�B2qk��0���{��DU��'�G@�`�����
�*Ɗ��������G��`�OW��8	=�����P�	��ysq�V'���l���(:��!�b�)Vڒ�~�
���eW���ia�t\�=�d&�,��O�M����)�v��.\>��ń��K���)]�5$��(Nèl!3�ۗ#ٜ����!�	sX��G�I�_�ջ[\B)�w�xi>�-,CP2o�-_zP�!l-����'7{E=�p&����ܵ3p�قIY� ���ç4N�rP�H�Ц`�W�F<_#���j�r|^���P��ΔT�(ZO�eC@&���{^r�rP��x��@rv�gc����;��(2O��b������;:���l��Un`�Wu���s�G���1��[�������D�:���)A'l�>8��T<�?^���DL[�1?���)����^'���"F�Y�W��'��R�ۀ'�nga	'�u��f8��!����F4�t�:{F\�X��'N�H��	��͹LUh��S��X��m<t��re2շ�Ϫ�;o�M$C�
:?�rP������s�8O[v���o���y�����T�8��BQ*"B�cz8T�S��\,�+��7/m�M��@2v�-�u	/�Vʧ)�f?>������@�7]������m�B����X�k�?{���1ٛo��u��¯�p�W���N�����ċ<�Zu����H[R< �K��fF����o�K��(�[D`T=�Bq>_3b�y�4�*���G-�6�np�k]̪A��H��o��	I�7EEC��O�}�b^���`q��ƞET�ٹ�0����Nτ��:�ޱ�s����=���;���_�X\�欟�@u�0�s�ȯH���m?Y�6�I���������wN/�GYze�:�(I'�a+��\�F9��jL����~Da�r�5�� ;��GH�B�n����3b��e���_2c�rc새�Gpz:��d������$J�+qM��F�͗�æ|�瀈q�t���N���Ri=6:|����D�y �,�sK�7�Y��q���� �H��NC3�?�x *mP�&!BH��[V�o��q�Ȣ��v��őf�N�
A"�����1:ƀ���'��^a��oi	9>Q���<�m�<���yS�W�B�ٍ��X�WIQ�W��l��H�&j�l�a1�Z*f�ԸqJ���MD!xk��D�d$��}�%Qn\b�W��j��Fa��T�����Zo7�LdUu���~&����P��Ժ�C1��oo<�Pm1<���RQ��o �Fs>y��2M���?�"���<�(jRf.�Ao�8�3-��:(�����Ԭ~�'�2�{�I��.��r�x�Vܲz�SJ����c�{G����%��C(�>Nmj^-�?k8*Ml�ibϓ��'(����������Ư[!�	 ��xak�ϰR~��d��x%-��|_֛��4�k�-k���3�<�R���*��`r���+஼��zD�4J[�YW�HBdЁg+�g�rn�6ͬ�C��i��-���J��"Eެi8m����� �t�W�{g���>�wAV�k.D���6��k%��q��mR��l�P���\�|Q0B6��5ze�ŭ%+!3nKz�a�|CA/	�((���Z#�ܢ��{��
�\p�I�]^��g��Ǚ���W�ڴx�Հ��νɑ��S�2
�M-�ؓ(���c��9�[;�q����0�d��L�o�����[�.��qa3I
ge�X&�}�?�d�;��t��Fw���\�H�mg���`9���P��U/C�r�ճ�z�"S�R4F/ub0!��fCxK9�3�s�n�t���Td�Y�]8���U	(;���� �%�8�8シ�S��$�oX�#'(�̤A�f�	��Mp��Z�ml]�6�SJY��`�hx�������f)����i�v��� FLr�U������3(Ȣ�z��W�)���i5����i�!��
@���t����ɾSD�3p�D�B��(�g���e��xO�7u:A)��f �s%��'��Ed�}�).�VW�a�T�-���?���$�CE�/�Pm�<��ӕ�R����ݶ��?���İg���?r��������H:���C�]�3�ܵ_��+����cu��?*�mF��r��:EC�{�Y
LAVo�㲛�CԢ���آ��!'�����k�a:�X�\�oO�x����?��Z�Q���E�dW����l/�9��
P���(�&i\)B���J��[��������D�/2�����lf��K����kH 6�+HZ�([;��QfZ�4����ag^;>׺���I�OX:Ū�����B2c\��9U6���Hh����MCy�J��!�͸��h��c�����KB�[�C7�:x��nu�t|�ζW��߈�rԞ�]�q����/?�R�&��JpΉs5��h��x���+�����FCV#��-���7�d	ar�&��S��Ƕ����Wv �"�'�ܗ`)pc3�h�����3��@��7-i`s�9��B�����i +y`��(�o��
)�
,���11quԉ�2�Ka�D��AP�Iv��vϰ�e¤ 7t�j�KL�`��}���=@O���7���@��uq��yTQ�,���M
]��[������NR���1���hQ��f�nqc���U�^��~����U��ĝw����90�ƫEx� )M���EE�����|rv�(]���|�v92FQ�Y�΃W�Ӄ���H�4ɀX/��85�z���~�ɋ�q0��/&�eG������f�V3|3j��|�p㑚��sM��ۋ�߲��o�"��O&���hd�J�-��_V>ڤ�L]�^�������T,)�y�l���h��P.����2�l	&aK"�WL���ޠ�Q$���Ș�C��(Dy>z�D��-6�@H�Ɩ|l��K���1�I@�>r�f�LF�tP
#^��E� '\�f�:w�8㽪��������J����{.�d\rJ(�5I���b�z�GZ�5֘eS�:�ys+3�����_$�Ƚ�&a_��#1u�ۣ����
��e�����V��F�ڧa���U}�3x��V��?�J������4��?.����P����&����7O,�Ag��x�1+ISe�0h���p�lcԃ�i�x���V^�\f
�F������^�{m��/X�e�Rà/�B�izC�qv�� ��C��&j�ȝ@h�q���ڈS �e^x�{�����-`�����I5�1���#��Ib�F/��� �{�F��h��4�cD~9�n_/�F�D�_��!������I~@�,[�u�S�����f���`���3����Yg�D�KC�_�o��Y$3�(��0����HU��D`����qN�����X������*6,�_! ��?���b�g����	�` է3
��]�{��k�0Y���?�my�ۂ'+�L�j�B��P�-=s��D�$�^���Wx�i��>�<��P�'̗�׌�Z٥�!�ԅ�W����[$�3��-��kW�C��3�l)��~��	�8��<%�˺��������{5��&�,�5�P/�G��7�-�s��35��M��� �9����L�~�[K�0gXzyS$>��n��#��?�ip,Zd�&d�}�\4)�e0�CR~������pb�ގ�r�U>y�,�W�5*��Q���GA� ��:����Jlr��:��5�ONfrfhBGsɭ�Ni�q=����h�(��h[��8�`���e������Ʃ�q���PJ3������=���3�G�*��%�ńHx${{�[<�ܿ����f�[�vͯ�1��	S�wN�8
	�q��U���m)(���*��1A����s��+ͩpU^z��Kc�����e`�iI�@`�)���^2���#}�d����%�.�8D�u⽮��������\)-l��Ό�3O��e�kHFę�t�zq1s#�Z����\`��R]B��*�pv�����ɢ���U���LB�O?�)�yr�z�Uoͬ�-w"	K��|ϺD)�a���u�%��� �jv�EH��d����4������T@r�}�G�+V�b��{�ŭq� uE�:�.�8󨵖��$��<��u�6%���Pj���i'�S�p��

���^�s�F��sި�I,t"�(��*ytNû�{-�zU�����^)��G(3x������!��L�ek������	���[�pG�

�p⃮q���(2���������ѽC|<k2m؈�����»��`"�JQ�G�R{��xطT�NtX!=��F��ӂ� *��^,GP���5�49��/skKa�o�G�?�_z�h�04^���N�z[� TAt��&Hr��<�d�p��EAX��/�zӥ>o�U!�uc8?������_���������|:�=�@Ώ��|*�.$�5g=��R���u������
�& Af�{
��}����q��Q%�A�@�a�M��1���ԱHd�]�H��×���n��!�p�LmA�Zu�Yg�B�L��и�^f���gTd28^�-e��-���M��E��}����D)���P�aPs/f�(�^N�KMAF�@@�|�m:|}�1SH{@oV��'+^\ڷ�}(0��\{Te�/q�ۙI�?�x�ҫᰆ�c�%��o�Z�1%�[�G�Y�<�b�p�<yӌ��d�E���ҾYD�q�? 3��g����P���B�����B�]���0�J ��]lhH��*h����]�1�|4��m!i�|����=��eĴ*p���ף���s�S����%�j�O�'f�N(�Q�ѮMwrQ��Nt���>i�[��JD5+��OI2��Y����!P$�ѫ�{�"]�[��-1tY��*��82������0�C̀WzX&pW����:������F��4��2��{��Ē{����%�E��~7hv� I�#��-���{Ǘ�wz��x]*{�Y�a�$��gS��g�o�\�
33H9Ē��d�匤J{[.��"����I�{�0�x��1�3�狣�M������V*�N�˻�^�1����C�8p�ɠ�0q ����We@o\ ~?����~������������5�©�r�n��=��w]^6��H��=��xk�� ���e���Ӯ�# 4���Tf˪��}��L���$��H���	j�n�+=-H0`��X��w��9�^D'���爈��M��#}���8��fl��%P���d�I���@a�1F LuFm?�<J��y���EO@�A�iV�:�VÝ���[b}H7����`?Q��+�kX�M�#�OVѢ?m'E�"��w\.�n��f���@��/]o�u�}���WG��"����0��bϤM�LJf�tj񣿳칙(lb0�xj�2����3��7f�@�ǐ�����f�"W�3�{P`5(=�>X�r������]��;���2(���m�ķ��ӻ���ݒ�0��� �?"v¦	V:]�H�8gĕ�,�B�Eg+��x©ְ;|y?�BVS�����,�%[b�ɷ�TtYMlR3��ɋ����d�\�PV虑���9-�9)t���h_i��e (ьN.U���w%�:�M)}3�(�Q�C�nr
�[�%l~b�~�B�����vf����"����ߩ(������Add�2OcY��O�?���8��\���X�¨lp���J����R�ɦ�Fj���~\0q����5>S���Q��kj�������ƣ�0/�	�W�^�^�E99W�o_�+�q�!Ĕ�Ϟ��6&޵"
��Q�V$e �]%��1Fn���jJ�n�d��l��6��������T���W�>�<��
����E}7��.=�Y.�.���NS���C�/���{?g�ޭ�!�	���Ž�p���<S;��Xӭ���SҨ�����	�ݸEu_/	�̣>�D�TxREx=�N��a&�������}������7�v�@�����H΁����N��C�}���N����`<b�@&��K�M{�&��kh��z>Ŵ��\�Z�wu���n�lz`1�a��`�u~�U^�+9��i�Z�'Ђ��C]���q���(I����0�r�(ez&�#~C�;_nn�l��Z�B���v���H~!���_R;|��Mb]50	!"�W�~��ci_N{�Y?�K�%�'ݙ��g���IH���P�	�wwZNs�#נ�29I�4u����ˉ�Ķ��|H�-b�(}��H++@��d�}<܁�!Xu:�~](����[������|XWrg�#�1�`	�UbB�#�f/���o��G�	�B��,v���][���2
T(*ւ��KӴ)1=	D�����ą�������:�� ��e��ȟ�05y���[��]`�s:S=<`��(gD���;�r��p�s5W��f�[�����E�����Iz��v���4Pj��2��Ab���WF�G��I������e �D��G�۾{�����t��W1�/:����x~$�UY��Ķ�����������BCF/��q�u�@���j���/I�mɞ��B� ����{���P=D����j��h��.��kJ�*wI�
��x��˩�������M��y�Ă�z���5%���4���QB�	=� �����iB�W��R�������2�M�C�M��k�:�A\Z�9�A��U??]vR0)��{��s���A�r��|jFu��C̸P���^�%j[ߒ��(nd{�n�2�� R�Ź�-����H"�fw<�G{�#m�#@w�̐���-�� 0��i�w��TU�;��MU.�=m�3�^ �sb�?�$ �X��~fUk�>�����5����X��Х��aGo�R��O�o�L���H�p��d�J�l�s������5~��Jיc=6��$+�F�m��).[�وk�@C3��+ �D�/''�# �YD� ?���KT�zc.�=F�;��'eSf�1�MS;�p�Lk�:Y�&n%)�hF���/��"z�$̖z=f�9���[#o�ުu�㦖���Ƌ䭕�+���b`E1�d(D��1�h���@3>�Ͻ�U�`����*'��8���z��vo�� 5�L�g2�K�:�ڜǂEm-b��7�� ������^p	�w����jlT,?e���LF��qw36��"i9�����ۨ�E��V��}�V4d<�M���ԶTKkv��)��"'=ʳ�8�Ӧ�.���y���R�k�J�g�'�as�5�F�{�G�bxQ�@���Z;�S*օ��r�>gج);]�V��|W#r��}�	D�r3"�`l���\�@ߑ=�ԋԸ�Py��_�nq8S��ng 	���m�Vԋ΋\�; v��5��Z�)�*+�Z9 H��~��d��3E}c-Ց�\�펠�gkQ��|���G[���KaЯ&��Y�c���B�]!b�0����k��\���^���W[�*�F�.Azz�C��V:�B�_kVVk�����a����������cX� ���|������~u�hÁ�m������@ɤ+��c��q��q��L�~�����o���U�Q��It��cƐk=-K`�Y�r�J��8�$c��k�d�x��%f'n3�?��k<�S�d�8������46^:�!#�\k4�`�ؙ��Զ�׎�W�h��hiɴ��F�s$�~�r�Wz2y��*�*�[#�w��m0A���\4d�F���4iLD�M����j2����Sv)�װ����L��Dv��\�����B�N�'��7sZM�N����%��p�q��MV����m��l�t�����ÓBdqpWa��\V3b���>k�(�߾�
���%I���Lh�֏J<��O�q���2R�b�2p%�Ʒ�������u�k{��Q�R^�8S$���f�a7q���P��
,�*	�%ḋ�}�����^;(���:���@C�o������R5k�%��B=a��r��3�Η$�C녘�;�Mt"�I�����B	`��L�zd��/Oӫ�X+�"�G,L|	��	uyɲ{�?���h�cb=ū�\c�%�Z?��0ٳ�h��~���F0��%�+	�Hj3���h�\<�	�q����*�u�I�Tk&6��8������>{�?%>*�-c~�,��}���`�X]�si8ڜCiRr�GY�6����8�@X"X�lic�碙3_O)s�XFPf�OT��f����qy���yt9�b�w?��iWH��Up�E�T�wQ{�_}&{������:v��v�0]��Î�A��yW���EH!��$�m8�\ڬ>�ǭE�K�ܮ���������������"C��9�� "k�������)�A:��b��"�⮞�����&-����'U;*�Fqk�L`ϹO`��b�O&	����`��2|��*���@@�Șp�J�����N����1�������"ɷ�y�MY��=�0�Ұ$Ȳv0��}��I4g��v |Ҧ�xD�Y��-�h�*�i���q���;Y7�7pr8�,�L�ˡ�Ӌ}�pW%9���]k،]�Ea���~eg������+ �
�Ϡ��"��i�"�V^���-�s_?�0ıfQ�j�Ɨ\�{�vCDC��>�C��	<��0���g��R(B~Joh��'0ӄ;�+���&�&?_�Ѡ�O�J}�9֣��J�g�Ux���i}�rc�3x���Cz`�t�Gc����D����dd@l�����[R���L#`Qn���Cb�N7B E8�*������O֧����C[٣� "턖;�VR��X�?�?7��스�%�:�пn��T����[���ȇ_�̣���-R9��y�4qg�U(|�U4��=��LS>�%)��p|[OW0�;���� �9�>A��i:0k�a�`5��[Q�y���4�����8�h��`���"����i����d��Fn��1c�p���F&�U��-��oݴ����U[4��t�}+/��t�S�2��{Z��RC�B5-/�f����_P��|����d�5�Gw��#k�Q�9��$��b�&��vx�
�	�`G���5����4$�%�Ǿ+c�4�9�c����eX���/�ڬ�ua��{3@�[;�9�<���}�_e�:4�������c�����{Yր��p=��Fu�o �j�=�zߠz���l+��KbIp�g����w�냖���D}	��� �?�}S1��}�2�Ʋ���qP��{��M�tvN�80�O_`bp�F+�f&�|�šU��V>fKʩ8@�����y"G��6N�����ڙ���:Hg��5<� }����8�O���Z��K�����߬(�ƫ*�7���2ONl��� e�o����yRW���V�bEԡ�WBZ��(!��a��|��g���9����u�ד-]6ň���I��G}��<��6;�p��d@���2(�K�'͝Q�Zz�
�LA'ZZUq��W�������[@X�9I�q�Ww�"L_�+�OJ:��w�z�F����̂@?��"X�d��� +�A���lPa���k� �O��x���p��Q��U���ˀ��m�\�A������RY�a�K|K�\��}JNRs+�I���+�e̵�}�����.���6���G��5��F�{E��YD&9�N�#c[�D���_>�g��q._Cuv1��]�v�<�~b����D��}��@�}�'�V\˦3�7�5�%kv����4]�  F���wm����4���
"?�x<���Ds,�Ǐd��5u�2E��Q`�ȴ%g�To����1 ^��s�BJv�9��,��߁�͌�����5�p���kD�*���ȓ��"��eg2��	�����:�QV���ſ��l"�l�Ϙ/���������.w�J݄���A���@BY�Z'�}d�F�����+�Jx���=Ǩ�����ұ�l����L�~D��FaőY@�hU��p����]�^��%���t#��dD�S-d���=�qMA��ww�����ɔ��I	�P���Z�&$�&��s׽Ž�b.xfƽ$P�
s�!9�s���_Km�'�K7�:��a�l�9�����<�Z�"�P��$�.�5��$@N�ә��yLW<Y,�&Y���GT���o�n�<P!�9�����m�|m�y��.0�݀�N����v���Ҧ�d�ra�V�^��P��ڼ��1�J��7� =�{�\�mr|K��8h��ď}�r4u�yk`�����̹Iu8Cp�[]��7*��g��9怟W:fVd��"^�����O�|������l��a�����8�:T2ء.A��0�w��p�jN���0�jI����ڡOB����jkb�23$,��"}�'&@D���G?ҴO�D믱���>`��KlU�" �	>'	ݴ�5��5<�8�m�l��<�P/�.Ʊ�Κ��Ňzn��yvm�X�1�2���=it�����g�5�1h�麧�a%S�+�8��sZFD1;�ѿ^96�?)1��+���u@���?�E.l�e+Kx�5�#[�+U�f5)����(�@X3a.���4��{*�v�����}3n1�����
�,���;�?3��]��0���	����2����Л���j�k/��Efv�]MuaS�"�f�9�j��h�@Q�2�u{��sCeēuRGE���H	LW��/ �U�[Ť!n��2�١�����ٲ��,.�*�P�� hzc����ޠ��u pPU���h�KaTȑ�S6iPw]u��g��Uq9B���Z�f�Z���Wqڳ}]�,\�0����m3{{�/?�4�Ӊ�d�jG�pn�B�d���|����s�
�+��pݰXO�����5��u���l:��T��ac��
�x;J�I-�����WA��fϯ������ɿ=1�?�~<JtG��/�~ܗ��O4���q��1�8�y�"�~�Z�s&J�kOx����:ڂ�úcz3��6DCe��h��X�


&���&����!x���
ۦv�ޑ����I��� �-WK��1�F�(���b�f��%	+�+}�G�d�n�㴢l%]C����[�_���q��Ĺ^텊c/����<�-�z"��Po�E�d�@����U�S�J��NP'A:�Wc�;���h�$�n0��+�<�ژn(H��]���wZW���n�@/P��BG6�.���[>�������B��l�Uh��x\�?ش.:n���	���b���cDHѬ���������2�/{�B��"�~ 4�R1�'PN���K���v6C��*@̈y�7�7Ǔ +�a��U��̔��������B�	"E�=c�4��<�L�C�X(mt�+ʗ��f;�7	��$�煖���j|j���x[T�bDp���FX#i�4Rl��������a]�ز�ĴS�ȀJ�8��2gR����'���
=N���-�쾬�'W+*~N�����R8r嬪�"9�T�,�F0�4���	�����.����#�ס۟�>��&�e������w�̌����1"�@R���!s�=�N(�iN�"w[^D}Jp��j؊���z��ܙ8$�Z+
��M��V���qQ`���N�c�Z����Ɏș�z�`�[h��͵N�lz����h��9Ө�����p����u�c�)�:�u@���}R��3E�D!��vD��$@+�mˋo�_O��I�Z73�Mk�t�k�mp>��A!� a�2F�]	���\@�GneƦ m��r�q�F%�U��>.߯P5���w���O)�'��f�?��`-�(^���!�?(-8z�t��>�*��'j������k�U"2�*S���9�=W��E��Qa.���`���/gAM���!�.���� �#?IB��:n�c��`�O�J�C�>s���-h ���)��?�S
��zXW6E�Q�I�,Wf��;��'�]E��l�3׆�@3�91�}���+�c�����y�>��-�~�QYc�E����M�H������78;�-��
^�[n��Ƣ�됷�������3�!a�e������p)�'1��W-���	Ե� B���W�ܔj.rN܌ݘ�T�ߕ��o�
���s��"�2���_�C|�$�!
z���q��4�tzű+T�6ۢ;¥ t�>��5Qv�ھ�"E�Īɯ���Y�-Y�(�	0�$_ӹ�vh ���ڪ�ݬѐ�on��DP/�ډ)���f��݉.J��`-t	!w�k����a��M3�&�T�S8d''����eƛ���`���E��}ˏ:��Ё7���]��M���+�:
���#�"�7�}H���D��%,zĮ�Z
�aD������倚񿌨\k\D;Ăr�;�Uo�Îfc<ą�%�{?��ز��r���I���_�S%�}��Q_���W��m�1g̈��!U-�� �b��?ŃgV��3U�g���q��qғ������pY�n�y�/��$�&Ĩ#�;.���R7p���浇�w�9#���m,��O
� �F�z�#��̩���<�-9}:�B)8|��,+6�_���8�����3�˚��ޠT����������Z��M'g�z�	Dk�7������-�A۩SXv�{��ߺgt�B����I,��ծ��{����p��QV(��2);�mC6���<.E�c�a�&�!�k)�}���
��v�q+�$Ep����{?��B�<��v>�W�@���Pk}��A�O�M��	��S��MK})�gc @�UrEz�19��m�/2�@AS׋�_�trAɰ������K���P� �M�g]ST*�z�ן�@�|p�K�r��������kF�"g�n�I��@K����l�\�;3�\��������;4�e-,4�zR�ѫ�Lʪ7�R�'��D�Y��B�P?RC�ܕ�Vsd��ͿY��Қ���޴Ϧt��AOcr�����vU��mV�S�G��`�
Vѕc<ȽL��ޤ�K�PH�Ƴ���6�H�����%|+�6���f!����qݰב:=ƽ�Dk�	E��.�;�����o�!�-�$���q��q_�ެ�(1�4��ݓ���zSE �]��7ߵ8/x�Kq��2ål���`��hn~L�:}I)K+���AN,�i�2��2�.�p�����[��NCG����[!��^�[�Q�Տ��%`���虀�ћ�\��b^l��dHR���SvS�L���iY��5kB�!D���|�BUI�puѓ�����Ak���U(���ӅvY�:c��4��(����D�5��JA�G�"�k�
���ک��4ħ3���\+>���p�DE��5`�C��4a����z�ge;�#�m�%��o�nܾ�Z��U�2(��R*]����Red�����z�l3���I�&�F����G����!���
[����Jh����X8*��ء�s��BCD�iCk\�z��%005�8��	Pz�Z���}����`Pҩ��x��J8d�O�H����s��X~�T9v2��b��g�L!��]ZLH���S=�8�5Q:Ja�Ղ/��5�j y�����zg��<�C7\�x�H$�@U?�s9�G���Y�f�J�I�5^��r��P�1%PqI����)�vc%�+z��x�.�����
�R�&C��b1��6����F�d�6K�u���
�v��]�\��͚M1 ��f����@狜!��+���ڊ�_ρ8�ꢺ���ڭ�d��L=����R�s�]���-2��"B�6���N����̭]����#��Pt���歴 l`Z����7E�T�8���QHkk#�h{Ql�"�羄�8?�}"NTf^�K����`:����h�E\OI���aȅ��*h��e��l��c������Q�EsI���_`(TM�J�[;�.,z�]l�'2B,�_��M��
�g�V�D?� �c�Ӄ��=l�b�:U�͔',������ ����u[�Pޓ��bF����h$׸8/�x&�� n�*%E* ��2 '��;z�Z��hђ��;�ރ B�K�^ o����_ ������蝵 �Q��_I�SOV�cK ۅ$��jv���(���[��뤦Z\��b�u���%������o��%��њF'RA{K
��3��ŎXҧ��ļHNj��y�xB����/�1&K��t�Mi*�GP����`��!f���k�O*�&W�|I8�d��o&�W �󷊆�C��2�ofz!P���x��gB/&'���Ӧ�;���p�v*��JfŪ�������I��4܉��:r:K_���s���;z��uh
�w���ɛ��vR��6�S�p��1���1:�g���[!I�,؆�ݴ݁��;��4��K*58]�_�z,yP��yCT��G{,�m�Wl�S:@�����.T3�����C���}��� ���T_��`�L����(����'��y�A���,��TU�X��s���C���{m��r���������S	}���0.�����ǡ�װd�o��#[\�^��=��nE�Yh��D�0G7:��P��M��h�@1����C�B[ɥ(��k�䯱�|3W������r�[��C�j�E�g�7qN6��C�0EC�U}ֱ��Y#�Qp�ӈ(v�ZgrϐZ��I��Ɛ�o�y�򛨧�1{B���=>�|��r�i����F]o؟b���⁢q�RC�"��_��1i3FI�k<��z&���ط%S����iI�Dv]�e�;Ak��Eqਧm*��^Pa��FN�By��?v�.{��F��^gP٭��i�������)r���*|�S��Z��)F�-<p��F�Iڙ�O�w�S&�λ�=��s���4<�M�E0���ʷ)Ī9$)~�C��h�G�T	o�<���w`hLvC�?Թ���������'�}�0p��	wZ��e��E���wauS��o�Rw�.���c��b�.V���zd{�=E��@�st>�ѝO��X���e�$w$�͈Jv6g��Bpń{��n|3��2T��lb�M��L�ֿ�.����4V�8k��)��J�x���haӣ��W-h¦� ��Z3��; ��/ň�#����F&�h.��n�S�=���F�s�����8�5�V [@G��`:�Ms �e��=>y��'�J�2/�o���u���(������s[�n4� �h6A��FbZI�!'�o|"[�J��n���?d>�?19���z��3��DQ��}g��GdC�,��m9���Y�H��� ���v(�F^t\~����O�Z��mA��=Yx��	c��L�7%��1��d�c]�q�c7���}	������)eO�N�l�<b1dVl�p*�u��W���\W�y:�o�c�����ff�]�ߞv'�G����G�	��@���jZ�G|=��-��`�Ƶ��U�H��0*Q����Ύ�C�����	����~k���*�83�$n�ug�V�㜩Q�Kq�w�8���.z�T�//Z�� '�1 `�$��ǚYnݩ� ���u����"���T6�ln��˦��m�R�Z���E�n�t?�X���xx�p��J:��*�S4pt�.����8:'vdI��*}`$���/��V��*��M�3��5�ϐI��Aiۥ��_�}��(�J{c-�sܬO����XVy��F�_�ׯ�wD���Q���nM����c�p�i�y���B���8=̘�	`Z�}}�Azw)���j w�X7�[Q�h�����]��W�6�7�a^�0tS D!�Cs��J�stz��{��1o���|�+�kA�(w�����w�6��n=�����M��.Ȳ�80oM?�M��˺�b��%OV�W�R�ϸDs[CO�Z��f�QC\Ia���^�;�\���[�k����hF@���'�hb�щ�crx*��-���K�_���<�	"��E�����D��;:]~A�YZ2���5U �{R/l�Q�Қ���7�q�c�H�JBm�l�o�.t,��\�L����[Ѓ��h/W�T��y�Hj�ߛ�R�(�������Γ6��f�w�X�f�0��3�\��8r8k�ob�Pr}��� #��	�u��i�9m/��I�Q4O����n�u��sM�g�R�/z�K~�|t�C��曜a�yQ�ܗAx#�A�^>�l�Z�*�����Op(�U��zG1�8�2S�ӺS�,1���6.�o�N9��Mn�O��G�3[�y�ߎq[��~!�K��uJb*���+�;�?tR2_�����J���2۱������5��x�5	^	E�u�O�&���5�yj�_+R'l��\�$�F�z�66���t��E��V-@J����/T��u�a6q��|�V_:�<O
7�ܙZ��oZ�aK�K՟���Kӷ�/��7� #"=n+�#_�
?����)iiW��mkg@c�V5�u~߇�ÍH@P�%,���c�@��P��w������Z��=;��+�z��Բo�"'��B��{������`�*T��1��CiDso�>����pBޘ��[L��o_ٟu�����K(�b�%�n��e�r�.&`�}�wz�&���/���"߁Ԉ��ǭM|2��K�ր����#���I�n9Z<�ј����p�>}jH��Ý��Fz �J���F��q�@�Z��w��O0#�&�]��m�Mz�a*Wޅ�Hy/.��ᒳj�S�B����]럫}�`q�f
�Ӂ�y�&㝂���BI�[q>=���F�Lb����H���ꎳ�������m�����(v��:�%%��r��o����6 }��]��.�"N�ڐ��cRd%���3qP���$8A�R6�7��O���y�8l�=�K"	MT�D���.�%1_�W6Z����P�K��uSqڦ��o����5���`��K&��m�|����!�6���.9'�}	�R�(�<��XB�D�N��Q3s{u�_���d�	��C^�	2o�통(L�T�WOȐ�Qr��V,��������H��-�{vz*��]lq=�B��ó���̪b��E65�t�~S��cBeQ���;�m�,K��i��Z]���DV�����ָ�X´�+ަs:����;�<*V�7O��������f)���Ma3E*���ReD�y��|St�����W����Ɍ��@?yILG����ѡ��ɒ�9�:!�������0
�c�i�:��NR���*Z����I\���ګf$�ߦDT�KT���7՗n?�,�w��'�,��z��vh�n�d7"��
�W�|��� �9;i3jN�����݂�����Py���po���jô��02F�b����D�^�_z����)=%	Vxx;'	8��b#�t�k��2�Si�s���t3CG�^8��,0��:X(��������k�H4��Jh1���m�jc�L�ӽ��oJ�(��P��異¾Ш����|��:B��}����ko�mZ��.@���_㭎�G^�q2�M�����U�� ��)y��YY��/��1��jfxBe��u���#�A���9�(��? �m�~�׾�?�i8C�
m�b���\���Dpxs���I/ CO��/Y:`�;�o�}�Yy���h��D��W=���xQ��jd[���$��s3ly��!ӏ��!΢�VF�@���uTxmS�չF���&�0@�{��E�2Y"R��jِ��0CS�������u�0z.�`U�ߏKV��w�pj��+ǈ�ݳ��X��� �"5�P@,�N��]��Fz��� �cӏۻ�e�¡��}��ȉ��z�"@)ܔ�i�y�;!��6�!A�s�n�>)�������~xL����c5�Xn�':OO��U����*�(���~6� q�%�o�I�;��تT��{*���Y����'`�J3�3e���X��L6��k$��e��t4�qY�Y��d1H<#��S2��s��{/��w����*0p�Jx� ^�vܷF��:�q���˜�f��ى=JȉD|����qLH���x�����fV{E�gF���$�	1 g�8��Ӷ�rڠ��B�הכ�Tx�(Ɣ�;�?i��إ� S kM��"��b����~��60K8XS�c:#ɼU�{~�g TO�zO H�Lbd�ӴJ�v���=ܓ�j2aTZ�-?�^���e����T/������ߑ�#���V�����1�6��y�i��j-�0E�����Yb��c]P�0m��/W�@{�oF`^��:��$+m[ѿ�(a9�)���#�;����!�[r��"��=�t�֓��b)�D�oX�n��)��"��q��u��¿{@���;D�>��}����'a�E?�	�M|3��Ւ�C֨�p��HP��wݥbP��3 g���K.L�4�����F�P���7aj�F�p���8Q�,T*u�����{�U�"5�ޕ%V��e�mL���Ĩ�&��1�˺