��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ�!��1g �n��ȓF�u�ǂ�|�H�0(@�8���A��C��l>�5� ����a�U�����T2�c4NbRmM�$Xrx�L.��j��CgüSu9�6`Ap�H������� �;LKr#GZ�ػ��b�[40O�א@���c��'V"�v�*0�럛v)��/���XH�K;�	�x��ж���tB��Y�x+���u����d�e�f���ﺆ�$	6Eiﺿ�6R�j�(H�?�n�P5��f�YR�>،+(�'����!��_*�CR}Ւ=�����!��J�F�ZY�)X	�ty�"�~���-3)�$�Q�Q ������{y�@w꩔����:��D��K�w�"f��&9��H�c�t٦Nm>S4D"�Se�w�u���+���y��!0#k�7��c�I�PǴ��	W�[������ˇ? s��ϑ�d�!JԔ���4����o|��.�=�셨����+�f�al'����������{�9h�:eQ̻��%��]ݺ�POqvVa��؍�UL�&z�ΪA�T�8���?;���+<>.?�W�s6P��
=��Οn� ���lS�1�B+J���In҃=�	���?FU��%�)��Q����*�*��ݸ�U~�X�ޡԏ��_��!�sC2�;:��FI���e
������n����1Z�p�56g�Щ�i�W(;Ni0��@�`��WYW���/�E,� �BΥz>P�Z�G��8��&8ͥ��!�;Xo�2-��I:=Gp�$�E�SK6jm���R��%z��������jc�M���}�
Q$����;]����^�VCnc\��Є�o�=$���#��@���Ȥ]����Gl�*)����mA�ԧ�ʪl;�	��Z2״�l5;F �������.�Ǘ��}���&�d`�'����XY�"����m�8"��"�Ա�X����R�EQ��rzi2������B,:r�[��%��[�}t�*B�3���?�w�.��4�,~�3R��C��:M,|�Lm��W�Y����@aaF~��Tfx���a-G4���]p��Z��H�c�k�9�ϒ�$��%�cj��l���.�G����A�r]�M%$�J�u�QI��3
���\"J�o"[*`;~�2Pd>����p������R�
ɉMx�+H�B��?i��u����)���}z��t��>&��T
���T�M��.��c#Ipܾ�@��g�,##��خ��f$�{���.:�	�2>Vm����6��I3��N1O�ށ �ǟ��������4���\�R^n�Y�����
A�cl�4W���?��F��f�ٞ\�SN/h2�}q��7�W1SC���)�pN1�nqT�]ɖ�ȫ�o��=�g7�P-� LƩ�]+�L�������O�SOy#2�i&D���aP�����r�$]�m�SEX<���$��OhcD���{�i}Z�:3�G��)��T����#=���`_�:��H�Y��[onX����B�7A�W�������Ȁl���?݇��m�A&�IA�U\�a�!��_��P[/��OFId8��|-��!�^5�������ι��ś{� �e)7hڋ�b���6vh,��&�r�V)�i��2�h1��Y�=-�L%xqR}yE~T#�*v�W�m�+[�_�e8�j[����Z����+OB{k��{�$�L`Xx�e����0j7�:0J1�T�*ZB}�b�øKߗ`��ޠ#7�5�i�f�ɱY19|a\�۴/��@�AOx�d#�`�`L^A�u<�Um)����}K��;S�]��\���].��(/*��9��j����J�I�Cc7]�d��s��j�/U�I�|;uF���#��m���X��uh�]�KWKY�m��Ȏ�.�}K5���R��f_��ߠz�u�ZX n�k�>�B*�f��2Q�vv*�fq�ŗxޥ0n
[�$��L������:Cp�?�V.}��f6Ѹ@���m��u,��/�s���W6M}��Ot-384�e�u��GVۼ��;Q��Q�V���:&g�)˷�JK�J˷iD�� �3���Ak?O2D���;� Z�?f(i�����FA�E�؜����d�^�Υ�k�I:=JNo�p��y-������-ҟ�wn 'G�?h8e��R�|�3��^2���ҡ�}JS�}{[]I�W��ɒE�=*T�=���DxϬ�Y�EM�����P((��խ��=�90u뼒��޸��Z��>+�O��R.��s�0qv�n�~t�M�~*Z5H8]cf�	ֵ��)��4��a���≁�:�OI��&�)Gb���ot>���b���gx%�B��;o퐜G5]\��>�6��M��ծ.d8b(&1�
��[������k�����&}`簜#Q��a`��PLW5c���v}��?�]HdJ�������:}���jի�����˜��V��J���}N�_V��0����b��Q6<�ڦ,ݢ�67<�
!Q�7�v@3>�H��s)�z�M��2r8I
o���p��������wR~C�Oq��WB���wE�2cx�&���ʸ=I*��������N��}q��VC#�Q!>2f|QI�b�$�oe��M�7�6��bj��J�'w4��9J>&����+8K�ۀF�VS-d�<3��{3�!j�:o����kv�)d2��օq�k~z�];�5;&�p�sZ�aN��3p% K�ǧ~�,8�ֈ�=��ll�թ�9qT?1p\I�|��$T��]�9A�ॎ�n�3�g졪��NB2��m��h�:|������M�4�o�+2;�����4)��`+9�Щ��Bd��N8�`�i�V���/[��\�"!�K>@�qa����QO�gvH+?1Xp}�m��O+6|I�ge��U�[F
%Ȫu��LB�Y!�<:DPyZ;�o�k�!1\��;p���~����>�d�_��I�2��Q����V�/�*A��%����-d�A�]��)@���V|��ơ���k}T�n��v�vR��e(H�s�ߏ��z�Wu����qb�p�lA�P��q�X\nΝ��r�<׬�J��E��&��M������n���9~Ž��X����}�wL����昘�+��)�Ү��<��s�@��D{f�U�bZ)�O�7W3q�mD�ֈtb\z�g��Ʊ6!����J\�s�-��T]���nA7�o9��������������|إ�օl�ҳ<}F9�0ikPh|6�ҿ	�]�������XW#�!�T0!K���r������w�N���i!:���nf�I�Ӱ�y���5[7;���f];c��$��U0����U��0F:�»l��Vk�D�[4�n6�N���ٶk�Ql^Bԋj6 !��d��IIQN*���,Q�G��]g���-#�e���1�BS{���W)?-��h;
��G@F�h=7˸�B����=cp�MɌ�Ȼ��i�'m.�69a �Ǻ���p�8�p��i��J�̀������J��H7��K��wK�������JNY/�ś�������F4́.��I#�`�R�E@^w����K<��� �Ju��6��D��_�^҆�NM�Z!����K* �I2Q�D7��D���+���h?B��V�������tGGC������+��C�	ŝ|"�V�1;��½��r��� �|&�yGc���>~��R)�r���zq���9��o�g����v����ȿ�?��l�,8�b���=r)�L�Y-���Z�D\C<�%7�gT�	��9��ө+L}�ܽh�[��r�
'�տ|��uV��1霮��9h�6ˡ��KD�_�Ql+���M��/���vq�� ��rc�G��I��zt����2��R'����l��x���ú+�[u�4��&��Q���C%x|�<r�l��ra�A?�B������JC�~�P $j^�.���=�IN�<�+~Gnu�ؑ�O@ �9�:�&�E�~�ko����w���Ux�l�[�D؋o{�}ߙ�1��#�Z�����������!:F5�Ul���$x��T��d�X`���'*�z��dT �7�1��>ZW)�uI�
Q*&��0}RԯpsddU붲X6�;���b�ZZ��