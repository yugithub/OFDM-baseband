��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛQ���b��E��.(�4�5/�vNK�QT���Bl+ѽ<�@X�ҝ�>�v�&Y�_�?eX[$�%�û�u��YэQv%�N����?��֎�znƑl`��&�~Gk��	4m��|�+���(ݕ�ZYT�g\\1a"fsLQ BӘ�zR��X��4ط���N�g�Y7*ʽϬ;�^���eb�#�=��
�;�Rޠ[��n���o���i�7Ip��8k��'s	����'Zw��6�m�|��.Őbɒ������G��O�a�X��Y)k�1o�N�m�Dm�}���zL��Wn4��@��3|hx�p�u�*r~��Ccʸj���WPp�H��W���uX�ǽ�s߿C�#�������|�҉�(>ɄCaVS����7�9t��&B`�y��q�2J�PQ��^��D�Yatg����1(����h���2���ʰ��!�>�=�-0�O׬P�q��)��)�"�1l��䶦�ph�Ԡ�ͧ&�0�X�q&l�	������l�:�ٻ�-��I�W_v�>;�>e,���#����`�h���nbsנ&��EK��F{��r>��� �ԊP��Kvc�DOk h^�8��c�����l��|%J���7'+��y����σ�D+yxQa����0N9�ի�U���Ź.7Yj����Ў�d��H�7�?;�`���l�^(�%-����XA��ʐ�-@sN��D�5�U ��/'г��{�I��]�)i�%�F�`1@#&#E��UN��	3TƑn�c
%0&kټ�~Ff��"e���
�0�N���-eG<�m~�H�����!LWc���O.ϬP�(���Q��	�l��D��Q%%��^ĒH��R��Q��6�(�����`%5K�C�'!Q�E����*����N��2�n�Q��.@0�`���Aa-א����_����,����	:�f����Fb�m�ʖ?ew��dw���t���'(�k����v���pFM&�ˣ�u�D��.��Ɔ�ŶS������+�$�"���Cl�"]P�Ɠ��Na�D����ʬ�碯!����R�S�)�@3�[�UC��h.�h@��)�9��^��0�/�����b�AmAjk�[��x��a/�u��j$�4]R�8�Ϫ���N�o[�9Kz�oC�-W�U�|i���3@޼��sv�al=�e k�K��V����߼����)!���gŝ�6�T�o�����m�{rߋ6�)k�S9,a���2���Tr7>�pZ�<Cx��&�9�hQ4��;�����5[�h��o���h?�hM��7K�X-qX3�M��v������J�T�D䇢��V��f,@��&��{��w�K
V�O{Qxw������st��O����Fk�~+׏A�S�n�Rw�",��Q��(Y�p�?s�5�d��B ���e�&��]w���:4� �J�?7�*�	���RI��j���UB�{�;aM��}(���7r�b{�Ib�����S�`�4�����Y��R�mE���Jz���yȋ��	q�=΋����lYƗ�f���}p?91B��}㔻Xp���RD�dX�ğa�W�'����]�/#�WR^km&�Q�&@����M�̔�}v�x^��[u�@�?����˹�|�#�:��ʽ�+T�����Dj6zþ���0`��Hc�"^�O5E�@���l0V^P�. �MQ�?(�5��t��ΠF�_����#��_�B�H�?>Lk�i�洑 ���f�=R�Q�����s)(�m`�˸�7qޟ�	)�f���%�!�J�)����^Tut��3s��#�d|,����gL�o]쩐ͭP[#F��@�SZ���O/B�ES��,�3����n�K>�3ޖ�W�[�t�Ip;�XW_����G�C_���N��c|���#��	�	e*�,A�'y�7
��ޠ�;3�[����u�4���3�e���t��Laq@�S1d�3�L���T+҂r��A� iwa˵��\�%t�U����UP웜N�|=�<}y+�D$n���:E��܌��l��p��9G�m�v;�3��ؼ��
\��m�n�c�h|y,*w}����3F'�S�4�w���Ib��Ql7��*巷/Ik�#��<.3�yC�-A���V���;���f�>��􋱑9��}�uE�@nB;������5]>[�-�����Bzz��EMD9��gT�f������*����S�tQ�>/it �H��(�&����	���K�u�{���_���Rq;�N;��X�=B0� �O�}CR��#`|���|�Y>�Ĥs'�N���_C�~��*}@�6��P]He��=�E��t���ڔ-SbS7Nܷ�(S��5�cޛyۀ�N����Ds��t�5�q����xvY�r�:G�L0����h�����ٶ��L��!��y��% Qa!�)����ˋ
��'(�	̤�`	��ӎ"��rj�Sm�å��.�PE�L��#Q�#4�px��9T0e��1���Ỿ?|z���8�D\)S7bڻ����V��k؊"w��O���"�I^�[��d��K�6%N����P(;& A��-�Ţ�����̅]�H�&oS2#e�(���[l� �@�=bF_�&�հ�=HZgȹ��R��z��u0V7�J~�7l��[e|�19���e=d{�����՜��FC�8o�BS�$\
MTq�L��_��St9Z#h��t�X��v�7�M�\z��C��#[�5��x̏q�'QEvꞿ��`����X|�X{�Ū��[�.����t�x�&L�����g�H��"�[�ގ^�3��Z�ⷍ_g�����n�8��4�B�o���z�L����;���I�ܰ�X�w�Pa_0(��u�k�@��L���N̫[{�dafj.��2�a^-������7ELY d�Z_���QN���f��k ��/�S�c[�b�y�,�hK�v�x`�_����ٟ�q:�����2�絣<��!1�B�Y,d��V��!��N�V���m�	¥�{@/�}:����9tL٪�s����;��K̠����2m ��+�"xy�Y���%���@R2�$
>o����N�^�y�I�ƀb -�Ia��k�F��v��%�����!aC��|�xÝn,N'0��M��I��[(��.
�zɰ�V=2��?����?�ȴ����<��g<�Jy�v�-c�P�Nq���X�X$�!��2��啐�'q����
�e`���L~��z�=V}�D����&�A{ �K��f�.^�e��&��kP�T���!e�y|��vĽ�9o�u������������k8\p;?r�/C���G�<r%~�R:u��2�!�� ZT^$�e���z�^�������E1����i�P����$�5y�s7#��Zr�"���v�C�`��"��+���י6�O̘\@��s]h�"j��HdC��_dG�޲�-���'o����Ƶc�	ۑ%�ˁ�{�"�{�Yଂ�+ &�:����j�Q�qԋ��u����kn8����ꉳ_����v�&��`SS�Zq�(eؾ�r�h9s*��ښ��k������8���f�7��$�Y�Nʷ8Λ��&�RA��gI+�ɡ�X�6H�σ�D�@�ލ����rpGXH�]���Q|A�"iS�B* �2�B,?\:!G��.2 ���U�%b
����!�^H&�~�Sr��aw�k��+����	��q�`��:�@��&�`s*Β��ͱ��(_n>cB6�������Q��_��j��Wv���k��Ep���i��E@�]
.��#(�*�L����?�(\3{:ss�N�(t�)�,L7�j���8z 
�XS�^�u������t��;�g>=S������K
���Kvf���ʑd�����C��ܺ)8|~pz��0����^:�L!?�$.SD���a��ցn�y�Sm��d�h�/q���Hձ���lf��9�+�`~�.�� j(���7G��"�8����۝Hr��ێ5,��P�i1�tX\	���7�Ҏ� ���bk\1V���!�7�A� S���Wa�-d����qT* ���8�t�|8g�>���o�/i�.��7�������!j�_9
����6#%��x�[�/*Y���5'�*�lh5�35�MX7~�X!k���;'�)�z^!�����<ؾ�ܣlW�[�LG�Ā��|Ar"����,�i��%�p��K�D�{�7��&�n<��1��-�l� ��`xD�#i�6!ڂ?�;��M!g
⎤s�{��1#(h�w�?L:Z�uh65X��n�������a�x�h�(.���{jk��c��1㯠���!���Qe���_\Z"C�~�1���la��{^�ڻ�'���i�o�P�<r�kC����Zo,�����N�2O(�YA�k�S��(��9x�g͈'�F�d>xb?w���\�I�@�����68�R�)���!���!j�:FS��]A���R(uZ�@��01�&��Gq�I�+SPH���&h���L�*�me|�j�F�e9�|ҳ���_2����*��J���*��b�z�E�1^;��5j�ȜC+]P�6n�Ŏot��:��a�/� ��?J�?�lԂ�3f���a����� +�4̉��Q�K�BPT�sW�᷵�_����o��z�7���yr ����H�~]�d4C4�jd��B<��%�Q?�6��t����(8@%�����*�|6�~�\OB��|���L��GS��h$�@2K>h$Q�\!e����t�����@���m�΃��v_�]y/�2#�3W�[�[����.A_�Ί�sm�����X1{��ɒ����(���;ab ��H��G>�R�l��$*�	-s��ud�ʘ�~Ч���:�I3|�?�
�]���js�~+����M��tO�]�Yt���¡ϐ�y���Zʹ���R��5����3'/*.�2��Q�pkW��TY��};x+�Xh�\RT|�B���o������,���R?�nX��P90I�f~y�-̢tˈ*d{�	(��a��t5�����h�W0
�zzH&^�t3���YÓO��6����W],V�G&�)���P"�
�֓�>�3�T|
O���}d�.�e� �(�M�PX�! d#$35��ʍ&T����GOo���c]��vOˬ#HC�h{���>��3<U@�!w��8�
�$�Q@���Ѭ"pݞ���^���<���aP+q+�_~D(	�!�cp1�;�o�\p�(?�G��1��� f�����I��I��܌z���R�6u�h	��]E�w���C����q��h���&��mK�_nd9��{X�ѼϘ�M8_��܂����4hB�|�n�kT�b��N�ّo�	��K�y�tFp�O�s��8K7-uH��n�~x�:�Ւ��|���~:��`�(�B)@�n�`���P�UGg��-v"��h�zi�*^��\+t��F�$�l���+,_v)�izN�9C��y�i�E
6���Ghj磣�ə��fͤs&�n5�3�P��'1;�4|>&��<g�ug�i]�ɝ���'9�&��>���D��<4���VE�A���w�a8����Ki[>�lּRO��NF��ou�8sVHb%l�'����f���76�Y�Ke���Z����ōr��#
��.�I�����M�T�I��:D(f�\'�F4���5�߯�����g��GԸ�''n�}w��O�-G�s��n��fEmt�r�r��܂��]����1�qDiFwAD�S�NtJYL2Ji�$ah��us�~;O
Ί����N@C���{�	I5}���Z���2����ע�kOrx(n����Z�����ߓGxj��s���'˿������p���� G6I��M$��0�K=�jLC��՜���"ӊr��QAp����t��� 2r���L)u�j>z�����ALI���.p��0Α3O���^4�B��vH����32��lЎ����E5v��?M���w��si?�L��ΨG�$���?���!�N[��2מ��d�a���|�p��RA*I�U�UK�3e����P���Wi�'���Y	.bf�����&�� �)ST�F��w�!![�Τف��/r�v�|�\�j��DG��~���	f�~Rk*�o�7��	����@��VCCe/��=�r�=D-��.[`Чsஹ���_z}XQXش��D8��2�bk 4���N�+���ss M�����D�����Ld��-yHv�ߐ��S�
�$�v�S�pW]_�F�|p�2�Ѿ%�:��|d��w#ƀ�����-$J���?�g�Zi���p�`:��U��J�L��v#z�OTf'��xMf���4��M9L��k�����`t���� ۨ��ʬ��x�ӡ\���:��Mx,�c l������e�&���)��̚�z$�Y����qo����I�w���,3!}��\c�tu�k�QV�ݣ�*����<����{(��T������vIy	�	b"�^"=�v�Iwb�Uw�6ta���	�g����Tn_ޤ�����P�#�@}P�جcZ9��X�S�i��"���������W��p:������	š�%l���|x?￫-zϤ�
��YT�@����V7��K�2�pFg$�ݕB�h������a�w}ޜ���Ll��Nķ $�	����KR��i�7^��͡��s��Q@�w�_z.FH�ӐPT=0
0��0���Oxl���-�-w��'���K�X�f�����4�9�SƇ�n'J�4 o:��� �
������J�8��
�	}��f� �l�����<�J�嬠v���;=�!վ�9�� ���{�n�-��)Ϳ���x����l�U����e3
ZTO��;���� N���'��R%�sy�{7�����HM	G~�fB�b>@�*��`��\���T�I5�Ȑ0f�zM ���L
��0I!�u˷�>yP������!�����:�����R�b����`�+�M����<LD�����~ żW02�3�1]{>ߏE��_�z����;JřQl�Ph�%�����;8�"�G�hG]{��*�R�e��j,_i��(�6�hG�r��˨����Hڲ���P��T�[�&�{�Ξ�Hx)�n��D�koگ��k2ۜG���܌�(~������$V��7k���V�~Ò8���i�AF�'��s��T�L���g��5f0#������SE=�;�\�sm{��	Q�w?	5����*�k�a����I�'���AV0�����d2�8~x���&b��q�;U���Xsg��X���NAs�1ك�P�'q���pu����u�y@�N��?s۽`��K�x$a_D���۠��TF���2���yQ������������	S�oMq�]S��� >�"Ҕ��9u#���f�u�_bt�V#�JJv��穭�� hqS)P5������c:)�r��ċq~�4R��Vؗ�pe$ws�$tz�T
s��<Vh/�� �O�����	kA^(b9	{�T���tg&���y&��`����1�Q��d�`o��8�n{���ԡ��D�Of�iH��mH��:�]5F?�L�����2 �ƙqR?�;�Ҹyx�Bi&kTj?�[Yu�M�"�(4&�?�5�� 5t8�\�Ԛa��GCb�Y�:��]W5�|�nw��hh�'��p �����N��$j��y��s`�X��7g�����g���=硥4zP(���\YfܱF;�z8�ړH+<2~����0x���h�CB�<Bn�7?G�����+,Q��dzC~r����0n�����5�P�]A�~ES��\[��$�D }#]=��8A.�j�v?��_7Z�����B0�zKR%��O�����#-�w������B�W#]����{�|���@����W4���n�Zќʬ�}x�m��E���A䞤\JU���׸�Tv=	��W��mĨ�m~���\�!���0+_�v�J���n�P�n�F���x�O aWO��E�k�$�,���� U*��3��1���X��G�XE��8J��gn����Z���l|��Ӿi��NGK��{�2�/l��'l9���$�}�y�b�7�Y��
u�ͅZ�T+9���RF/�I�����{>`�G�Ǧ!�����횼�+j(��q�kQ�ݫ��N�M�v)lzKΒ�u׉���4nٜ	�x8ظE��	P���!ᔩG����j�ea6��ySH���$7�X��f~� �>�ҟ�����s��3��O\fm�@ �l{�cXĄܥ�?�G��Q�,K�`kވ�������r�p	� |����Cg�J8R�'�9	���;(�\�DK?�}(�C��t�4� B�����>���ܲ���l�ž/��,��-^H��%a�CM���ޗ�MfC�h}�6?����Q9d� ���.�
�'�.Q�nxC����Ŀ�Z	hH!�[�e��3i�U_���7ӝ�~j��N�A�0�{zɊXn7[2�l�P����Z��<��Ҋ�n��E�c�$����L����c�-��:�����	��rI���R�𜏳E P�u�}�>VÎ���$�y������w�;���Ď{b}���}�g�U��:�8���9���/��F�����hV��U��yN��?U��"LBKl㤾?�yr�o"�Ҡ�^�SEq�,������z�g;���&E)��C�"Z)ph����IZQ�bsI�6��7ì=���G��Ha�|2b���Q��':�K���^~�*�W������S�'�!!$zu%MN2�b�*��e����C���`�.�	O�n��`B��:U9�&ݫ!5{�NE=��ݪ�0�g@�wǣ�,U��r����$��(��:0��l�^[ʕ�?�R2�'at�.jA���w�F��g���q��uф���i��@��_Wmv���J@�N�q����Eވ�`�*��(5�;�_`zL�(������s��� ���� �g��z��E�f�zSe;!pO�|R�"���y*�����.FxN�m�QP~d���)��~h"+ǩTB\ ��n���UCB��c�Rs�0��X��MqZ��ICK���o��'L�ل�E��U $&�N~�f�[�[lݓ���L���P�=ʲ���=>�d^�q	|cܵ�����*�x�|w�=�%���G��")����l�[��H �>���f�˾y�M�|JQ����`Y]c<IԅD��4%Bj����õk����{���6z��I5՚�L�N9[�@��+��:1my�vW�1n�$h"uB��V������V�U)�4H���G�Iֲn�V�8�+�lp��=Ξ���g`���{��6�>�5{)c�Զ�&�ř��W?�_)vh��)zP����HT�&4�7W���zF�{ЪX	u�\����-Axb�J� �<L�SmL��wIЋ?R�l.��/��DV��W�xA�F*p6�T�h$@e2����;2H=X�#䠅:&�de�.��F�<4��}!��_+�-� *�#ed�N}¼�E;��Y�Y2��2�J�x���hPl%D�%�E>��������KmR)a����Z{�օ2HϕEK�F�5#�q�}�]P��*�g��@I�۸�T�Ȇ0p.Y�����o2�s�[��q%��c�jYJh��;�J�H0/��Ʃz$r�h�<�W�i��D�B��M��(I� �̯~�����S��3N��@z�1���3:��>z�DN�����>e�)ɞT<��o�������p�_'cDQ9��c��}�N��i��|o�[t�v�d�¯Cu����̋lE����� �c�3���Ŭ��I]��6��O��9h����Lnyu�7������e����i�ǜl���3�QU��&�f�<��f&�l��Z�|�}�������g�Vе�i(�l������
�~�83?,l8Ar��V�=�!y��Xfǽ�l��H�r.*�B�[�cհ��X��)#�Y�y3�����^�`g�ե�Gb!YP%o�	=ɡP��ga�i���Æ[xn,������-�Ԡ��=L���f&�%N���:3������X,�Q���jܷO�~�:%�E
9�;�FC�n�0x:�ϨGvU=�B9M�-BlI���	l(�Nw`�����}�N���tB�e3�e`���ti?5�ySΡ-�a�� �B�A��}�~2m�E������!ՙ����V��^z��aJM���e�%��+�bZ�M�KQ�����s�����o�ᵜvȊ������J�+����Bݢ��O?�э�
s
բR'RRs[l���.��;�/<����;D�$p 0d=Cio]��D8}ط͎gO��J��M��������X�|���(Sa��ޱ�b�=��L�l���I���՛����4��U`5��v�S��$h"�%��,�(S��a*H���Oª1A���z��όxU�v��i<w��l�<��]i�~4�ϽK׀�*ʔ��������������*�Z���|��ҘiE/h�񤑷�߿1W���`�����r����[��c
�A�0��;������	uۨ���\�q޸�3����������-�[����C�;k����Q��D~����e�X�NȀ���p[Lk]3�U�0�F(ѹ���i�����q�Mu�S~Z�	7B�<Y��l�-�%���Eh=����US�Zh�cd��a���� �x)^�3�2�⼻9"SG��9$��"�H	�3���>7��n�Bf�����N�y=G�4���(�E�[��/�x��n����Ъ��
Č&}IAx��-�`u�r���E�ݔ���·[Ǚ��W�Q�
Q�s��J����m�H���u��KZ�OԉE���2	0#��םª=��M�`ּx���I