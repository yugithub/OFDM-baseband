��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ���6'��Y�8ֺ�L��|sqwɦ~�b�̼ީ{>I�󠗂+���֒���*V�'�A�t����w�)��#ƶ.RS��)�g�k���~�X;G`A���.�BԼ޲�CĄf�S�#����߰��&�U�u6i�#*P#�O�j���\�Gbv�w�ʖ=%m_W;�u�g�Xr���ġ>��+@��MG/��fDVA�Rx�+�
: G65
)2�}(�JS�?�L����l�G}v31S�y-5�?^7?�sri��s��V����Fmi#��
\)�9�kr�LFE-�X�d��wK�22Mn��?;2�zg�k�&�X�OY��r�)-h��l�]`�u}�̊��2_x��W��8p��?��K�B5���N���8|�(h�A2�!��{���a���=��Z��`�Z]WdlS�_>H�>��n`o^��h���-f!<1��.!F���#s�� ���8���.Ê����j�"�.��ܔΑf'=_���-l�=�#ǭ���c��<I�cl�H�PC��ɋ�A�BT_\FO��8ͥɻ@Hod��-��)�Ⱥa�<��,?$��5-��&���V�¶.�f�X$�O�m0l���?f�N٠�ω|[��9�Ne�-��E�q�Z�LѸ�љ �L��H��G�<�	~���Q�1�[漻��h���'��;����z��qB������j#0Ԭ���nܨE����r��x8�ko���k�	*#O#$� C�)?������'��Mu엾���F�	���M�\^��(+����Jx���O���пq��C��h���Xc�%c�T��_��`6���k�M|�`N��Z� "<�gJS�q�V�Y1������<���J@)J��
/��ᚒ%���A�a��j9?UQK'D޻�hY��O��l��Ҡ_�h�Δ��%�}� VC�Եy��)њ�c�yͷ ���k��v
}�:؂q�x�O�D�g�cj�MА����Wr�@
�N����� ��Wt��<���@j{���FX�#�{���š�Nl3NҙP��q����������U���X��|Q��hi�:���=�?�YV��䣎����$&��q� ���cG�NLM�l	?gt&ʎļƧ�M�==7�svW���cZ�tBz%ɷO�K��R�;J����Ր��ײ��z4�U3���Q�B�a4��P-��>�U�TԮ@�G�"&*;JR��s�P%j�;����q�R���C��(���uB����C��~����
��w�Tg��]����R�Igg_Pp6��:���'�!*��Ϋ�����;}�k�?(�r�tq&�p�7
#-�����b2;�vZ��g��?���v�7��v�K[�):�}Ϭ��>cg@T��j)����}Dx<\��Վ=eZ�-Z�/Vrb���r�w�Vgkx��%j?xQP��"z�ï$�Ϲ}e1�M/��p�E�h�`��)@��7�0Qv�����0��n�n�$[}���0�����%�^���_�����������}(��Wc~x$��H�"W;\>!��>�8]�R=i�k��"�,7�����d=�n<�Zԙr�?�D=_GK���j������4{�;��^E�m4����H���W��x{���{kH���"�*��>MSgbr,ʟS�Q9I��4¸#s�iΤ�-R@pn+ q��(U�-�tRRS�w��w�^Մ����Ni��^�ţ����L�nuwLܮ._��'�#:�H��G>X*aGA8�fn�2HA��*�#�3c��ӋB!��㹶b��{?���E�$��ȿjE:��C���S!͋V�����|�;�уy��
j�g�ˢ��XVe�#�ꀵ�b��𣇶?+���D�~&J��m�{|�|�@����}����}�!|�9��|D��)u�ݫ��#�E@���\_���%�ն�����O�4FG�����|D�r�\@�n����b=c.���Wخ���E{���$�` Ls�ahN
hz[|Ƨ-�O�5����-�R��Z�����.���%��f�F��m�Я8��*,�'�'���Y^1�+�%���ѬG- �8C�+����[�ˉ:!�dJ}�'�.g�W]OF��T�C
��m8��M��\��6�����Dr���3IB��������ʘD|� &��R��螷IqŪ���Z#&Ǜ��S�=jB&O"o����ˌ+AVyZ}} L�����m����!hP	�Km5���mW�1�ȉ��L?��\<t:�4����Mluw9Bu�)|.��mDha�4AH����u&79M$U� ���j6��p�hq������gNB���"9"�-�-X��H�;�pç��3d5�c�'��WJ��/N�8ub��wd8��m�M��m���"�Ԍ��`�w�B ]�1�Z@�G�h����9[������b��3z@�]OR}(;����zb�7���?K�̑�*�78S�eZz���J�Y����h9i���B�[6�Ŧ���+c⥑|MS$�o��#^㹝"A&�@&���+˒��&`|��z��`�=�ٮQ�����xcږE���`W�b3m�)Q�\oH,JV|5j:>��s̱^�9�f ����ab_��2A~OMY�K�D=j�M�����z
�Py����3�w^aM]`��Ks!5�#�+H������� o!�T&�T�+>��\��}b�H�Ƶ���o��,���3��`��Q�~�Mi��<��{���T�ӧc)1h���k&����_XwQ)�ÿ��2u����A��[�"��G�z��
�QӰx�K2���},���Շ痙��\>�Fۋkb
��o�����6����i��݈�K R�~����_�SJo�I����OD[�vy����1�_	~��Bڟ:a�o_fd=T њԢ�/���) w�ې�X�[]�XM�b��m�^+�mcI���~�E�|�Y�?=1�a�g���J�2��ᄑ� �	��n���j<�[�e��[�|�p�����i���; �֕Av` ٺ�z�w��	�u8?ݕ,��m�*���y��}	����g�s��[��Z_v������U�  ��0���)�3<�T6� f�c:��$).�J�m;d�S�(���o:lW�f����*���-Q8O���F�%�?+������ �Λ�+!�ӥ�؏ʏ�N�16���P�2�PρN]dW�I֜冋ň��f&y��Ή
���'02B�),K(tu0�y�����/l����M�┣IV�`���E�OY��[������b��FY�n�
_��G+�ƒ�#�=ī���frToˎ(�"��P��w'GA�NP���z�����V�����'7��2�����(�ǎ��A坅턉��٨��ķ����/�*"#��M[��R<�V�2���F]؂�'���y��+�����f�U�HCc�>�+�`�ۅzXxTr����Q��/�Rgfh�2�����B�'��*�:پ���a���ȇ���>{zzpk��ϥE>������^�zs�� ����}��v~�mr�Y���p�Ӭu�s�7�2���rrg���\d�xcgs~�w4��ͺ:%"�ƒ���s��7��w[n���qx �6�}����?Q�HhC��[�"y�z��c!M�'.00*ؽ�:����6t���z��on��W�ū�ܾ#|�����;���`��TwM��na|�|'uC��&#�q"&P�Iu��q�ϓ�a��X�E�:��E]Y��Q�x�lJ\��MZUxy�c2�8��h���Ў�}�$��xt�̫_�G���C��T�g��Z͢F��`���*�ߘ�J'=2�=��J�L#V�:��mp�n��IY~%�`�Q8A0�l$�.�F.l���q�;�k=�Ҳ�,X �ģ/+�������?Ip&�7�ª���/9y��F�7
a�դ"za��c)e�5 ���S�x'8c3���Zŀ��upz���?�S�#��(}��nէp^����ɑX:�MH��i�W��d�؏��W��/XT
�QQ+^��ĸf��"�Z��E����C�09��q�.wk�@�m�3_�
{^�<��93�T�!��*�+������*_�СO�x�љ�{��U{ʳ\ߤ�#��)��b`Ak|�R�.���&c��u�;��4��2��|i1�������I,E��
�(-��*�r^��`̅��ie<�d�H݂ ��C�"e���ssd7��,��蟟�-'�b��|���R�Ho�H�AQ>%)a�֮��$��8X~��%��Ҁ����±GG���/��̵'[��^ӭ	��nЧ� �W�L��;�j���(!�K������C0ja����uMH>�t�w��hL��Zƻ�S��]+��	�z3u�[��$H/�h0��~����XI�����k�hZ���x�����w ��L�&�=����ȕ��y8��G�؂��w_����b�R���4�����	�yI�A$�%��xN���#<��e�7��'Ph<œ9W������'{I��)�F�Y���)�s�.�7�O�9���m�,	On�U�8ǩT2������hw��'�I}L��W�t�̥|3��;̸�h�j3�������������٬���]��@'2�p����4�_#ֵ8����DtǾ�
��'+�
�޸������FT�4!�n��&�����k�r!H��Id�M�"��)���O@6�]}����m���Qb�|��8g-��lnw�ߤ**[SZ����ؤ��~s�1��v_
v�U~J�4��M��}�R��$-#��%����w��%�3gRT6�����GI���ׄf�)��SF�+:�E�&� q������u,������ Y}`�����%����j�O���B$�˧XV����
���2o��~��8��b3�}K��`~dʻ�H�&�O��.����8/kC)@m�S�:+17 (�i�E�^���5ʛ|�dl�b��1��Y��Bwy�G���y�"(�2��3�wCE&��)�%bv|B�to"�m����������9������0����=�g�&H"ny��锛+�	�Vl���Bօ�E�DS�R��'�0��5z�^�k���mf$�%����b����{�C��<���1�a����v��-�}�\�6I7-�M�ŏ5�0�,[&�c��QV��,&3/�ڪ�m]��l����3�B$l��^b[����;��_����z�!IrD���|�n��{���Q��t���I�k�m�`F:2��i4�iG�m^����u� X�5aM�D�Uy�g�x�M�P՗p�i���丫�q����Pq��c��~�#���Yރt0t�u�y�H�0[n��l	�o��^fǊ�,rr��DWn$��Ѷ�;sM�ݎ�b��R,K���!�����t� 8v��1	K�� �V��N���Iŝ ���J��E�,��Yi�'S1��=s��J$��@k��--��h�8h��<��k�ʣT�mH���u $y���+����] ^ě�>���B�>d�<���g~�Z���-H�������BGN2��X��e{�.u4�]�Z��Q��I�vC����99��J�g?B��-�
�|7
�8�	j��"�Z4QC�ע:�Y��7nҨ@$y!c��@�Q7��МZ������9�K�:�0Z�N7���޴~�4�M�2����� ȣ�s��/�n^(��� ��k�y�)�4���+�����B4�䉍)t�*r���
.3�veVL;�o���[g���¸8�r@h`�40cjT8,Qg5�}������.x�=ba�C=H�Nt ��禅�hE>c[�j@\�.���t{�v(tKY�Vgj�;����)�/��-;��_�3�e�p��1��}��:Q�"9�7�bA]f���(��Xv�dϤ3�xw���;�������q�V#�?^��O5$���R�2A�m��ɛ��2x�2�қ[�%�� ���s}�iB�á6���lhŷZ2�/���h% ��9�y��w�~������ ��=g`Ȋ�n՗�0z	��� �P6���g�r9Q5�sWn`
�^G;l��w}�a�˞�­_�8x�/�I �����Խ���M������4J%?&$	������,��&<����.���F߾��o;�]�[��C�9�*qe��c=6�y�HQ���n1-4P٪��K�� �	A��	#d�u�Ji�ْ��ӧu���qI׮e��i/��J�Y��l�I����*Bi�e���@��h��MОw)ohP�
^8f��ԞS'�<�}�sh�
!�4�V�Gb�5�i��J���Q�ށ�5�F�K��Q��L���	'�aLq��V� ���+�9(Pz.b%ӣe��H|�opp�j�X�\ �&֫#c��hvP���R���Ƃ�Wι�Ʉ�kA�E��)�E иN��f��k�n��R҆���R_��A�:��5ąD�J���(�IxH�?2��q��ԏ��=xe��(+��U|�
Τ�-���vDJ��U���8$%�f	T���}�Á����~�{�̅w�v�-O�Z���_*�ߍ{t���y�G�*!J����
�|!
��F~*V5,��/������u}�s�f��uY�q8�{�5�_��M���G?ë%폭jV8
��(�s=��{�3i!�����gG�VL�)�3������D��[��oV�\��G�"�&��sJ�O��k���:���<�y�4���A{���`c3w�F1}�_�m�p��{k*}�K����ڴ�p�[;��uF�*V���O`}F�+Shf�]��7I!���Ҿ@�d�F�ܵgsF���Oܑ�*�[��e5'�ϝ��`l�a���]�<������wZO~��3��m�i 4�3���7Q��Q��;���[i1!Y�o���z��9�lR~M=Q�D�ƻ������u�ml}��%���T��+za=KAV��>%>5��F�N,�D�#n-wM�Y2��V<�^�N���X�wn��������۞�!�(�)��D�<�Y;(�NYSJ��50D�)�*�n��W�:��*t&6�l\b� �6��ԋ�H���n4���(�p�Ho`�/�Q�tvK�-��!����T�q'`(C���tnQ�ye����ʔ6^A\0jRK��eт_���FB�L�l̝o����� �瑷Xb}j�,�S��8�C%5�yԱ�$B�!��?JZ���;|�΀Q["���j�ByK�	�3���H�Z`����H]XۣX�!�Fo��{��k�����9�VƠ~%ّmh��ճ�/�[����s�칉�Œl��Jd�Ed盋ut����Q�<�pPo2e<ځǈ��r�O�_�w~B�:�^Գ��Y@A��3�Ea3Gˣ��ƆlL����=���
�t���=��z�~O*��f໾���su"�ڰ�3k�[ ��٘iϜ�w�B&��"�2�^�,1�aЗ���Zќ�.E��{"�\	�7�������f~��o{��L��J��,��n��p���C����F>~W��8��KQ�PYa�l�SXd���gSdc5��NDb$$���n�	ʩG�=��.b&�ҸU���*
�`�Ռ>�ƻ=V�3l[m-O0��q��x�LI���<-!�u�T��s�~F���Q43����|�c�.�٨7�X��_1�p�h�8C��P	�Z�	I���ٕ��;� � p�a:i��۩�h�o}�:�{��a��w���{c�_��\X��Uy��i�����V��]-��o��N��i@H���{�Co��m�"I橠���sU(e���"ɱ��^
w���e͖W����~�~�3y�+,K�&��-�󙦌�.�<���-�.͙�w�4���N��8'45VIݰ"2�ۊC�mf�M� ��S�<4�ˡ�!�Q9&�Fhԉ��]V���~���l=㔺��h ��pYs�<$�7�'ac	�#�,�m<�+Z�NB�=x���$8�p���}��7l����� qt�q��$Úr|#D%Ƭ�J,��9t�D1�4��3_|���AZ�ڟ��[���A �&Szc�l|�[�$[�O{6�v�^��]-+�$a��-�{ŵK�1��ANe��8�u�w��;k���X:�53��/K����(6���B<�W}҄B�\0b��y&�$zڀ4Zj��f�K<�y*J��F��B����N�q/�w��ÝH���H���1>��?��1?�p��{����ɵ�i؅N+��tr�Ŕ��5�LA�� .\HN=iN��P�Y�� w�*ܶ��T�<���y�1���[f�v�������V������z֐(
���1��_>$XiM>k���ڮ���v�Ņ$禉�U���V�9?�E���H�"{i����J}�.�{ r#$]B�X�G�4 �7z���L"��/��zD%�=��ŖD���Z�Á�Ԧ�,��4""��JmF�Ķ�0�*�8�J�|���D]���W�6�?O|����0��fk9�}W�Ǽ(ˌ���y�F!����5nǯ��/�+�&�G�@mo��U��W~��:B��v�uS�b�S��hJ�*j�fD�8�?c����3i����[�!�WD
{����
����=$ԜV5!��L��7�ڽZW�9���ַ�[�̿��o��]j ��v� ��2��)�fw��$M˼��C"��G���t�.K@~��G�o!t�WJ