��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q�SOj
[��%�F� I��F��Ul�Q�(�F.�ՁZGL��	pHDJ�ȷ6������s����<)y3`�]\�G�:��u�փr�&�����:Cb�#ޡ$<��\|��t숶Ų���0']�t�z��7�g(�R3'v� �U��	�_Y3�.(���W�K��=�h}�%2���y�y�-T��d�f��A�J��T��ێ=�s�,����qm�Q�cK���� AƮ��ph=�p�y�h�ϚN?���Sb�_c̡u��u򜱢��޶""?�b���,�Z�1M.6�0�b���t���Q� ��|�9\1#b<�	؃
����L�w�U�*՗z��q̻*����&VW�����i��B���A0�wL�sH� ��j�])t��;i��S�YA5FMNx\�K+��M��;◪wni 
��Wi�K�Q����(�I+���NŁ�����4̌��*��%��$рE]|��A��R��Ձ:��Fe�M��]Xx\F�q�����-T �����;ּꌾ���c�l�33(7@�=�����
�)��w�$J�Em_9d���D���7�N>���EQ�����;�t��K�¤X�!n�fp@���u�i���J���Cn�r��~�_�ރ=��x/V���3�%ZA�X��;I��rA�@��F�ѐ�#w�:���N����{�53��E"�!S��i�Q����ӡ�
օ�j)'��ݴ��ZFǀ�'$.M�O����D��h�%d*0�6�c��e0��캾/y���N/G)���}�@g�~9��ʇi�7:�G?�oM�+a�a��M�������A�ق��p���<�ϭM�b���s|i���#�(*rwNJ��MM1 ��R\������%`���>�l��7Wמ q-�dn�9���&Xچ�0��8���~��e�:?aq��E�[I�8�p��;�����T��Z�-��:uT,���;��!G�H��:��Y��p5g�M�������ʞr��S����oV�m�w����30c{��G�a�Q��㕵�%�K�����,q.��Y#H^iF���)- ��R%0��pƪ.�ߺ݂�"�PϘm��hM3�b�R����[SQ)B�Z�Ca�ؒ`"�3�042\_��i������]�9�>���$�駿a���in�k���e�ߧ�P�,����
}[ݸ��k�A+I�>����H�/[�w����#�Ob0UDy��b����Q,q �=�#(6 6�3(bH�?�k7��Q�,5����=�?��k���2�ko����[�a���<Մ=��z��ei�k��Øy�Y�z@���u�o���8�qɛ��|��ć�`;ϲǑr��W�
�7doV���w��A���p�Q$	�AK�zn�3e(��$Ԉ���/���Nu��{M6��2�:��C& D�����`��6�*��,*��E7�.G��j>`(Z����^s��ֵ�-���+��ڸ�%H�Ѐ^�F�Ėm<h.��s�WeY��kI���#؄Z�
��Xn�3}$P��\��5oY��R([	+�Rr�=��*�c��(��k8����{%#o�	1\��6��m*��v���1�4BՓ_=OdRz����h������n�.q�},>p�$!sy���do�Z��%A�QyJwq٬Ŕ``�ٴ��3�+}��V<��k�x'W����1V#~�a�J<ќ�}�d��8�r�ԅ�����A�Wxd��Ƭ	���4.�pQTd�"G�������W���w0����O�n�:u�J�QZ��=�Ԍ[r��0d�7����0���B�_���d�7�!�E*���j�c�۽�Fşs'(q?�~<�*��/�XAa�<��mMf�M��,du�b��|��t��KPj�F�	4U�l1=h<")L�\�"���ϱJ$�x%�}Q�	+��49).b�ж��8�L����-&�zP *O�{�ʲ10n�Oj� �`QLB���ش%M?�M9��P�]e�{�;Td�~�A0/���h�:�f���H���,�½��w�ҿpw괷JWP�;����8�o7�&I�|?�<�}�-_n�V����e7� ��x�s~(�U�;ǖ��\������q_����k[MZ6��I�����9i���"�V�u�^ʜ(�_��ȹ�R�#������c�����/zc;���Brt�"�1��v
�ً�0�A~��
�9-\���"
b���$�"n���ȡ�(m��H[K��<:��/����[['i�'#��]����8�h�Vb��A��о����b�e���*�xe�����, �p�l�n��a�@�a����ǡ�F1 ��K[H�DJ�dc�lǪ *w�m&�_;�5鏒fdW	�D}X=a�ǵ�M�gwc
(�-I��h#: O1# 40���`�I��
�}�; uQ|i�TN\����ʈ���i�Bh��n�9N�j2CðG-K2؟<s&F�-�ٝ��Ks�i�(^%*>ń�%B�g�6o����f9�a�,��S�nhx¸я��)в����G�Y��imÃ�8���AS�D�iEGV�uHv!��uTܩZ}9`'�֤��a�#���s��^�KY�*���Sl�fpl��~<U�+��Ũ(��o���<e4?�E�K <���Z�T��7
�q�ٽiϨ � M��{3,J�w/͍W������Z���.)Ʉ����84�v�A���B
z�d�)4�ļ��G"�t�+�@K��:�>Rn+���F�}�f��CR!:�	J��)Ǻ��⚹*ԣ������쏬̢8�w烗O�N�ХZ��>����it�S���a��1�V=�t��n�k�M�b�	|Fa�9	eb�ѻ�-�su�D�D�w�Ru!PZ��F�XC`��HCuf�	q.�6u�ƐsP��X���ᰄL�e�k������/����섿�B+�
�����y)�4���8���^"�P��D�X�D������c^d!:�QY�D�a�����+�K�������0�zEbX~�L�A�t� ��qw�*���*����[#�z�1��L�Ȉ-\P�m1lB�Xu�8��b��� �>�?X��$+��뻩����j�)�lj �a3�>0����w�o�X�