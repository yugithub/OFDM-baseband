��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f����qL��\|���@��#A����Lߡؘ��mO��|���jO��ϛ���6'���w���g��T�st�����U
��r��v�C��v[���v�Z��Ã�p�	���4$�g��d�2����90�Xyi��< $��d}��j������ !�ɏMn�f4�K���C��3�k����R6:�z��u�l����f��<��ƺ��W�H��g��qo�A���2/3���mM6�'��Zd8��7���G�>I>��ɢ�h��#$��
ҭ)��1>6�I}����H��k�M��3%��f^�����P] ���S~f"S����V�-�J� ���j1��6���/������!��E�Yz�ح<��=�:1��� �~W	�u���~
����R~轃G�鶖����Pt�D������?��ԓd_B��e�8�{�|�T��V��(�3�偻UCI״�g/�IP���0w��ݕXn0g��� Z�{k��X/I��j�@� E���$!����A��JL��(����S��V�\��)�N��n����w������[5@a,�*O��ě�w��N֌[R�L����H=���ѹ�^�Ǒ���F��Ԟ`��U�%�I���`7��FZ^C�{��2���::�[k��Y~���ft�+j<m��P�iT�%�>f�e�o�7e��W�$���ِ1��'��K�eM�>�~�⭧�njeH�s����B-�A*�.�cd¸�b[���.UE�@YH�#��t�����o.k,��zf�H�N���+�<Q�Ѽ�E��C�X2���ؘ���@��/>Z6�~bQ��"[�������K��k�?������"�F#>5��~J����A�H���J�J]� ::c��5�MxFn9�m�'��vwpJм�Qn^_���+L�5���(]`����1�D�K�C�<1y8��Y빑q��5)=~�wGk���Q܀y�iRuy�ѱ�a��8�^�f+8ԇW�����h��N�u�(-+Ѵ�,XctQ���se��s�R�P,��A�:�\(w�eVG IDl��Z��o-�:i	�&F�\B���2��0n|�_-O	B�b,�X%�f1>�����`U	�*��x��3�xpY%�%%.}#9,�)��ةa�a9E�lo3������ G��P7��9�_�!�$l:��ؘ^�ʼk�m��.p�9�4�zs�\u��/��t�'���/(#�,��a�6�)���i��悪��k����RJF����A�F��;��<�#H$OB��p�����ʚ�/|?a�|���&j \�#h6�aG�'a��k�N�����e���^y$�]��h�+���km��JE�w?O:{��1;����9f'5��>��k���,��W�tŖ�IL�7Me1��X��xHV��m:��ި�K��~���} �=T���dr��<���2����^x�R
ԉd�6*�heҺb+�\<��R}�-��󍜠%w��;�,�%\�^_C�p�B���s'��C�O̝�SD��	�O�sq���>�^�e��,G�y�"�"��v�Y��mC�"����Bk�Onq��r]I�Z���c��c8
�h�����G�����ـ�gx�r7>}��`	�!�)v�Ub�[g�2��c��� j��k�y����ָ��BHY;��v��7}�' �A�=���#�^�5V~|��Q��l0ߚvi�`��ʕ�� ������N��"s"nEa\͗I�Ȉ���)�l+֭��g��Ⱦ�ǆ]wc�0��0�!� �D�	2�]N�"��6��l�S Չ��ze�ިXlJ�4�y��L�=��K�f�.�邠钚�]� c;~b�Dp\��yp=i�� ��/i�8H��
�|0sT��C=�2u���'�lK[�tw	�Ԟ:�����&���`�
VD���:��	�]���w�\�y����
����)�D�j�L�"['���g����jkS<�B��h���-ej�@�2���ϣC*\ξ��uwY�L��*Zd�֙Ӂ�D�
�(,��7��蔽����CFI��B5oN����~ޣ�%�ͧ*lŧ�쐛z�o��s��8�����0�j��J��[Zc�����b�vg�dEKY�_:!�.�H��nxsN��7t���E� U�RR��
�$���
����]�1�M��J�I�p�^�a+x��ʑ��d�'���lǇ�GnҚR=�TT)�84o�խ5'6�n<��M�O�U�d��ჲ�g�-R��d
�N�t��c)���z��j�Ş�b�݌���`����������TI�e� C�5��&q�0����:�����R�H� ���P{q�#g��mM���)�	����9ء���#�f�؈t�Ҕ�\��c�% �ߜ��OvM	#]
� ,;2���M���ʦn43�L��l����NMk�q&5�&�t��#J���ő+��:�h8A���D��_���t;��vs����<�M;�O���i_Qf}	}hB���i*_}���Č��xfdȥ!I|��-�NL�b��U����'F���E�3>FX:|�3(껧/[2���Ԋ�������@"K���k��`��PKQ��3u�!_%U��XX��]P�3XF�d*��F�,�*�S��c�e�Gm�&as˳��CCZ]>�m��#���t-D���v�D�h�h�C?�{�����ưA��W��G�\%����j��O�X9 b$����϶��}��d�ME�Mğ�J�VG���'�wsS0,��8G?njms�/;�W�L�L����|�iY9����ۥހ��"jZт�g1P{Z�� 2G[sa �ɥ�p�(����L�Q�������*B�R�Xl�Q-R:��!�4��=���?�?Iz]����zj��qƖk�j[�;{~6N��p�!�ߞ��Q
��Pn�	~(�tg;��<�q��v���t��s��l�> F%hs&�/��Uŵ���ʘ�(�(����?�eTuj�V�s���v�������#����s(=��݄Hٴ���� +v�ʶ���1��?����
��+�]^���ti��d#V�`L����n�Tve	˵������]���gg7āl�k�!�Ǯ|��옟ƽ��'��\���&�0�u���Dj��h��SJDl��	N��i�:�a!�|�AR10õ����o�~ˑc���!�>]Q�Z�����b@��qu���z�@���l�o"��b��ˏ������c���$׼����=�EQ/d�����x!���dۡRС��Xlrz���֦T�d^N'�u
v����ք�Ľ��ٵ��!)$���� :����� ����ĕ�����c��@a��)"j������v|VKK��U�u�ֳO4���.��#��z�F�Y&�~C�V6���ȉ�~"<�@�.�k%*&�F��ʢ���>0䲴QV)��Ʃ��JX���1��tqCqp���d�2UHɠ����&:��o�PD`��3gĥĽ;p���C8y f�W�T.6L�P#h�a�Rp)�5$2��b��u�-:����x�.�� �6Q`���nO}���߫�uLcSd����[����D�
�U���]Q>sAvpN�`Ӡ�|j0 ��V&S&�Î�����1 �@@Q(z����w�Ƨ����U&��?&�>`g]��Ʌ�(	n��݂)�\#M;�(<FGW��-cQH�A�w��7y��YB����bIc-���WsjZ��g�`եr���(�,FC�'֎��-�:���O"Q�|�@{��5'#pS�v�Զ����b&�3-�mr�����j��)RO�$S��jbufۅ��o����fX�u��b1e};ۮ`������Q _�	Lp���m�\�YJ�Έ��Y�q+h�٭��[9rn����p�g	�(1�R�4=����w󋐇~��4S�����P���0�]V��9|��C�~�'�t�#�ݔ�U����iq�D���x���5���aTX�8rY!@�7�,*�z%)�� ���S��gP?` �X��a	=��īon�-"_T.޿8�XΎs�M�@oNw���Xeϋ�<�׽{zu�7���D^'� ����-��F��ڴ2o5��*R�$�at��k�����it��k���Xq[jp*��-~
0��穋Uc&�8�*��V�-�I��T�n����a�x/�����b��\��x~���Kdؚk*��^J��!N���-S�-�����fIzx�P1q$r3z7[�Tm�M#�V�}��������<*�:>��
��G��x1���d�}��	�@�O�W�����"�7���F6x��:�&g�[�Y�ekT��a�/tQVs�t��v�R�CM<�4o��I�?@9j��x"��h�5DH�������e�����o(ݫ5�+���2�#��7���}}������׼��`^c �UN�ͥ-��u�z��X��G]���h�6���a��`�s�K�c_���}�9
<�q��\26�ء�"���H�1\W�7T��?7�A��/E����Ǚ��{A�RG9�'�B�*�2�T78U����U��Xn��K�*-WV*�O"� Vf��ʥ�f�